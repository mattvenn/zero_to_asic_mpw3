magic
tech sky130A
magscale 1 2
timestamp 1635332755
<< metal1 >>
rect 191742 703332 191748 703384
rect 191800 703372 191806 703384
rect 283834 703372 283840 703384
rect 191800 703344 283840 703372
rect 191800 703332 191806 703344
rect 283834 703332 283840 703344
rect 283892 703332 283898 703384
rect 273898 703264 273904 703316
rect 273956 703304 273962 703316
rect 348786 703304 348792 703316
rect 273956 703276 348792 703304
rect 273956 703264 273962 703276
rect 348786 703264 348792 703276
rect 348844 703264 348850 703316
rect 215202 703196 215208 703248
rect 215260 703236 215266 703248
rect 364978 703236 364984 703248
rect 215260 703208 364984 703236
rect 215260 703196 215266 703208
rect 364978 703196 364984 703208
rect 365036 703196 365042 703248
rect 240778 703128 240784 703180
rect 240836 703168 240842 703180
rect 332502 703168 332508 703180
rect 240836 703140 332508 703168
rect 240836 703128 240842 703140
rect 332502 703128 332508 703140
rect 332560 703128 332566 703180
rect 249702 703060 249708 703112
rect 249760 703100 249766 703112
rect 413646 703100 413652 703112
rect 249760 703072 413652 703100
rect 249760 703060 249766 703072
rect 413646 703060 413652 703072
rect 413704 703060 413710 703112
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 220078 702992 220084 703044
rect 220136 703032 220142 703044
rect 267642 703032 267648 703044
rect 220136 703004 267648 703032
rect 220136 702992 220142 703004
rect 267642 702992 267648 703004
rect 267700 702992 267706 703044
rect 282178 702992 282184 703044
rect 282236 703032 282242 703044
rect 462314 703032 462320 703044
rect 282236 703004 462320 703032
rect 282236 702992 282242 703004
rect 462314 702992 462320 703004
rect 462372 702992 462378 703044
rect 104802 702924 104808 702976
rect 104860 702964 104866 702976
rect 300118 702964 300124 702976
rect 104860 702936 300124 702964
rect 104860 702924 104866 702936
rect 300118 702924 300124 702936
rect 300176 702924 300182 702976
rect 24302 702856 24308 702908
rect 24360 702896 24366 702908
rect 86218 702896 86224 702908
rect 24360 702868 86224 702896
rect 24360 702856 24366 702868
rect 86218 702856 86224 702868
rect 86276 702856 86282 702908
rect 90358 702856 90364 702908
rect 90416 702896 90422 702908
rect 235166 702896 235172 702908
rect 90416 702868 235172 702896
rect 90416 702856 90422 702868
rect 235166 702856 235172 702868
rect 235224 702856 235230 702908
rect 271138 702856 271144 702908
rect 271196 702896 271202 702908
rect 478506 702896 478512 702908
rect 271196 702868 478512 702896
rect 271196 702856 271202 702868
rect 478506 702856 478512 702868
rect 478564 702856 478570 702908
rect 70302 702788 70308 702840
rect 70360 702828 70366 702840
rect 154114 702828 154120 702840
rect 70360 702800 154120 702828
rect 70360 702788 70366 702800
rect 154114 702788 154120 702800
rect 154172 702788 154178 702840
rect 213178 702788 213184 702840
rect 213236 702828 213242 702840
rect 429838 702828 429844 702840
rect 213236 702800 429844 702828
rect 213236 702788 213242 702800
rect 429838 702788 429844 702800
rect 429896 702788 429902 702840
rect 40494 702720 40500 702772
rect 40552 702760 40558 702772
rect 94682 702760 94688 702772
rect 40552 702732 94688 702760
rect 40552 702720 40558 702732
rect 94682 702720 94688 702732
rect 94740 702720 94746 702772
rect 173802 702720 173808 702772
rect 173860 702760 173866 702772
rect 397454 702760 397460 702772
rect 173860 702732 397460 702760
rect 173860 702720 173866 702732
rect 397454 702720 397460 702732
rect 397512 702720 397518 702772
rect 8110 702652 8116 702704
rect 8168 702692 8174 702704
rect 96614 702692 96620 702704
rect 8168 702664 96620 702692
rect 8168 702652 8174 702664
rect 96614 702652 96620 702664
rect 96672 702652 96678 702704
rect 280798 702652 280804 702704
rect 280856 702692 280862 702704
rect 543458 702692 543464 702704
rect 280856 702664 543464 702692
rect 280856 702652 280862 702664
rect 543458 702652 543464 702664
rect 543516 702652 543522 702704
rect 84102 702584 84108 702636
rect 84160 702624 84166 702636
rect 202782 702624 202788 702636
rect 84160 702596 202788 702624
rect 84160 702584 84166 702596
rect 202782 702584 202788 702596
rect 202840 702584 202846 702636
rect 215938 702584 215944 702636
rect 215996 702624 216002 702636
rect 527082 702624 527088 702636
rect 215996 702596 527088 702624
rect 215996 702584 216002 702596
rect 527082 702584 527088 702596
rect 527140 702584 527146 702636
rect 66162 702516 66168 702568
rect 66220 702556 66226 702568
rect 170306 702556 170312 702568
rect 66220 702528 170312 702556
rect 66220 702516 66226 702528
rect 170306 702516 170312 702528
rect 170364 702516 170370 702568
rect 177942 702516 177948 702568
rect 178000 702556 178006 702568
rect 580902 702556 580908 702568
rect 178000 702528 580908 702556
rect 178000 702516 178006 702528
rect 580902 702516 580908 702528
rect 580960 702516 580966 702568
rect 77202 702448 77208 702500
rect 77260 702488 77266 702500
rect 494790 702488 494796 702500
rect 77260 702460 494796 702488
rect 77260 702448 77266 702460
rect 494790 702448 494796 702460
rect 494848 702448 494854 702500
rect 79962 700272 79968 700324
rect 80020 700312 80026 700324
rect 89162 700312 89168 700324
rect 80020 700284 89168 700312
rect 80020 700272 80026 700284
rect 89162 700272 89168 700284
rect 89220 700272 89226 700324
rect 218974 700272 218980 700324
rect 219032 700312 219038 700324
rect 241514 700312 241520 700324
rect 219032 700284 241520 700312
rect 219032 700272 219038 700284
rect 241514 700272 241520 700284
rect 241572 700272 241578 700324
rect 3418 683136 3424 683188
rect 3476 683176 3482 683188
rect 39298 683176 39304 683188
rect 3476 683148 39304 683176
rect 3476 683136 3482 683148
rect 39298 683136 39304 683148
rect 39356 683136 39362 683188
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 14458 670732 14464 670744
rect 3568 670704 14464 670732
rect 3568 670692 3574 670704
rect 14458 670692 14464 670704
rect 14516 670692 14522 670744
rect 3418 656888 3424 656940
rect 3476 656928 3482 656940
rect 74534 656928 74540 656940
rect 3476 656900 74540 656928
rect 3476 656888 3482 656900
rect 74534 656888 74540 656900
rect 74592 656888 74598 656940
rect 68922 625812 68928 625864
rect 68980 625852 68986 625864
rect 104894 625852 104900 625864
rect 68980 625824 104900 625852
rect 68980 625812 68986 625824
rect 104894 625812 104900 625824
rect 104952 625812 104958 625864
rect 3510 618264 3516 618316
rect 3568 618304 3574 618316
rect 11698 618304 11704 618316
rect 3568 618276 11704 618304
rect 3568 618264 3574 618276
rect 11698 618264 11704 618276
rect 11756 618264 11762 618316
rect 2774 605888 2780 605940
rect 2832 605928 2838 605940
rect 4798 605928 4804 605940
rect 2832 605900 4804 605928
rect 2832 605888 2838 605900
rect 4798 605888 4804 605900
rect 4856 605888 4862 605940
rect 79318 592016 79324 592068
rect 79376 592056 79382 592068
rect 79962 592056 79968 592068
rect 79376 592028 79968 592056
rect 79376 592016 79382 592028
rect 79962 592016 79968 592028
rect 80020 592056 80026 592068
rect 112438 592056 112444 592068
rect 80020 592028 112444 592056
rect 80020 592016 80026 592028
rect 112438 592016 112444 592028
rect 112496 592016 112502 592068
rect 76466 590384 76472 590436
rect 76524 590424 76530 590436
rect 77202 590424 77208 590436
rect 76524 590396 77208 590424
rect 76524 590384 76530 590396
rect 77202 590384 77208 590396
rect 77260 590384 77266 590436
rect 76466 589296 76472 589348
rect 76524 589336 76530 589348
rect 124398 589336 124404 589348
rect 76524 589308 124404 589336
rect 76524 589296 76530 589308
rect 124398 589296 124404 589308
rect 124456 589296 124462 589348
rect 67726 588344 67732 588396
rect 67784 588384 67790 588396
rect 68922 588384 68928 588396
rect 67784 588356 68928 588384
rect 67784 588344 67790 588356
rect 68922 588344 68928 588356
rect 68980 588344 68986 588396
rect 68922 587868 68928 587920
rect 68980 587908 68986 587920
rect 128354 587908 128360 587920
rect 68980 587880 128360 587908
rect 68980 587868 68986 587880
rect 128354 587868 128360 587880
rect 128412 587868 128418 587920
rect 81802 587188 81808 587240
rect 81860 587228 81866 587240
rect 84102 587228 84108 587240
rect 81860 587200 84108 587228
rect 81860 587188 81866 587200
rect 84102 587188 84108 587200
rect 84160 587228 84166 587240
rect 143534 587228 143540 587240
rect 84160 587200 143540 587228
rect 84160 587188 84166 587200
rect 143534 587188 143540 587200
rect 143592 587188 143598 587240
rect 4798 587120 4804 587172
rect 4856 587160 4862 587172
rect 96706 587160 96712 587172
rect 4856 587132 96712 587160
rect 4856 587120 4862 587132
rect 96706 587120 96712 587132
rect 96764 587120 96770 587172
rect 121454 585760 121460 585812
rect 121512 585800 121518 585812
rect 582834 585800 582840 585812
rect 121512 585772 582840 585800
rect 121512 585760 121518 585772
rect 582834 585760 582840 585772
rect 582892 585760 582898 585812
rect 87506 585216 87512 585268
rect 87564 585256 87570 585268
rect 121454 585256 121460 585268
rect 87564 585228 121460 585256
rect 87564 585216 87570 585228
rect 121454 585216 121460 585228
rect 121512 585216 121518 585268
rect 72418 585148 72424 585200
rect 72476 585188 72482 585200
rect 116578 585188 116584 585200
rect 72476 585160 116584 585188
rect 72476 585148 72482 585160
rect 116578 585148 116584 585160
rect 116636 585148 116642 585200
rect 74258 583788 74264 583840
rect 74316 583828 74322 583840
rect 98638 583828 98644 583840
rect 74316 583800 98644 583828
rect 74316 583788 74322 583800
rect 98638 583788 98644 583800
rect 98696 583788 98702 583840
rect 88242 583720 88248 583772
rect 88300 583760 88306 583772
rect 115198 583760 115204 583772
rect 88300 583732 115204 583760
rect 88300 583720 88306 583732
rect 115198 583720 115204 583732
rect 115256 583720 115262 583772
rect 78122 582632 78128 582684
rect 78180 582672 78186 582684
rect 79318 582672 79324 582684
rect 78180 582644 79324 582672
rect 78180 582632 78186 582644
rect 79318 582632 79324 582644
rect 79376 582632 79382 582684
rect 57882 582564 57888 582616
rect 57940 582604 57946 582616
rect 90450 582604 90456 582616
rect 57940 582576 90456 582604
rect 57940 582564 57946 582576
rect 90450 582564 90456 582576
rect 90508 582564 90514 582616
rect 86218 582496 86224 582548
rect 86276 582536 86282 582548
rect 100202 582536 100208 582548
rect 86276 582508 100208 582536
rect 86276 582496 86282 582508
rect 100202 582496 100208 582508
rect 100260 582496 100266 582548
rect 50982 582428 50988 582480
rect 51040 582468 51046 582480
rect 69934 582468 69940 582480
rect 51040 582440 69940 582468
rect 51040 582428 51046 582440
rect 69934 582428 69940 582440
rect 69992 582428 69998 582480
rect 79042 582360 79048 582412
rect 79100 582400 79106 582412
rect 86862 582400 86868 582412
rect 79100 582372 86868 582400
rect 79100 582360 79106 582372
rect 86862 582360 86868 582372
rect 86920 582360 86926 582412
rect 90266 582360 90272 582412
rect 90324 582400 90330 582412
rect 95970 582400 95976 582412
rect 90324 582372 95976 582400
rect 90324 582360 90330 582372
rect 95970 582360 95976 582372
rect 96028 582360 96034 582412
rect 76282 581068 76288 581120
rect 76340 581108 76346 581120
rect 108298 581108 108304 581120
rect 76340 581080 108304 581108
rect 76340 581068 76346 581080
rect 108298 581068 108304 581080
rect 108356 581068 108362 581120
rect 59262 581000 59268 581052
rect 59320 581040 59326 581052
rect 82998 581040 83004 581052
rect 59320 581012 83004 581040
rect 59320 581000 59326 581012
rect 82998 581000 83004 581012
rect 83056 581000 83062 581052
rect 93762 581000 93768 581052
rect 93820 581040 93826 581052
rect 148318 581040 148324 581052
rect 93820 581012 148324 581040
rect 93820 581000 93826 581012
rect 148318 581000 148324 581012
rect 148376 581000 148382 581052
rect 69014 580660 69020 580712
rect 69072 580660 69078 580712
rect 86862 580660 86868 580712
rect 86920 580700 86926 580712
rect 86920 580672 93854 580700
rect 86920 580660 86926 580672
rect 3510 580184 3516 580236
rect 3568 580224 3574 580236
rect 8110 580224 8116 580236
rect 3568 580196 8116 580224
rect 3568 580184 3574 580196
rect 8110 580184 8116 580196
rect 8168 580184 8174 580236
rect 64782 579708 64788 579760
rect 64840 579748 64846 579760
rect 66530 579748 66536 579760
rect 64840 579720 66536 579748
rect 64840 579708 64846 579720
rect 66530 579708 66536 579720
rect 66588 579708 66594 579760
rect 53558 579640 53564 579692
rect 53616 579680 53622 579692
rect 69032 579680 69060 580660
rect 93826 580292 93854 580672
rect 94682 580456 94688 580508
rect 94740 580496 94746 580508
rect 95878 580496 95884 580508
rect 94740 580468 95884 580496
rect 94740 580456 94746 580468
rect 95878 580456 95884 580468
rect 95936 580456 95942 580508
rect 102778 580292 102784 580304
rect 93826 580264 102784 580292
rect 102778 580252 102784 580264
rect 102836 580252 102842 580304
rect 53616 579652 69060 579680
rect 53616 579640 53622 579652
rect 97166 578212 97172 578264
rect 97224 578252 97230 578264
rect 134518 578252 134524 578264
rect 97224 578224 134524 578252
rect 97224 578212 97230 578224
rect 134518 578212 134524 578224
rect 134576 578212 134582 578264
rect 97166 576852 97172 576904
rect 97224 576892 97230 576904
rect 122834 576892 122840 576904
rect 97224 576864 122840 576892
rect 97224 576852 97230 576864
rect 122834 576852 122840 576864
rect 122892 576852 122898 576904
rect 187602 576852 187608 576904
rect 187660 576892 187666 576904
rect 580166 576892 580172 576904
rect 187660 576864 580172 576892
rect 187660 576852 187666 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 3418 576784 3424 576836
rect 3476 576824 3482 576836
rect 67634 576824 67640 576836
rect 3476 576796 67640 576824
rect 3476 576784 3482 576796
rect 67634 576784 67640 576796
rect 67692 576784 67698 576836
rect 97902 576104 97908 576156
rect 97960 576144 97966 576156
rect 104802 576144 104808 576156
rect 97960 576116 104808 576144
rect 97960 576104 97966 576116
rect 104802 576104 104808 576116
rect 104860 576144 104866 576156
rect 125594 576144 125600 576156
rect 104860 576116 125600 576144
rect 104860 576104 104866 576116
rect 125594 576104 125600 576116
rect 125652 576104 125658 576156
rect 95970 574744 95976 574796
rect 96028 574784 96034 574796
rect 104158 574784 104164 574796
rect 96028 574756 104164 574784
rect 96028 574744 96034 574756
rect 104158 574744 104164 574756
rect 104216 574744 104222 574796
rect 95878 573316 95884 573368
rect 95936 573356 95942 573368
rect 120074 573356 120080 573368
rect 95936 573328 120080 573356
rect 95936 573316 95942 573328
rect 120074 573316 120080 573328
rect 120132 573316 120138 573368
rect 63402 572704 63408 572756
rect 63460 572744 63466 572756
rect 66530 572744 66536 572756
rect 63460 572716 66536 572744
rect 63460 572704 63466 572716
rect 66530 572704 66536 572716
rect 66588 572704 66594 572756
rect 41322 571344 41328 571396
rect 41380 571384 41386 571396
rect 66530 571384 66536 571396
rect 41380 571356 66536 571384
rect 41380 571344 41386 571356
rect 66530 571344 66536 571356
rect 66588 571344 66594 571396
rect 96798 571344 96804 571396
rect 96856 571384 96862 571396
rect 106918 571384 106924 571396
rect 96856 571356 106924 571384
rect 96856 571344 96862 571356
rect 106918 571344 106924 571356
rect 106976 571344 106982 571396
rect 61930 569984 61936 570036
rect 61988 570024 61994 570036
rect 66898 570024 66904 570036
rect 61988 569996 66904 570024
rect 61988 569984 61994 569996
rect 66898 569984 66904 569996
rect 66956 569984 66962 570036
rect 97902 569916 97908 569968
rect 97960 569956 97966 569968
rect 115290 569956 115296 569968
rect 97960 569928 115296 569956
rect 97960 569916 97966 569928
rect 115290 569916 115296 569928
rect 115348 569916 115354 569968
rect 97902 568624 97908 568676
rect 97960 568664 97966 568676
rect 104434 568664 104440 568676
rect 97960 568636 104440 568664
rect 97960 568624 97966 568636
rect 104434 568624 104440 568636
rect 104492 568624 104498 568676
rect 62022 565836 62028 565888
rect 62080 565876 62086 565888
rect 66162 565876 66168 565888
rect 62080 565848 66168 565876
rect 62080 565836 62086 565848
rect 66162 565836 66168 565848
rect 66220 565836 66226 565888
rect 56502 564408 56508 564460
rect 56560 564448 56566 564460
rect 66530 564448 66536 564460
rect 56560 564420 66536 564448
rect 56560 564408 56566 564420
rect 66530 564408 66536 564420
rect 66588 564408 66594 564460
rect 52362 563048 52368 563100
rect 52420 563088 52426 563100
rect 66530 563088 66536 563100
rect 52420 563060 66536 563088
rect 52420 563048 52426 563060
rect 66530 563048 66536 563060
rect 66588 563048 66594 563100
rect 107010 562912 107016 562964
rect 107068 562952 107074 562964
rect 111058 562952 111064 562964
rect 107068 562924 111064 562952
rect 107068 562912 107074 562924
rect 111058 562912 111064 562924
rect 111116 562912 111122 562964
rect 96798 561688 96804 561740
rect 96856 561728 96862 561740
rect 117314 561728 117320 561740
rect 96856 561700 117320 561728
rect 96856 561688 96862 561700
rect 117314 561688 117320 561700
rect 117372 561688 117378 561740
rect 48038 560260 48044 560312
rect 48096 560300 48102 560312
rect 66714 560300 66720 560312
rect 48096 560272 66720 560300
rect 48096 560260 48102 560272
rect 66714 560260 66720 560272
rect 66772 560260 66778 560312
rect 48222 558900 48228 558952
rect 48280 558940 48286 558952
rect 66714 558940 66720 558952
rect 48280 558912 66720 558940
rect 48280 558900 48286 558912
rect 66714 558900 66720 558912
rect 66772 558900 66778 558952
rect 96798 558900 96804 558952
rect 96856 558940 96862 558952
rect 112714 558940 112720 558952
rect 96856 558912 112720 558940
rect 96856 558900 96862 558912
rect 112714 558900 112720 558912
rect 112772 558900 112778 558952
rect 44082 557540 44088 557592
rect 44140 557580 44146 557592
rect 66714 557580 66720 557592
rect 44140 557552 66720 557580
rect 44140 557540 44146 557552
rect 66714 557540 66720 557552
rect 66772 557540 66778 557592
rect 96982 554752 96988 554804
rect 97040 554792 97046 554804
rect 129734 554792 129740 554804
rect 97040 554764 129740 554792
rect 97040 554752 97046 554764
rect 129734 554752 129740 554764
rect 129792 554752 129798 554804
rect 3326 553392 3332 553444
rect 3384 553432 3390 553444
rect 29638 553432 29644 553444
rect 3384 553404 29644 553432
rect 3384 553392 3390 553404
rect 29638 553392 29644 553404
rect 29696 553392 29702 553444
rect 57790 553392 57796 553444
rect 57848 553432 57854 553444
rect 66530 553432 66536 553444
rect 57848 553404 66536 553432
rect 57848 553392 57854 553404
rect 66530 553392 66536 553404
rect 66588 553392 66594 553444
rect 96982 552032 96988 552084
rect 97040 552072 97046 552084
rect 108482 552072 108488 552084
rect 97040 552044 108488 552072
rect 97040 552032 97046 552044
rect 108482 552032 108488 552044
rect 108540 552032 108546 552084
rect 97902 550604 97908 550656
rect 97960 550644 97966 550656
rect 115934 550644 115940 550656
rect 97960 550616 115940 550644
rect 97960 550604 97966 550616
rect 115934 550604 115940 550616
rect 115992 550604 115998 550656
rect 55122 549244 55128 549296
rect 55180 549284 55186 549296
rect 66530 549284 66536 549296
rect 55180 549256 66536 549284
rect 55180 549244 55186 549256
rect 66530 549244 66536 549256
rect 66588 549244 66594 549296
rect 64690 547884 64696 547936
rect 64748 547924 64754 547936
rect 66806 547924 66812 547936
rect 64748 547896 66812 547924
rect 64748 547884 64754 547896
rect 66806 547884 66812 547896
rect 66864 547884 66870 547936
rect 63310 545096 63316 545148
rect 63368 545136 63374 545148
rect 66714 545136 66720 545148
rect 63368 545108 66720 545136
rect 63368 545096 63374 545108
rect 66714 545096 66720 545108
rect 66772 545096 66778 545148
rect 97074 543736 97080 543788
rect 97132 543776 97138 543788
rect 104342 543776 104348 543788
rect 97132 543748 104348 543776
rect 97132 543736 97138 543748
rect 104342 543736 104348 543748
rect 104400 543736 104406 543788
rect 39298 543668 39304 543720
rect 39356 543708 39362 543720
rect 67266 543708 67272 543720
rect 39356 543680 67272 543708
rect 39356 543668 39362 543680
rect 67266 543668 67272 543680
rect 67324 543668 67330 543720
rect 97166 540948 97172 541000
rect 97224 540988 97230 541000
rect 130378 540988 130384 541000
rect 97224 540960 130384 540988
rect 97224 540948 97230 540960
rect 130378 540948 130384 540960
rect 130436 540948 130442 541000
rect 11698 540200 11704 540252
rect 11756 540240 11762 540252
rect 11756 540212 64874 540240
rect 11756 540200 11762 540212
rect 64846 539832 64874 540212
rect 73154 539832 73160 539844
rect 64846 539804 73160 539832
rect 73154 539792 73160 539804
rect 73212 539792 73218 539844
rect 91002 539792 91008 539844
rect 91060 539832 91066 539844
rect 96706 539832 96712 539844
rect 91060 539804 96712 539832
rect 91060 539792 91066 539804
rect 96706 539792 96712 539804
rect 96764 539792 96770 539844
rect 59170 539588 59176 539640
rect 59228 539628 59234 539640
rect 66438 539628 66444 539640
rect 59228 539600 66444 539628
rect 59228 539588 59234 539600
rect 66438 539588 66444 539600
rect 66496 539588 66502 539640
rect 86218 539588 86224 539640
rect 86276 539628 86282 539640
rect 94314 539628 94320 539640
rect 86276 539600 94320 539628
rect 86276 539588 86282 539600
rect 94314 539588 94320 539600
rect 94372 539588 94378 539640
rect 67818 539044 67824 539096
rect 67876 539084 67882 539096
rect 71866 539084 71872 539096
rect 67876 539056 71872 539084
rect 67876 539044 67882 539056
rect 71866 539044 71872 539056
rect 71924 539044 71930 539096
rect 82722 538840 82728 538892
rect 82780 538880 82786 538892
rect 95510 538880 95516 538892
rect 82780 538852 95516 538880
rect 82780 538840 82786 538852
rect 95510 538840 95516 538852
rect 95568 538840 95574 538892
rect 4798 538228 4804 538280
rect 4856 538268 4862 538280
rect 93946 538268 93952 538280
rect 4856 538240 93952 538268
rect 4856 538228 4862 538240
rect 93946 538228 93952 538240
rect 94004 538228 94010 538280
rect 29638 538160 29644 538212
rect 29696 538200 29702 538212
rect 70670 538200 70676 538212
rect 29696 538172 70676 538200
rect 29696 538160 29702 538172
rect 70670 538160 70676 538172
rect 70728 538160 70734 538212
rect 90358 538160 90364 538212
rect 90416 538200 90422 538212
rect 136634 538200 136640 538212
rect 90416 538172 136640 538200
rect 90416 538160 90422 538172
rect 136634 538160 136640 538172
rect 136692 538160 136698 538212
rect 75822 537480 75828 537532
rect 75880 537520 75886 537532
rect 96890 537520 96896 537532
rect 75880 537492 96896 537520
rect 75880 537480 75886 537492
rect 96890 537480 96896 537492
rect 96948 537480 96954 537532
rect 3418 536732 3424 536784
rect 3476 536772 3482 536784
rect 69014 536772 69020 536784
rect 3476 536744 69020 536772
rect 3476 536732 3482 536744
rect 69014 536732 69020 536744
rect 69072 536732 69078 536784
rect 73430 536732 73436 536784
rect 73488 536772 73494 536784
rect 76558 536772 76564 536784
rect 73488 536744 76564 536772
rect 73488 536732 73494 536744
rect 76558 536732 76564 536744
rect 76616 536732 76622 536784
rect 82170 536120 82176 536172
rect 82228 536160 82234 536172
rect 95326 536160 95332 536172
rect 82228 536132 95332 536160
rect 82228 536120 82234 536132
rect 95326 536120 95332 536132
rect 95384 536120 95390 536172
rect 67726 536052 67732 536104
rect 67784 536092 67790 536104
rect 83458 536092 83464 536104
rect 67784 536064 83464 536092
rect 67784 536052 67790 536064
rect 83458 536052 83464 536064
rect 83516 536052 83522 536104
rect 86678 535508 86684 535560
rect 86736 535548 86742 535560
rect 87690 535548 87696 535560
rect 86736 535520 87696 535548
rect 86736 535508 86742 535520
rect 87690 535508 87696 535520
rect 87748 535508 87754 535560
rect 50798 534692 50804 534744
rect 50856 534732 50862 534744
rect 87138 534732 87144 534744
rect 50856 534704 87144 534732
rect 50856 534692 50862 534704
rect 87138 534692 87144 534704
rect 87196 534692 87202 534744
rect 88334 533400 88340 533452
rect 88392 533440 88398 533452
rect 88886 533440 88892 533452
rect 88392 533412 88892 533440
rect 88392 533400 88398 533412
rect 88886 533400 88892 533412
rect 88944 533400 88950 533452
rect 91094 533400 91100 533452
rect 91152 533440 91158 533452
rect 91830 533440 91836 533452
rect 91152 533412 91836 533440
rect 91152 533400 91158 533412
rect 91830 533400 91836 533412
rect 91888 533400 91894 533452
rect 55030 533332 55036 533384
rect 55088 533372 55094 533384
rect 96798 533372 96804 533384
rect 55088 533344 96804 533372
rect 55088 533332 55094 533344
rect 96798 533332 96804 533344
rect 96856 533332 96862 533384
rect 65886 531972 65892 532024
rect 65944 532012 65950 532024
rect 107010 532012 107016 532024
rect 65944 531984 107016 532012
rect 65944 531972 65950 531984
rect 107010 531972 107016 531984
rect 107068 531972 107074 532024
rect 93762 531224 93768 531276
rect 93820 531264 93826 531276
rect 94498 531264 94504 531276
rect 93820 531236 94504 531264
rect 93820 531224 93826 531236
rect 94498 531224 94504 531236
rect 94556 531224 94562 531276
rect 70670 530544 70676 530596
rect 70728 530584 70734 530596
rect 141418 530584 141424 530596
rect 70728 530556 141424 530584
rect 70728 530544 70734 530556
rect 141418 530544 141424 530556
rect 141476 530544 141482 530596
rect 3418 529184 3424 529236
rect 3476 529224 3482 529236
rect 93762 529224 93768 529236
rect 3476 529196 93768 529224
rect 3476 529184 3482 529196
rect 93762 529184 93768 529196
rect 93820 529184 93826 529236
rect 3510 527824 3516 527876
rect 3568 527864 3574 527876
rect 122834 527864 122840 527876
rect 3568 527836 122840 527864
rect 3568 527824 3574 527836
rect 122834 527824 122840 527836
rect 122892 527824 122898 527876
rect 64598 526396 64604 526448
rect 64656 526436 64662 526448
rect 84194 526436 84200 526448
rect 64656 526408 84200 526436
rect 64656 526396 64662 526408
rect 84194 526396 84200 526408
rect 84252 526396 84258 526448
rect 67358 525036 67364 525088
rect 67416 525076 67422 525088
rect 113174 525076 113180 525088
rect 67416 525048 113180 525076
rect 67416 525036 67422 525048
rect 113174 525036 113180 525048
rect 113232 525036 113238 525088
rect 104342 521568 104348 521620
rect 104400 521608 104406 521620
rect 108390 521608 108396 521620
rect 104400 521580 108396 521608
rect 104400 521568 104406 521580
rect 108390 521568 108396 521580
rect 108448 521568 108454 521620
rect 64690 520888 64696 520940
rect 64748 520928 64754 520940
rect 69658 520928 69664 520940
rect 64748 520900 69664 520928
rect 64748 520888 64754 520900
rect 69658 520888 69664 520900
rect 69716 520888 69722 520940
rect 53650 518168 53656 518220
rect 53708 518208 53714 518220
rect 97994 518208 98000 518220
rect 53708 518180 98000 518208
rect 53708 518168 53714 518180
rect 97994 518168 98000 518180
rect 98052 518168 98058 518220
rect 3510 514768 3516 514820
rect 3568 514808 3574 514820
rect 7558 514808 7564 514820
rect 3568 514780 7564 514808
rect 3568 514768 3574 514780
rect 7558 514768 7564 514780
rect 7616 514768 7622 514820
rect 108482 506948 108488 507000
rect 108540 506988 108546 507000
rect 112530 506988 112536 507000
rect 108540 506960 112536 506988
rect 108540 506948 108546 506960
rect 112530 506948 112536 506960
rect 112588 506948 112594 507000
rect 66070 501576 66076 501628
rect 66128 501616 66134 501628
rect 125778 501616 125784 501628
rect 66128 501588 125784 501616
rect 66128 501576 66134 501588
rect 125778 501576 125784 501588
rect 125836 501576 125842 501628
rect 88426 498788 88432 498840
rect 88484 498828 88490 498840
rect 124306 498828 124312 498840
rect 88484 498800 124312 498828
rect 88484 498788 88490 498800
rect 124306 498788 124312 498800
rect 124364 498788 124370 498840
rect 63310 496068 63316 496120
rect 63368 496108 63374 496120
rect 123478 496108 123484 496120
rect 63368 496080 123484 496108
rect 63368 496068 63374 496080
rect 123478 496068 123484 496080
rect 123536 496068 123542 496120
rect 76558 493280 76564 493332
rect 76616 493320 76622 493332
rect 102870 493320 102876 493332
rect 76616 493292 102876 493320
rect 76616 493280 76622 493292
rect 102870 493280 102876 493292
rect 102928 493280 102934 493332
rect 64782 490560 64788 490612
rect 64840 490600 64846 490612
rect 92474 490600 92480 490612
rect 64840 490572 92480 490600
rect 64840 490560 64846 490572
rect 92474 490560 92480 490572
rect 92532 490560 92538 490612
rect 73798 487772 73804 487824
rect 73856 487812 73862 487824
rect 99374 487812 99380 487824
rect 73856 487784 99380 487812
rect 73856 487772 73862 487784
rect 99374 487772 99380 487784
rect 99432 487772 99438 487824
rect 102134 487772 102140 487824
rect 102192 487812 102198 487824
rect 102778 487812 102784 487824
rect 102192 487784 102784 487812
rect 102192 487772 102198 487784
rect 102778 487772 102784 487784
rect 102836 487812 102842 487824
rect 240778 487812 240784 487824
rect 102836 487784 240784 487812
rect 102836 487772 102842 487784
rect 240778 487772 240784 487784
rect 240836 487772 240842 487824
rect 77294 486412 77300 486464
rect 77352 486452 77358 486464
rect 108482 486452 108488 486464
rect 77352 486424 108488 486452
rect 77352 486412 77358 486424
rect 108482 486412 108488 486424
rect 108540 486412 108546 486464
rect 77938 485052 77944 485104
rect 77996 485092 78002 485104
rect 91186 485092 91192 485104
rect 77996 485064 91192 485092
rect 77996 485052 78002 485064
rect 91186 485052 91192 485064
rect 91244 485052 91250 485104
rect 188982 484372 188988 484424
rect 189040 484412 189046 484424
rect 580166 484412 580172 484424
rect 189040 484384 580172 484412
rect 189040 484372 189046 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 112438 483624 112444 483676
rect 112496 483664 112502 483676
rect 125686 483664 125692 483676
rect 112496 483636 125692 483664
rect 112496 483624 112502 483636
rect 125686 483624 125692 483636
rect 125744 483624 125750 483676
rect 87690 481584 87696 481636
rect 87748 481624 87754 481636
rect 88242 481624 88248 481636
rect 87748 481596 88248 481624
rect 87748 481584 87754 481596
rect 88242 481584 88248 481596
rect 88300 481584 88306 481636
rect 241514 481584 241520 481636
rect 241572 481624 241578 481636
rect 242158 481624 242164 481636
rect 241572 481596 242164 481624
rect 241572 481584 241578 481596
rect 242158 481584 242164 481596
rect 242216 481584 242222 481636
rect 88242 480904 88248 480956
rect 88300 480944 88306 480956
rect 242158 480944 242164 480956
rect 88300 480916 242164 480944
rect 88300 480904 88306 480916
rect 242158 480904 242164 480916
rect 242216 480904 242222 480956
rect 67726 479476 67732 479528
rect 67784 479516 67790 479528
rect 96982 479516 96988 479528
rect 67784 479488 96988 479516
rect 67784 479476 67790 479488
rect 96982 479476 96988 479488
rect 97040 479476 97046 479528
rect 90450 478864 90456 478916
rect 90508 478904 90514 478916
rect 91002 478904 91008 478916
rect 90508 478876 91008 478904
rect 90508 478864 90514 478876
rect 91002 478864 91008 478876
rect 91060 478904 91066 478916
rect 218054 478904 218060 478916
rect 91060 478876 218060 478904
rect 91060 478864 91066 478876
rect 218054 478864 218060 478876
rect 218112 478864 218118 478916
rect 106918 478116 106924 478168
rect 106976 478156 106982 478168
rect 128446 478156 128452 478168
rect 106976 478128 128452 478156
rect 106976 478116 106982 478128
rect 128446 478116 128452 478128
rect 128504 478116 128510 478168
rect 2774 476076 2780 476128
rect 2832 476116 2838 476128
rect 3418 476116 3424 476128
rect 2832 476088 3424 476116
rect 2832 476076 2838 476088
rect 3418 476076 3424 476088
rect 3476 476116 3482 476128
rect 4798 476116 4804 476128
rect 3476 476088 4804 476116
rect 3476 476076 3482 476088
rect 4798 476076 4804 476088
rect 4856 476076 4862 476128
rect 104158 476076 104164 476128
rect 104216 476116 104222 476128
rect 241514 476116 241520 476128
rect 104216 476088 241520 476116
rect 104216 476076 104222 476088
rect 241514 476076 241520 476088
rect 241572 476076 241578 476128
rect 78674 475396 78680 475448
rect 78732 475436 78738 475448
rect 98730 475436 98736 475448
rect 78732 475408 98736 475436
rect 78732 475396 78738 475408
rect 98730 475396 98736 475408
rect 98788 475396 98794 475448
rect 98638 475328 98644 475380
rect 98696 475368 98702 475380
rect 121546 475368 121552 475380
rect 98696 475340 121552 475368
rect 98696 475328 98702 475340
rect 121546 475328 121552 475340
rect 121604 475328 121610 475380
rect 104250 475192 104256 475244
rect 104308 475232 104314 475244
rect 104802 475232 104808 475244
rect 104308 475204 104808 475232
rect 104308 475192 104314 475204
rect 104802 475192 104808 475204
rect 104860 475192 104866 475244
rect 104802 474716 104808 474768
rect 104860 474756 104866 474768
rect 255406 474756 255412 474768
rect 104860 474728 255412 474756
rect 104860 474716 104866 474728
rect 255406 474716 255412 474728
rect 255464 474716 255470 474768
rect 93946 473832 93952 473884
rect 94004 473872 94010 473884
rect 94682 473872 94688 473884
rect 94004 473844 94688 473872
rect 94004 473832 94010 473844
rect 94682 473832 94688 473844
rect 94740 473832 94746 473884
rect 94682 473356 94688 473408
rect 94740 473396 94746 473408
rect 227806 473396 227812 473408
rect 94740 473368 227812 473396
rect 94740 473356 94746 473368
rect 227806 473356 227812 473368
rect 227864 473356 227870 473408
rect 88334 472608 88340 472660
rect 88392 472648 88398 472660
rect 118694 472648 118700 472660
rect 88392 472620 118700 472648
rect 88392 472608 88398 472620
rect 118694 472608 118700 472620
rect 118752 472608 118758 472660
rect 118694 471996 118700 472048
rect 118752 472036 118758 472048
rect 255590 472036 255596 472048
rect 118752 472008 255596 472036
rect 118752 471996 118758 472008
rect 255590 471996 255596 472008
rect 255648 471996 255654 472048
rect 108482 471248 108488 471300
rect 108540 471288 108546 471300
rect 117406 471288 117412 471300
rect 108540 471260 117412 471288
rect 108540 471248 108546 471260
rect 117406 471248 117412 471260
rect 117464 471248 117470 471300
rect 117406 470568 117412 470620
rect 117464 470608 117470 470620
rect 262214 470608 262220 470620
rect 117464 470580 262220 470608
rect 117464 470568 117470 470580
rect 262214 470568 262220 470580
rect 262272 470568 262278 470620
rect 82814 469820 82820 469872
rect 82872 469860 82878 469872
rect 109678 469860 109684 469872
rect 82872 469832 109684 469860
rect 82872 469820 82878 469832
rect 109678 469820 109684 469832
rect 109736 469820 109742 469872
rect 159358 469276 159364 469328
rect 159416 469316 159422 469328
rect 253934 469316 253940 469328
rect 159416 469288 253940 469316
rect 159416 469276 159422 469288
rect 253934 469276 253940 469288
rect 253992 469276 253998 469328
rect 112438 469208 112444 469260
rect 112496 469248 112502 469260
rect 142890 469248 142896 469260
rect 112496 469220 142896 469248
rect 112496 469208 112502 469220
rect 142890 469208 142896 469220
rect 142948 469248 142954 469260
rect 252554 469248 252560 469260
rect 142948 469220 252560 469248
rect 142948 469208 142954 469220
rect 252554 469208 252560 469220
rect 252612 469208 252618 469260
rect 71682 468528 71688 468580
rect 71740 468568 71746 468580
rect 91094 468568 91100 468580
rect 71740 468540 91100 468568
rect 71740 468528 71746 468540
rect 91094 468528 91100 468540
rect 91152 468528 91158 468580
rect 85574 468460 85580 468512
rect 85632 468500 85638 468512
rect 113358 468500 113364 468512
rect 85632 468472 113364 468500
rect 85632 468460 85638 468472
rect 113358 468460 113364 468472
rect 113416 468460 113422 468512
rect 108390 467848 108396 467900
rect 108448 467888 108454 467900
rect 245654 467888 245660 467900
rect 108448 467860 245660 467888
rect 108448 467848 108454 467860
rect 245654 467848 245660 467860
rect 245712 467848 245718 467900
rect 82722 466488 82728 466540
rect 82780 466528 82786 466540
rect 211154 466528 211160 466540
rect 82780 466500 211160 466528
rect 82780 466488 82786 466500
rect 211154 466488 211160 466500
rect 211212 466488 211218 466540
rect 102410 466420 102416 466472
rect 102468 466460 102474 466472
rect 102870 466460 102876 466472
rect 102468 466432 102876 466460
rect 102468 466420 102474 466432
rect 102870 466420 102876 466432
rect 102928 466460 102934 466472
rect 240870 466460 240876 466472
rect 102928 466432 240876 466460
rect 102928 466420 102934 466432
rect 240870 466420 240876 466432
rect 240928 466420 240934 466472
rect 87598 465672 87604 465724
rect 87656 465712 87662 465724
rect 126974 465712 126980 465724
rect 87656 465684 126980 465712
rect 87656 465672 87662 465684
rect 126974 465672 126980 465684
rect 127032 465672 127038 465724
rect 188338 465128 188344 465180
rect 188396 465168 188402 465180
rect 256694 465168 256700 465180
rect 188396 465140 256700 465168
rect 188396 465128 188402 465140
rect 256694 465128 256700 465140
rect 256752 465128 256758 465180
rect 137278 465060 137284 465112
rect 137336 465100 137342 465112
rect 240134 465100 240140 465112
rect 137336 465072 240140 465100
rect 137336 465060 137342 465072
rect 240134 465060 240140 465072
rect 240192 465060 240198 465112
rect 57698 464992 57704 465044
rect 57756 465032 57762 465044
rect 57882 465032 57888 465044
rect 57756 465004 57888 465032
rect 57756 464992 57762 465004
rect 57882 464992 57888 465004
rect 57940 464992 57946 465044
rect 86862 464312 86868 464364
rect 86920 464352 86926 464364
rect 95234 464352 95240 464364
rect 86920 464324 95240 464352
rect 86920 464312 86926 464324
rect 95234 464312 95240 464324
rect 95292 464312 95298 464364
rect 141418 463768 141424 463820
rect 141476 463808 141482 463820
rect 259546 463808 259552 463820
rect 141476 463780 259552 463808
rect 141476 463768 141482 463780
rect 259546 463768 259552 463780
rect 259604 463768 259610 463820
rect 57698 463700 57704 463752
rect 57756 463740 57762 463752
rect 186958 463740 186964 463752
rect 57756 463712 186964 463740
rect 57756 463700 57762 463712
rect 186958 463700 186964 463712
rect 187016 463700 187022 463752
rect 191190 463700 191196 463752
rect 191248 463740 191254 463752
rect 231118 463740 231124 463752
rect 191248 463712 231124 463740
rect 191248 463700 191254 463712
rect 231118 463700 231124 463712
rect 231176 463700 231182 463752
rect 77202 462952 77208 463004
rect 77260 462992 77266 463004
rect 90358 462992 90364 463004
rect 77260 462964 90364 462992
rect 77260 462952 77266 462964
rect 90358 462952 90364 462964
rect 90416 462952 90422 463004
rect 92382 462408 92388 462460
rect 92440 462448 92446 462460
rect 225598 462448 225604 462460
rect 92440 462420 225604 462448
rect 92440 462408 92446 462420
rect 225598 462408 225604 462420
rect 225656 462408 225662 462460
rect 3510 462340 3516 462392
rect 3568 462380 3574 462392
rect 32398 462380 32404 462392
rect 3568 462352 32404 462380
rect 3568 462340 3574 462352
rect 32398 462340 32404 462352
rect 32456 462340 32462 462392
rect 223574 462340 223580 462392
rect 223632 462380 223638 462392
rect 291194 462380 291200 462392
rect 223632 462352 291200 462380
rect 223632 462340 223638 462352
rect 291194 462340 291200 462352
rect 291252 462340 291258 462392
rect 80054 461592 80060 461644
rect 80112 461632 80118 461644
rect 113266 461632 113272 461644
rect 80112 461604 113272 461632
rect 80112 461592 80118 461604
rect 113266 461592 113272 461604
rect 113324 461592 113330 461644
rect 285674 461592 285680 461644
rect 285732 461632 285738 461644
rect 583202 461632 583208 461644
rect 285732 461604 583208 461632
rect 285732 461592 285738 461604
rect 583202 461592 583208 461604
rect 583260 461592 583266 461644
rect 166902 460980 166908 461032
rect 166960 461020 166966 461032
rect 233234 461020 233240 461032
rect 166960 460992 233240 461020
rect 166960 460980 166966 460992
rect 233234 460980 233240 460992
rect 233292 460980 233298 461032
rect 75178 460912 75184 460964
rect 75236 460952 75242 460964
rect 75822 460952 75828 460964
rect 75236 460924 75828 460952
rect 75236 460912 75242 460924
rect 75822 460912 75828 460924
rect 75880 460952 75886 460964
rect 195974 460952 195980 460964
rect 75880 460924 195980 460952
rect 75880 460912 75886 460924
rect 195974 460912 195980 460924
rect 196032 460912 196038 460964
rect 202138 460912 202144 460964
rect 202196 460952 202202 460964
rect 285674 460952 285680 460964
rect 202196 460924 285680 460952
rect 202196 460912 202202 460924
rect 285674 460912 285680 460924
rect 285732 460912 285738 460964
rect 184842 459620 184848 459672
rect 184900 459660 184906 459672
rect 233326 459660 233332 459672
rect 184900 459632 233332 459660
rect 184900 459620 184906 459632
rect 233326 459620 233332 459632
rect 233384 459620 233390 459672
rect 119338 459552 119344 459604
rect 119396 459592 119402 459604
rect 258258 459592 258264 459604
rect 119396 459564 258264 459592
rect 119396 459552 119402 459564
rect 258258 459552 258264 459564
rect 258316 459552 258322 459604
rect 95234 458260 95240 458312
rect 95292 458300 95298 458312
rect 197078 458300 197084 458312
rect 95292 458272 197084 458300
rect 95292 458260 95298 458272
rect 197078 458260 197084 458272
rect 197136 458300 197142 458312
rect 227714 458300 227720 458312
rect 197136 458272 227720 458300
rect 197136 458260 197142 458272
rect 227714 458260 227720 458272
rect 227772 458260 227778 458312
rect 85482 458192 85488 458244
rect 85540 458232 85546 458244
rect 86218 458232 86224 458244
rect 85540 458204 86224 458232
rect 85540 458192 85546 458204
rect 86218 458192 86224 458204
rect 86276 458192 86282 458244
rect 148318 458192 148324 458244
rect 148376 458232 148382 458244
rect 256786 458232 256792 458244
rect 148376 458204 256792 458232
rect 148376 458192 148382 458204
rect 256786 458192 256792 458204
rect 256844 458192 256850 458244
rect 192478 456900 192484 456952
rect 192536 456940 192542 456952
rect 218882 456940 218888 456952
rect 192536 456912 218888 456940
rect 192536 456900 192542 456912
rect 218882 456900 218888 456912
rect 218940 456900 218946 456952
rect 72418 456832 72424 456884
rect 72476 456872 72482 456884
rect 157334 456872 157340 456884
rect 72476 456844 157340 456872
rect 72476 456832 72482 456844
rect 157334 456832 157340 456844
rect 157392 456872 157398 456884
rect 197354 456872 197360 456884
rect 157392 456844 197360 456872
rect 157392 456832 157398 456844
rect 197354 456832 197360 456844
rect 197412 456832 197418 456884
rect 226426 456832 226432 456884
rect 226484 456872 226490 456884
rect 260834 456872 260840 456884
rect 226484 456844 260840 456872
rect 226484 456832 226490 456844
rect 260834 456832 260840 456844
rect 260892 456832 260898 456884
rect 78674 456764 78680 456816
rect 78732 456804 78738 456816
rect 175182 456804 175188 456816
rect 78732 456776 175188 456804
rect 78732 456764 78738 456776
rect 175182 456764 175188 456776
rect 175240 456764 175246 456816
rect 204438 456764 204444 456816
rect 204496 456804 204502 456816
rect 247402 456804 247408 456816
rect 204496 456776 247408 456804
rect 204496 456764 204502 456776
rect 247402 456764 247408 456776
rect 247460 456764 247466 456816
rect 288342 456764 288348 456816
rect 288400 456804 288406 456816
rect 580166 456804 580172 456816
rect 288400 456776 580172 456804
rect 288400 456764 288406 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 68922 456016 68928 456068
rect 68980 456056 68986 456068
rect 80054 456056 80060 456068
rect 68980 456028 80060 456056
rect 68980 456016 68986 456028
rect 80054 456016 80060 456028
rect 80112 456016 80118 456068
rect 190362 455472 190368 455524
rect 190420 455512 190426 455524
rect 204530 455512 204536 455524
rect 190420 455484 204536 455512
rect 190420 455472 190426 455484
rect 204530 455472 204536 455484
rect 204588 455472 204594 455524
rect 235994 455472 236000 455524
rect 236052 455512 236058 455524
rect 260098 455512 260104 455524
rect 236052 455484 260104 455512
rect 236052 455472 236058 455484
rect 260098 455472 260104 455484
rect 260156 455472 260162 455524
rect 192570 455404 192576 455456
rect 192628 455444 192634 455456
rect 213178 455444 213184 455456
rect 192628 455416 213184 455444
rect 192628 455404 192634 455416
rect 213178 455404 213184 455416
rect 213236 455404 213242 455456
rect 237374 455404 237380 455456
rect 237432 455444 237438 455456
rect 273346 455444 273352 455456
rect 237432 455416 273352 455444
rect 237432 455404 237438 455416
rect 273346 455404 273352 455416
rect 273404 455404 273410 455456
rect 74534 455336 74540 455388
rect 74592 455376 74598 455388
rect 75362 455376 75368 455388
rect 74592 455348 75368 455376
rect 74592 455336 74598 455348
rect 75362 455336 75368 455348
rect 75420 455336 75426 455388
rect 88242 454656 88248 454708
rect 88300 454696 88306 454708
rect 104894 454696 104900 454708
rect 88300 454668 104900 454696
rect 88300 454656 88306 454668
rect 104894 454656 104900 454668
rect 104952 454656 104958 454708
rect 75362 454112 75368 454164
rect 75420 454152 75426 454164
rect 151078 454152 151084 454164
rect 75420 454124 151084 454152
rect 75420 454112 75426 454124
rect 151078 454112 151084 454124
rect 151136 454112 151142 454164
rect 193398 454112 193404 454164
rect 193456 454152 193462 454164
rect 237834 454152 237840 454164
rect 193456 454124 237840 454152
rect 193456 454112 193462 454124
rect 237834 454112 237840 454124
rect 237892 454112 237898 454164
rect 240778 454112 240784 454164
rect 240836 454152 240842 454164
rect 276014 454152 276020 454164
rect 240836 454124 276020 454152
rect 240836 454112 240842 454124
rect 276014 454112 276020 454124
rect 276072 454112 276078 454164
rect 116670 454044 116676 454096
rect 116728 454084 116734 454096
rect 245746 454084 245752 454096
rect 116728 454056 245752 454084
rect 116728 454044 116734 454056
rect 245746 454044 245752 454056
rect 245804 454044 245810 454096
rect 239214 453976 239220 454028
rect 239272 454016 239278 454028
rect 240778 454016 240784 454028
rect 239272 453988 240784 454016
rect 239272 453976 239278 453988
rect 240778 453976 240784 453988
rect 240836 453976 240842 454028
rect 240134 453432 240140 453484
rect 240192 453472 240198 453484
rect 240870 453472 240876 453484
rect 240192 453444 240876 453472
rect 240192 453432 240198 453444
rect 240870 453432 240876 453444
rect 240928 453432 240934 453484
rect 231670 453364 231676 453416
rect 231728 453404 231734 453416
rect 237374 453404 237380 453416
rect 231728 453376 237380 453404
rect 231728 453364 231734 453376
rect 237374 453364 237380 453376
rect 237432 453364 237438 453416
rect 232590 452752 232596 452804
rect 232648 452792 232654 452804
rect 232648 452764 238754 452792
rect 232648 452752 232654 452764
rect 82814 452684 82820 452736
rect 82872 452724 82878 452736
rect 168282 452724 168288 452736
rect 82872 452696 168288 452724
rect 82872 452684 82878 452696
rect 168282 452684 168288 452696
rect 168340 452724 168346 452736
rect 200390 452724 200396 452736
rect 168340 452696 200396 452724
rect 168340 452684 168346 452696
rect 200390 452684 200396 452696
rect 200448 452684 200454 452736
rect 201586 452684 201592 452736
rect 201644 452724 201650 452736
rect 205910 452724 205916 452736
rect 201644 452696 205916 452724
rect 201644 452684 201650 452696
rect 205910 452684 205916 452696
rect 205968 452684 205974 452736
rect 75270 452616 75276 452668
rect 75328 452656 75334 452668
rect 201310 452656 201316 452668
rect 75328 452628 201316 452656
rect 75328 452616 75334 452628
rect 201310 452616 201316 452628
rect 201368 452616 201374 452668
rect 202782 452616 202788 452668
rect 202840 452656 202846 452668
rect 209774 452656 209780 452668
rect 202840 452628 209780 452656
rect 202840 452616 202846 452628
rect 209774 452616 209780 452628
rect 209832 452616 209838 452668
rect 227714 452616 227720 452668
rect 227772 452656 227778 452668
rect 229646 452656 229652 452668
rect 227772 452628 229652 452656
rect 227772 452616 227778 452628
rect 229646 452616 229652 452628
rect 229704 452616 229710 452668
rect 238726 452656 238754 452764
rect 240134 452684 240140 452736
rect 240192 452724 240198 452736
rect 259454 452724 259460 452736
rect 240192 452696 259460 452724
rect 240192 452684 240198 452696
rect 259454 452684 259460 452696
rect 259512 452684 259518 452736
rect 269114 452656 269120 452668
rect 238726 452628 269120 452656
rect 269114 452616 269120 452628
rect 269172 452616 269178 452668
rect 111794 452548 111800 452600
rect 111852 452588 111858 452600
rect 112438 452588 112444 452600
rect 111852 452560 112444 452588
rect 111852 452548 111858 452560
rect 112438 452548 112444 452560
rect 112496 452548 112502 452600
rect 191098 451868 191104 451920
rect 191156 451908 191162 451920
rect 202782 451908 202788 451920
rect 191156 451880 202788 451908
rect 191156 451868 191162 451880
rect 202782 451868 202788 451880
rect 202840 451868 202846 451920
rect 104250 451324 104256 451376
rect 104308 451364 104314 451376
rect 137278 451364 137284 451376
rect 104308 451336 137284 451364
rect 104308 451324 104314 451336
rect 137278 451324 137284 451336
rect 137336 451324 137342 451376
rect 248782 451324 248788 451376
rect 248840 451364 248846 451376
rect 254026 451364 254032 451376
rect 248840 451336 254032 451364
rect 248840 451324 248846 451336
rect 254026 451324 254032 451336
rect 254084 451324 254090 451376
rect 39298 451256 39304 451308
rect 39356 451296 39362 451308
rect 111794 451296 111800 451308
rect 39356 451268 111800 451296
rect 39356 451256 39362 451268
rect 111794 451256 111800 451268
rect 111852 451256 111858 451308
rect 122098 451256 122104 451308
rect 122156 451296 122162 451308
rect 142062 451296 142068 451308
rect 122156 451268 142068 451296
rect 122156 451256 122162 451268
rect 142062 451256 142068 451268
rect 142120 451256 142126 451308
rect 184382 451256 184388 451308
rect 184440 451296 184446 451308
rect 199286 451296 199292 451308
rect 184440 451268 199292 451296
rect 184440 451256 184446 451268
rect 199286 451256 199292 451268
rect 199344 451256 199350 451308
rect 204070 451256 204076 451308
rect 204128 451296 204134 451308
rect 277394 451296 277400 451308
rect 204128 451268 277400 451296
rect 204128 451256 204134 451268
rect 277394 451256 277400 451268
rect 277452 451256 277458 451308
rect 87598 449964 87604 450016
rect 87656 450004 87662 450016
rect 214190 450004 214196 450016
rect 87656 449976 214196 450004
rect 87656 449964 87662 449976
rect 214190 449964 214196 449976
rect 214248 449964 214254 450016
rect 218606 449964 218612 450016
rect 218664 450004 218670 450016
rect 270494 450004 270500 450016
rect 218664 449976 270500 450004
rect 218664 449964 218670 449976
rect 270494 449964 270500 449976
rect 270552 449964 270558 450016
rect 67266 449896 67272 449948
rect 67324 449936 67330 449948
rect 94774 449936 94780 449948
rect 67324 449908 94780 449936
rect 67324 449896 67330 449908
rect 94774 449896 94780 449908
rect 94832 449936 94838 449948
rect 95142 449936 95148 449948
rect 94832 449908 95148 449936
rect 94832 449896 94838 449908
rect 95142 449896 95148 449908
rect 95200 449896 95206 449948
rect 98638 449896 98644 449948
rect 98696 449936 98702 449948
rect 232222 449936 232228 449948
rect 98696 449908 232228 449936
rect 98696 449896 98702 449908
rect 232222 449896 232228 449908
rect 232280 449896 232286 449948
rect 233142 449896 233148 449948
rect 233200 449936 233206 449948
rect 244550 449936 244556 449948
rect 233200 449908 244556 449936
rect 233200 449896 233206 449908
rect 244550 449896 244556 449908
rect 244608 449936 244614 449948
rect 262858 449936 262864 449948
rect 244608 449908 262864 449936
rect 244608 449896 244614 449908
rect 262858 449896 262864 449908
rect 262916 449896 262922 449948
rect 191466 449828 191472 449880
rect 191524 449868 191530 449880
rect 246022 449868 246028 449880
rect 191524 449840 246028 449868
rect 191524 449828 191530 449840
rect 246022 449828 246028 449840
rect 246080 449828 246086 449880
rect 251818 449692 251824 449744
rect 251876 449732 251882 449744
rect 251876 449704 258074 449732
rect 251876 449692 251882 449704
rect 41322 449148 41328 449200
rect 41380 449188 41386 449200
rect 106918 449188 106924 449200
rect 41380 449160 106924 449188
rect 41380 449148 41386 449160
rect 106918 449148 106924 449160
rect 106976 449148 106982 449200
rect 185578 449148 185584 449200
rect 185636 449188 185642 449200
rect 193398 449188 193404 449200
rect 185636 449160 193404 449188
rect 185636 449148 185642 449160
rect 193398 449148 193404 449160
rect 193456 449148 193462 449200
rect 258046 448984 258074 449704
rect 281626 448984 281632 448996
rect 258046 448956 281632 448984
rect 281626 448944 281632 448956
rect 281684 448944 281690 448996
rect 3142 448536 3148 448588
rect 3200 448576 3206 448588
rect 11698 448576 11704 448588
rect 3200 448548 11704 448576
rect 3200 448536 3206 448548
rect 11698 448536 11704 448548
rect 11756 448536 11762 448588
rect 61930 448536 61936 448588
rect 61988 448576 61994 448588
rect 169018 448576 169024 448588
rect 61988 448548 169024 448576
rect 61988 448536 61994 448548
rect 169018 448536 169024 448548
rect 169076 448536 169082 448588
rect 176562 448536 176568 448588
rect 176620 448576 176626 448588
rect 191650 448576 191656 448588
rect 176620 448548 191656 448576
rect 176620 448536 176626 448548
rect 191650 448536 191656 448548
rect 191708 448536 191714 448588
rect 67634 448332 67640 448384
rect 67692 448372 67698 448384
rect 75362 448372 75368 448384
rect 67692 448344 75368 448372
rect 67692 448332 67698 448344
rect 75362 448332 75368 448344
rect 75420 448332 75426 448384
rect 73246 447788 73252 447840
rect 73304 447828 73310 447840
rect 82814 447828 82820 447840
rect 73304 447800 82820 447828
rect 73304 447788 73310 447800
rect 82814 447788 82820 447800
rect 82872 447788 82878 447840
rect 95142 447788 95148 447840
rect 95200 447828 95206 447840
rect 170398 447828 170404 447840
rect 95200 447800 170404 447828
rect 95200 447788 95206 447800
rect 170398 447788 170404 447800
rect 170456 447788 170462 447840
rect 178954 447788 178960 447840
rect 179012 447828 179018 447840
rect 192570 447828 192576 447840
rect 179012 447800 192576 447828
rect 179012 447788 179018 447800
rect 192570 447788 192576 447800
rect 192628 447788 192634 447840
rect 82906 447108 82912 447160
rect 82964 447148 82970 447160
rect 83458 447148 83464 447160
rect 82964 447120 83464 447148
rect 82964 447108 82970 447120
rect 83458 447108 83464 447120
rect 83516 447148 83522 447160
rect 178954 447148 178960 447160
rect 83516 447120 178960 447148
rect 83516 447108 83522 447120
rect 178954 447108 178960 447120
rect 179012 447148 179018 447160
rect 179230 447148 179236 447160
rect 179012 447120 179236 447148
rect 179012 447108 179018 447120
rect 179230 447108 179236 447120
rect 179288 447108 179294 447160
rect 172422 446360 172428 446412
rect 172480 446400 172486 446412
rect 192478 446400 192484 446412
rect 172480 446372 192484 446400
rect 172480 446360 172486 446372
rect 192478 446360 192484 446372
rect 192536 446360 192542 446412
rect 253842 446360 253848 446412
rect 253900 446400 253906 446412
rect 267734 446400 267740 446412
rect 253900 446372 267740 446400
rect 253900 446360 253906 446372
rect 267734 446360 267740 446372
rect 267792 446360 267798 446412
rect 37090 445816 37096 445868
rect 37148 445856 37154 445868
rect 77294 445856 77300 445868
rect 37148 445828 77300 445856
rect 37148 445816 37154 445828
rect 77294 445816 77300 445828
rect 77352 445856 77358 445868
rect 77938 445856 77944 445868
rect 77352 445828 77944 445856
rect 77352 445816 77358 445828
rect 77938 445816 77944 445828
rect 77996 445816 78002 445868
rect 66162 445748 66168 445800
rect 66220 445788 66226 445800
rect 191742 445788 191748 445800
rect 66220 445760 191748 445788
rect 66220 445748 66226 445760
rect 191742 445748 191748 445760
rect 191800 445748 191806 445800
rect 50982 445680 50988 445732
rect 51040 445720 51046 445732
rect 95142 445720 95148 445732
rect 51040 445692 95148 445720
rect 51040 445680 51046 445692
rect 95142 445680 95148 445692
rect 95200 445680 95206 445732
rect 83458 444388 83464 444440
rect 83516 444428 83522 444440
rect 176654 444428 176660 444440
rect 83516 444400 176660 444428
rect 83516 444388 83522 444400
rect 176654 444388 176660 444400
rect 176712 444428 176718 444440
rect 191742 444428 191748 444440
rect 176712 444400 191748 444428
rect 176712 444388 176718 444400
rect 191742 444388 191748 444400
rect 191800 444388 191806 444440
rect 188430 444320 188436 444372
rect 188488 444360 188494 444372
rect 190454 444360 190460 444372
rect 188488 444332 190460 444360
rect 188488 444320 188494 444332
rect 190454 444320 190460 444332
rect 190512 444320 190518 444372
rect 69106 443640 69112 443692
rect 69164 443680 69170 443692
rect 166258 443680 166264 443692
rect 69164 443652 166264 443680
rect 69164 443640 69170 443652
rect 166258 443640 166264 443652
rect 166316 443640 166322 443692
rect 255682 443640 255688 443692
rect 255740 443680 255746 443692
rect 284294 443680 284300 443692
rect 255740 443652 284300 443680
rect 255740 443640 255746 443652
rect 284294 443640 284300 443652
rect 284352 443640 284358 443692
rect 33778 442960 33784 443012
rect 33836 443000 33842 443012
rect 95326 443000 95332 443012
rect 33836 442972 95332 443000
rect 33836 442960 33842 442972
rect 95326 442960 95332 442972
rect 95384 442960 95390 443012
rect 255406 442960 255412 443012
rect 255464 443000 255470 443012
rect 258810 443000 258816 443012
rect 255464 442972 258816 443000
rect 255464 442960 255470 442972
rect 258810 442960 258816 442972
rect 258868 442960 258874 443012
rect 88426 442892 88432 442944
rect 88484 442932 88490 442944
rect 92566 442932 92572 442944
rect 88484 442904 92572 442932
rect 88484 442892 88490 442904
rect 92566 442892 92572 442904
rect 92624 442892 92630 442944
rect 48130 442212 48136 442264
rect 48188 442252 48194 442264
rect 52362 442252 52368 442264
rect 48188 442224 52368 442252
rect 48188 442212 48194 442224
rect 52362 442212 52368 442224
rect 52420 442252 52426 442264
rect 88426 442252 88432 442264
rect 52420 442224 88432 442252
rect 52420 442212 52426 442224
rect 88426 442212 88432 442224
rect 88484 442212 88490 442264
rect 254670 442212 254676 442264
rect 254728 442252 254734 442264
rect 271874 442252 271880 442264
rect 254728 442224 271880 442252
rect 254728 442212 254734 442224
rect 271874 442212 271880 442224
rect 271932 442212 271938 442264
rect 67450 441600 67456 441652
rect 67508 441640 67514 441652
rect 162118 441640 162124 441652
rect 67508 441612 162124 441640
rect 67508 441600 67514 441612
rect 162118 441600 162124 441612
rect 162176 441600 162182 441652
rect 7558 441532 7564 441584
rect 7616 441572 7622 441584
rect 104158 441572 104164 441584
rect 7616 441544 104164 441572
rect 7616 441532 7622 441544
rect 104158 441532 104164 441544
rect 104216 441532 104222 441584
rect 161382 440852 161388 440904
rect 161440 440892 161446 440904
rect 191282 440892 191288 440904
rect 161440 440864 191288 440892
rect 161440 440852 161446 440864
rect 191282 440852 191288 440864
rect 191340 440852 191346 440904
rect 63310 440240 63316 440292
rect 63368 440280 63374 440292
rect 191190 440280 191196 440292
rect 63368 440252 191196 440280
rect 63368 440240 63374 440252
rect 191190 440240 191196 440252
rect 191248 440240 191254 440292
rect 67174 439492 67180 439544
rect 67232 439532 67238 439544
rect 83458 439532 83464 439544
rect 67232 439504 83464 439532
rect 67232 439492 67238 439504
rect 83458 439492 83464 439504
rect 83516 439492 83522 439544
rect 104802 439492 104808 439544
rect 104860 439532 104866 439544
rect 114646 439532 114652 439544
rect 104860 439504 114652 439532
rect 104860 439492 104866 439504
rect 114646 439492 114652 439504
rect 114704 439492 114710 439544
rect 255406 439492 255412 439544
rect 255464 439532 255470 439544
rect 258258 439532 258264 439544
rect 255464 439504 258264 439532
rect 255464 439492 255470 439504
rect 258258 439492 258264 439504
rect 258316 439532 258322 439544
rect 288618 439532 288624 439544
rect 258316 439504 288624 439532
rect 258316 439492 258322 439504
rect 288618 439492 288624 439504
rect 288676 439532 288682 439544
rect 582926 439532 582932 439544
rect 288676 439504 582932 439532
rect 288676 439492 288682 439504
rect 582926 439492 582932 439504
rect 582984 439492 582990 439544
rect 73982 438880 73988 438932
rect 74040 438920 74046 438932
rect 75270 438920 75276 438932
rect 74040 438892 75276 438920
rect 74040 438880 74046 438892
rect 75270 438880 75276 438892
rect 75328 438880 75334 438932
rect 82906 438880 82912 438932
rect 82964 438920 82970 438932
rect 180058 438920 180064 438932
rect 82964 438892 180064 438920
rect 82964 438880 82970 438892
rect 180058 438880 180064 438892
rect 180116 438880 180122 438932
rect 48038 438812 48044 438864
rect 48096 438852 48102 438864
rect 74718 438852 74724 438864
rect 48096 438824 74724 438852
rect 48096 438812 48102 438824
rect 74718 438812 74724 438824
rect 74776 438852 74782 438864
rect 75362 438852 75368 438864
rect 74776 438824 75368 438852
rect 74776 438812 74782 438824
rect 75362 438812 75368 438824
rect 75420 438812 75426 438864
rect 94498 438812 94504 438864
rect 94556 438852 94562 438864
rect 97350 438852 97356 438864
rect 94556 438824 97356 438852
rect 94556 438812 94562 438824
rect 97350 438812 97356 438824
rect 97408 438812 97414 438864
rect 255498 438812 255504 438864
rect 255556 438852 255562 438864
rect 262214 438852 262220 438864
rect 255556 438824 262220 438852
rect 255556 438812 255562 438824
rect 262214 438812 262220 438824
rect 262272 438812 262278 438864
rect 70486 437452 70492 437504
rect 70544 437492 70550 437504
rect 191742 437492 191748 437504
rect 70544 437464 191748 437492
rect 70544 437452 70550 437464
rect 191742 437452 191748 437464
rect 191800 437452 191806 437504
rect 262214 437452 262220 437504
rect 262272 437492 262278 437504
rect 263686 437492 263692 437504
rect 262272 437464 263692 437492
rect 262272 437452 262278 437464
rect 263686 437452 263692 437464
rect 263744 437452 263750 437504
rect 82814 437384 82820 437436
rect 82872 437424 82878 437436
rect 83918 437424 83924 437436
rect 82872 437396 83924 437424
rect 82872 437384 82878 437396
rect 83918 437384 83924 437396
rect 83976 437424 83982 437436
rect 87598 437424 87604 437436
rect 83976 437396 87604 437424
rect 83976 437384 83982 437396
rect 87598 437384 87604 437396
rect 87656 437384 87662 437436
rect 97350 437384 97356 437436
rect 97408 437424 97414 437436
rect 98638 437424 98644 437436
rect 97408 437396 98644 437424
rect 97408 437384 97414 437396
rect 98638 437384 98644 437396
rect 98696 437384 98702 437436
rect 98730 437384 98736 437436
rect 98788 437424 98794 437436
rect 103698 437424 103704 437436
rect 98788 437396 103704 437424
rect 98788 437384 98794 437396
rect 103698 437384 103704 437396
rect 103756 437424 103762 437436
rect 104250 437424 104256 437436
rect 103756 437396 104256 437424
rect 103756 437384 103762 437396
rect 104250 437384 104256 437396
rect 104308 437384 104314 437436
rect 108298 437384 108304 437436
rect 108356 437424 108362 437436
rect 122098 437424 122104 437436
rect 108356 437396 122104 437424
rect 108356 437384 108362 437396
rect 122098 437384 122104 437396
rect 122156 437384 122162 437436
rect 255498 437384 255504 437436
rect 255556 437424 255562 437436
rect 582374 437424 582380 437436
rect 255556 437396 582380 437424
rect 255556 437384 255562 437396
rect 582374 437384 582380 437396
rect 582432 437384 582438 437436
rect 107378 436704 107384 436756
rect 107436 436744 107442 436756
rect 116670 436744 116676 436756
rect 107436 436716 116676 436744
rect 107436 436704 107442 436716
rect 116670 436704 116676 436716
rect 116728 436704 116734 436756
rect 87322 436432 87328 436484
rect 87380 436472 87386 436484
rect 90450 436472 90456 436484
rect 87380 436444 90456 436472
rect 87380 436432 87386 436444
rect 90450 436432 90456 436444
rect 90508 436432 90514 436484
rect 53742 436160 53748 436212
rect 53800 436200 53806 436212
rect 69842 436200 69848 436212
rect 53800 436172 69848 436200
rect 53800 436160 53806 436172
rect 69842 436160 69848 436172
rect 69900 436160 69906 436212
rect 70854 436200 70860 436212
rect 70366 436172 70860 436200
rect 17218 436092 17224 436144
rect 17276 436132 17282 436144
rect 70366 436132 70394 436172
rect 70854 436160 70860 436172
rect 70912 436200 70918 436212
rect 75178 436200 75184 436212
rect 70912 436172 75184 436200
rect 70912 436160 70918 436172
rect 75178 436160 75184 436172
rect 75236 436160 75242 436212
rect 75638 436160 75644 436212
rect 75696 436200 75702 436212
rect 78030 436200 78036 436212
rect 75696 436172 78036 436200
rect 75696 436160 75702 436172
rect 78030 436160 78036 436172
rect 78088 436160 78094 436212
rect 17276 436104 70394 436132
rect 17276 436092 17282 436104
rect 71682 436092 71688 436144
rect 71740 436132 71746 436144
rect 72418 436132 72424 436144
rect 71740 436104 72424 436132
rect 71740 436092 71746 436104
rect 72418 436092 72424 436104
rect 72476 436092 72482 436144
rect 72510 436092 72516 436144
rect 72568 436132 72574 436144
rect 77478 436132 77484 436144
rect 72568 436104 77484 436132
rect 72568 436092 72574 436104
rect 77478 436092 77484 436104
rect 77536 436092 77542 436144
rect 92382 436092 92388 436144
rect 92440 436132 92446 436144
rect 94222 436132 94228 436144
rect 92440 436104 94228 436132
rect 92440 436092 92446 436104
rect 94222 436092 94228 436104
rect 94280 436092 94286 436144
rect 107562 435412 107568 435464
rect 107620 435452 107626 435464
rect 116026 435452 116032 435464
rect 107620 435424 116032 435452
rect 107620 435412 107626 435424
rect 116026 435412 116032 435424
rect 116084 435412 116090 435464
rect 55030 435344 55036 435396
rect 55088 435384 55094 435396
rect 191742 435384 191748 435396
rect 55088 435356 191748 435384
rect 55088 435344 55094 435356
rect 191742 435344 191748 435356
rect 191800 435344 191806 435396
rect 255406 435344 255412 435396
rect 255464 435384 255470 435396
rect 259546 435384 259552 435396
rect 255464 435356 259552 435384
rect 255464 435344 255470 435356
rect 259546 435344 259552 435356
rect 259604 435384 259610 435396
rect 274634 435384 274640 435396
rect 259604 435356 274640 435384
rect 259604 435344 259610 435356
rect 274634 435344 274640 435356
rect 274692 435344 274698 435396
rect 137370 434868 137376 434920
rect 137428 434908 137434 434920
rect 141418 434908 141424 434920
rect 137428 434880 141424 434908
rect 137428 434868 137434 434880
rect 141418 434868 141424 434880
rect 141476 434868 141482 434920
rect 64690 434732 64696 434784
rect 64748 434772 64754 434784
rect 73982 434772 73988 434784
rect 64748 434744 73988 434772
rect 64748 434732 64754 434744
rect 73982 434732 73988 434744
rect 74040 434732 74046 434784
rect 115014 434664 115020 434716
rect 115072 434704 115078 434716
rect 178678 434704 178684 434716
rect 115072 434676 178684 434704
rect 115072 434664 115078 434676
rect 178678 434664 178684 434676
rect 178736 434664 178742 434716
rect 188430 434664 188436 434716
rect 188488 434704 188494 434716
rect 188890 434704 188896 434716
rect 188488 434676 188896 434704
rect 188488 434664 188494 434676
rect 188890 434664 188896 434676
rect 188948 434704 188954 434716
rect 191742 434704 191748 434716
rect 188948 434676 191748 434704
rect 188948 434664 188954 434676
rect 191742 434664 191748 434676
rect 191800 434664 191806 434716
rect 255406 434596 255412 434648
rect 255464 434636 255470 434648
rect 258074 434636 258080 434648
rect 255464 434608 258080 434636
rect 255464 434596 255470 434608
rect 258074 434596 258080 434608
rect 258132 434636 258138 434648
rect 265066 434636 265072 434648
rect 258132 434608 265072 434636
rect 258132 434596 258138 434608
rect 265066 434596 265072 434608
rect 265124 434596 265130 434648
rect 100202 433984 100208 434036
rect 100260 434024 100266 434036
rect 115382 434024 115388 434036
rect 100260 433996 115388 434024
rect 100260 433984 100266 433996
rect 115382 433984 115388 433996
rect 115440 433984 115446 434036
rect 96586 433724 106274 433752
rect 64782 433304 64788 433356
rect 64840 433344 64846 433356
rect 96586 433344 96614 433724
rect 64840 433316 96614 433344
rect 106246 433344 106274 433724
rect 191650 433344 191656 433356
rect 106246 433316 191656 433344
rect 64840 433304 64846 433316
rect 191650 433304 191656 433316
rect 191708 433304 191714 433356
rect 68646 433236 68652 433288
rect 68704 433276 68710 433288
rect 188890 433276 188896 433288
rect 68704 433248 80054 433276
rect 68704 433236 68710 433248
rect 80026 433140 80054 433248
rect 102520 433248 103514 433276
rect 102520 433140 102548 433248
rect 103486 433208 103514 433248
rect 113146 433248 188896 433276
rect 113146 433208 113174 433248
rect 188890 433236 188896 433248
rect 188948 433236 188954 433288
rect 103486 433180 113174 433208
rect 80026 433112 102548 433140
rect 255958 432624 255964 432676
rect 256016 432664 256022 432676
rect 262214 432664 262220 432676
rect 256016 432636 262220 432664
rect 256016 432624 256022 432636
rect 262214 432624 262220 432636
rect 262272 432624 262278 432676
rect 254578 432556 254584 432608
rect 254636 432596 254642 432608
rect 283006 432596 283012 432608
rect 254636 432568 283012 432596
rect 254636 432556 254642 432568
rect 283006 432556 283012 432568
rect 283064 432556 283070 432608
rect 187418 431944 187424 431996
rect 187476 431984 187482 431996
rect 191098 431984 191104 431996
rect 187476 431956 191104 431984
rect 187476 431944 187482 431956
rect 191098 431944 191104 431956
rect 191156 431944 191162 431996
rect 115290 431264 115296 431316
rect 115348 431304 115354 431316
rect 118694 431304 118700 431316
rect 115348 431276 118700 431304
rect 115348 431264 115354 431276
rect 118694 431264 118700 431276
rect 118752 431264 118758 431316
rect 171042 431196 171048 431248
rect 171100 431236 171106 431248
rect 180150 431236 180156 431248
rect 171100 431208 180156 431236
rect 171100 431196 171106 431208
rect 180150 431196 180156 431208
rect 180208 431196 180214 431248
rect 115842 430244 115848 430296
rect 115900 430284 115906 430296
rect 119430 430284 119436 430296
rect 115900 430256 119436 430284
rect 115900 430244 115906 430256
rect 119430 430244 119436 430256
rect 119488 430244 119494 430296
rect 255130 429836 255136 429888
rect 255188 429876 255194 429888
rect 258718 429876 258724 429888
rect 255188 429848 258724 429876
rect 255188 429836 255194 429848
rect 258718 429836 258724 429848
rect 258776 429836 258782 429888
rect 258810 429836 258816 429888
rect 258868 429876 258874 429888
rect 270586 429876 270592 429888
rect 258868 429848 270592 429876
rect 258868 429836 258874 429848
rect 270586 429836 270592 429848
rect 270644 429836 270650 429888
rect 61930 429088 61936 429140
rect 61988 429128 61994 429140
rect 66806 429128 66812 429140
rect 61988 429100 66812 429128
rect 61988 429088 61994 429100
rect 66806 429088 66812 429100
rect 66864 429088 66870 429140
rect 151078 429088 151084 429140
rect 151136 429128 151142 429140
rect 191558 429128 191564 429140
rect 151136 429100 191564 429128
rect 151136 429088 151142 429100
rect 191558 429088 191564 429100
rect 191616 429088 191622 429140
rect 115842 428408 115848 428460
rect 115900 428448 115906 428460
rect 122926 428448 122932 428460
rect 115900 428420 122932 428448
rect 115900 428408 115906 428420
rect 122926 428408 122932 428420
rect 122984 428448 122990 428460
rect 123478 428448 123484 428460
rect 122984 428420 123484 428448
rect 122984 428408 122990 428420
rect 123478 428408 123484 428420
rect 123536 428408 123542 428460
rect 46842 427796 46848 427848
rect 46900 427836 46906 427848
rect 66254 427836 66260 427848
rect 46900 427808 66260 427836
rect 46900 427796 46906 427808
rect 66254 427796 66260 427808
rect 66312 427796 66318 427848
rect 255406 427796 255412 427848
rect 255464 427836 255470 427848
rect 264974 427836 264980 427848
rect 255464 427808 264980 427836
rect 255464 427796 255470 427808
rect 264974 427796 264980 427808
rect 265032 427796 265038 427848
rect 115842 427728 115848 427780
rect 115900 427768 115906 427780
rect 159358 427768 159364 427780
rect 115900 427740 159364 427768
rect 115900 427728 115906 427740
rect 159358 427728 159364 427740
rect 159416 427728 159422 427780
rect 255498 427728 255504 427780
rect 255556 427768 255562 427780
rect 260926 427768 260932 427780
rect 255556 427740 260932 427768
rect 255556 427728 255562 427740
rect 260926 427728 260932 427740
rect 260984 427768 260990 427780
rect 262122 427768 262128 427780
rect 260984 427740 262128 427768
rect 260984 427728 260990 427740
rect 262122 427728 262128 427740
rect 262180 427728 262186 427780
rect 169018 427048 169024 427100
rect 169076 427088 169082 427100
rect 176746 427088 176752 427100
rect 169076 427060 176752 427088
rect 169076 427048 169082 427060
rect 176746 427048 176752 427060
rect 176804 427048 176810 427100
rect 262122 427048 262128 427100
rect 262180 427088 262186 427100
rect 279326 427088 279332 427100
rect 262180 427060 279332 427088
rect 262180 427048 262186 427060
rect 279326 427048 279332 427060
rect 279384 427048 279390 427100
rect 50890 426436 50896 426488
rect 50948 426476 50954 426488
rect 66898 426476 66904 426488
rect 50948 426448 66904 426476
rect 50948 426436 50954 426448
rect 66898 426436 66904 426448
rect 66956 426436 66962 426488
rect 176746 426436 176752 426488
rect 176804 426476 176810 426488
rect 177850 426476 177856 426488
rect 176804 426448 177856 426476
rect 176804 426436 176810 426448
rect 177850 426436 177856 426448
rect 177908 426476 177914 426488
rect 191558 426476 191564 426488
rect 177908 426448 191564 426476
rect 177908 426436 177914 426448
rect 191558 426436 191564 426448
rect 191616 426436 191622 426488
rect 279326 426436 279332 426488
rect 279384 426476 279390 426488
rect 582650 426476 582656 426488
rect 279384 426448 582656 426476
rect 279384 426436 279390 426448
rect 582650 426436 582656 426448
rect 582708 426436 582714 426488
rect 115290 426096 115296 426148
rect 115348 426136 115354 426148
rect 119338 426136 119344 426148
rect 115348 426108 119344 426136
rect 115348 426096 115354 426108
rect 119338 426096 119344 426108
rect 119396 426096 119402 426148
rect 57882 425688 57888 425740
rect 57940 425728 57946 425740
rect 66070 425728 66076 425740
rect 57940 425700 66076 425728
rect 57940 425688 57946 425700
rect 66070 425688 66076 425700
rect 66128 425728 66134 425740
rect 66622 425728 66628 425740
rect 66128 425700 66628 425728
rect 66128 425688 66134 425700
rect 66622 425688 66628 425700
rect 66680 425688 66686 425740
rect 181438 425076 181444 425128
rect 181496 425116 181502 425128
rect 191006 425116 191012 425128
rect 181496 425088 191012 425116
rect 181496 425076 181502 425088
rect 191006 425076 191012 425088
rect 191064 425076 191070 425128
rect 115290 424940 115296 424992
rect 115348 424980 115354 424992
rect 117406 424980 117412 424992
rect 115348 424952 117412 424980
rect 115348 424940 115354 424952
rect 117406 424940 117412 424952
rect 117464 424940 117470 424992
rect 157242 424328 157248 424380
rect 157300 424368 157306 424380
rect 181530 424368 181536 424380
rect 157300 424340 181536 424368
rect 157300 424328 157306 424340
rect 181530 424328 181536 424340
rect 181588 424328 181594 424380
rect 256786 424328 256792 424380
rect 256844 424368 256850 424380
rect 266354 424368 266360 424380
rect 256844 424340 266360 424368
rect 256844 424328 256850 424340
rect 266354 424328 266360 424340
rect 266412 424328 266418 424380
rect 114646 423716 114652 423768
rect 114704 423756 114710 423768
rect 116026 423756 116032 423768
rect 114704 423728 116032 423756
rect 114704 423716 114710 423728
rect 116026 423716 116032 423728
rect 116084 423716 116090 423768
rect 55030 423648 55036 423700
rect 55088 423688 55094 423700
rect 66806 423688 66812 423700
rect 55088 423660 66812 423688
rect 55088 423648 55094 423660
rect 66806 423648 66812 423660
rect 66864 423648 66870 423700
rect 3510 423580 3516 423632
rect 3568 423620 3574 423632
rect 39298 423620 39304 423632
rect 3568 423592 39304 423620
rect 3568 423580 3574 423592
rect 39298 423580 39304 423592
rect 39356 423580 39362 423632
rect 52362 423580 52368 423632
rect 52420 423620 52426 423632
rect 54938 423620 54944 423632
rect 52420 423592 54944 423620
rect 52420 423580 52426 423592
rect 54938 423580 54944 423592
rect 54996 423620 55002 423632
rect 66622 423620 66628 423632
rect 54996 423592 66628 423620
rect 54996 423580 55002 423592
rect 66622 423580 66628 423592
rect 66680 423580 66686 423632
rect 115842 423580 115848 423632
rect 115900 423620 115906 423632
rect 137370 423620 137376 423632
rect 115900 423592 137376 423620
rect 115900 423580 115906 423592
rect 137370 423580 137376 423592
rect 137428 423580 137434 423632
rect 137922 422900 137928 422952
rect 137980 422940 137986 422952
rect 148318 422940 148324 422952
rect 137980 422912 148324 422940
rect 137980 422900 137986 422912
rect 148318 422900 148324 422912
rect 148376 422900 148382 422952
rect 170398 422900 170404 422952
rect 170456 422940 170462 422952
rect 170950 422940 170956 422952
rect 170456 422912 170956 422940
rect 170456 422900 170462 422912
rect 170950 422900 170956 422912
rect 171008 422940 171014 422952
rect 190822 422940 190828 422952
rect 171008 422912 190828 422940
rect 171008 422900 171014 422912
rect 190822 422900 190828 422912
rect 190880 422900 190886 422952
rect 255498 422288 255504 422340
rect 255556 422328 255562 422340
rect 276106 422328 276112 422340
rect 255556 422300 276112 422328
rect 255556 422288 255562 422300
rect 276106 422288 276112 422300
rect 276164 422288 276170 422340
rect 64782 422220 64788 422272
rect 64840 422260 64846 422272
rect 66806 422260 66812 422272
rect 64840 422232 66812 422260
rect 64840 422220 64846 422232
rect 66806 422220 66812 422232
rect 66864 422220 66870 422272
rect 48038 421540 48044 421592
rect 48096 421580 48102 421592
rect 57698 421580 57704 421592
rect 48096 421552 57704 421580
rect 48096 421540 48102 421552
rect 57698 421540 57704 421552
rect 57756 421540 57762 421592
rect 255498 420928 255504 420980
rect 255556 420968 255562 420980
rect 280154 420968 280160 420980
rect 255556 420940 280160 420968
rect 255556 420928 255562 420940
rect 280154 420928 280160 420940
rect 280212 420928 280218 420980
rect 173158 419568 173164 419620
rect 173216 419608 173222 419620
rect 191558 419608 191564 419620
rect 173216 419580 191564 419608
rect 173216 419568 173222 419580
rect 191558 419568 191564 419580
rect 191616 419568 191622 419620
rect 63126 419500 63132 419552
rect 63184 419540 63190 419552
rect 66898 419540 66904 419552
rect 63184 419512 66904 419540
rect 63184 419500 63190 419512
rect 66898 419500 66904 419512
rect 66956 419500 66962 419552
rect 115842 419500 115848 419552
rect 115900 419540 115906 419552
rect 180150 419540 180156 419552
rect 115900 419512 180156 419540
rect 115900 419500 115906 419512
rect 180150 419500 180156 419512
rect 180208 419500 180214 419552
rect 255590 419500 255596 419552
rect 255648 419540 255654 419552
rect 266446 419540 266452 419552
rect 255648 419512 266452 419540
rect 255648 419500 255654 419512
rect 266446 419500 266452 419512
rect 266504 419500 266510 419552
rect 63310 419432 63316 419484
rect 63368 419472 63374 419484
rect 66806 419472 66812 419484
rect 63368 419444 66812 419472
rect 63368 419432 63374 419444
rect 66806 419432 66812 419444
rect 66864 419432 66870 419484
rect 286042 418752 286048 418804
rect 286100 418792 286106 418804
rect 583018 418792 583024 418804
rect 286100 418764 583024 418792
rect 286100 418752 286106 418764
rect 583018 418752 583024 418764
rect 583076 418752 583082 418804
rect 184290 418140 184296 418192
rect 184348 418180 184354 418192
rect 191558 418180 191564 418192
rect 184348 418152 191564 418180
rect 184348 418140 184354 418152
rect 191558 418140 191564 418152
rect 191616 418140 191622 418192
rect 255498 418140 255504 418192
rect 255556 418180 255562 418192
rect 285674 418180 285680 418192
rect 255556 418152 285680 418180
rect 255556 418140 255562 418152
rect 285674 418140 285680 418152
rect 285732 418180 285738 418192
rect 286042 418180 286048 418192
rect 285732 418152 286048 418180
rect 285732 418140 285738 418152
rect 286042 418140 286048 418152
rect 286100 418140 286106 418192
rect 115198 418072 115204 418124
rect 115256 418112 115262 418124
rect 188338 418112 188344 418124
rect 115256 418084 188344 418112
rect 115256 418072 115262 418084
rect 188338 418072 188344 418084
rect 188396 418072 188402 418124
rect 115842 418004 115848 418056
rect 115900 418044 115906 418056
rect 133138 418044 133144 418056
rect 115900 418016 133144 418044
rect 115900 418004 115906 418016
rect 133138 418004 133144 418016
rect 133196 418004 133202 418056
rect 263778 417460 263784 417512
rect 263836 417500 263842 417512
rect 271138 417500 271144 417512
rect 263836 417472 271144 417500
rect 263836 417460 263842 417472
rect 271138 417460 271144 417472
rect 271196 417460 271202 417512
rect 167638 417392 167644 417444
rect 167696 417432 167702 417444
rect 184382 417432 184388 417444
rect 167696 417404 184388 417432
rect 167696 417392 167702 417404
rect 184382 417392 184388 417404
rect 184440 417392 184446 417444
rect 262122 417392 262128 417444
rect 262180 417432 262186 417444
rect 583110 417432 583116 417444
rect 262180 417404 583116 417432
rect 262180 417392 262186 417404
rect 583110 417392 583116 417404
rect 583168 417392 583174 417444
rect 255590 416848 255596 416900
rect 255648 416888 255654 416900
rect 260926 416888 260932 416900
rect 255648 416860 260932 416888
rect 255648 416848 255654 416860
rect 260926 416848 260932 416860
rect 260984 416888 260990 416900
rect 262122 416888 262128 416900
rect 260984 416860 262128 416888
rect 260984 416848 260990 416860
rect 262122 416848 262128 416860
rect 262180 416848 262186 416900
rect 187694 416780 187700 416832
rect 187752 416820 187758 416832
rect 191558 416820 191564 416832
rect 187752 416792 191564 416820
rect 187752 416780 187758 416792
rect 191558 416780 191564 416792
rect 191616 416780 191622 416832
rect 255498 416780 255504 416832
rect 255556 416820 255562 416832
rect 263778 416820 263784 416832
rect 255556 416792 263784 416820
rect 255556 416780 255562 416792
rect 263778 416780 263784 416792
rect 263836 416780 263842 416832
rect 179322 416100 179328 416152
rect 179380 416140 179386 416152
rect 188982 416140 188988 416152
rect 179380 416112 188988 416140
rect 179380 416100 179386 416112
rect 188982 416100 188988 416112
rect 189040 416140 189046 416152
rect 191006 416140 191012 416152
rect 189040 416112 191012 416140
rect 189040 416100 189046 416112
rect 191006 416100 191012 416112
rect 191064 416100 191070 416152
rect 118694 416032 118700 416084
rect 118752 416072 118758 416084
rect 137922 416072 137928 416084
rect 118752 416044 137928 416072
rect 118752 416032 118758 416044
rect 137922 416032 137928 416044
rect 137980 416032 137986 416084
rect 159450 416032 159456 416084
rect 159508 416072 159514 416084
rect 187694 416072 187700 416084
rect 159508 416044 187700 416072
rect 159508 416032 159514 416044
rect 187694 416032 187700 416044
rect 187752 416032 187758 416084
rect 39942 415420 39948 415472
rect 40000 415460 40006 415472
rect 57790 415460 57796 415472
rect 40000 415432 57796 415460
rect 40000 415420 40006 415432
rect 57790 415420 57796 415432
rect 57848 415460 57854 415472
rect 66898 415460 66904 415472
rect 57848 415432 66904 415460
rect 57848 415420 57854 415432
rect 66898 415420 66904 415432
rect 66956 415420 66962 415472
rect 115842 415420 115848 415472
rect 115900 415460 115906 415472
rect 118694 415460 118700 415472
rect 115900 415432 118700 415460
rect 115900 415420 115906 415432
rect 118694 415420 118700 415432
rect 118752 415420 118758 415472
rect 130378 414672 130384 414724
rect 130436 414712 130442 414724
rect 191558 414712 191564 414724
rect 130436 414684 191564 414712
rect 130436 414672 130442 414684
rect 191558 414672 191564 414684
rect 191616 414672 191622 414724
rect 64782 413992 64788 414044
rect 64840 414032 64846 414044
rect 66714 414032 66720 414044
rect 64840 414004 66720 414032
rect 64840 413992 64846 414004
rect 66714 413992 66720 414004
rect 66772 413992 66778 414044
rect 115842 413788 115848 413840
rect 115900 413828 115906 413840
rect 117314 413828 117320 413840
rect 115900 413800 117320 413828
rect 115900 413788 115906 413800
rect 117314 413788 117320 413800
rect 117372 413788 117378 413840
rect 49602 413244 49608 413296
rect 49660 413284 49666 413296
rect 59262 413284 59268 413296
rect 49660 413256 59268 413284
rect 49660 413244 49666 413256
rect 59262 413244 59268 413256
rect 59320 413284 59326 413296
rect 66254 413284 66260 413296
rect 59320 413256 66260 413284
rect 59320 413244 59326 413256
rect 66254 413244 66260 413256
rect 66312 413244 66318 413296
rect 50798 412564 50804 412616
rect 50856 412604 50862 412616
rect 66806 412604 66812 412616
rect 50856 412576 66812 412604
rect 50856 412564 50862 412576
rect 66806 412564 66812 412576
rect 66864 412564 66870 412616
rect 162118 412020 162124 412072
rect 162176 412060 162182 412072
rect 162762 412060 162768 412072
rect 162176 412032 162768 412060
rect 162176 412020 162182 412032
rect 162762 412020 162768 412032
rect 162820 412020 162826 412072
rect 41322 411884 41328 411936
rect 41380 411924 41386 411936
rect 50798 411924 50804 411936
rect 41380 411896 50804 411924
rect 41380 411884 41386 411896
rect 50798 411884 50804 411896
rect 50856 411884 50862 411936
rect 162762 411884 162768 411936
rect 162820 411924 162826 411936
rect 191466 411924 191472 411936
rect 162820 411896 191472 411924
rect 162820 411884 162826 411896
rect 191466 411884 191472 411896
rect 191524 411884 191530 411936
rect 255498 411544 255504 411596
rect 255556 411584 255562 411596
rect 258074 411584 258080 411596
rect 255556 411556 258080 411584
rect 255556 411544 255562 411556
rect 258074 411544 258080 411556
rect 258132 411544 258138 411596
rect 2958 411204 2964 411256
rect 3016 411244 3022 411256
rect 33778 411244 33784 411256
rect 3016 411216 33784 411244
rect 3016 411204 3022 411216
rect 33778 411204 33784 411216
rect 33836 411204 33842 411256
rect 50982 410524 50988 410576
rect 51040 410564 51046 410576
rect 62022 410564 62028 410576
rect 51040 410536 62028 410564
rect 51040 410524 51046 410536
rect 62022 410524 62028 410536
rect 62080 410564 62086 410576
rect 66898 410564 66904 410576
rect 62080 410536 66904 410564
rect 62080 410524 62086 410536
rect 66898 410524 66904 410536
rect 66956 410524 66962 410576
rect 255498 409912 255504 409964
rect 255556 409952 255562 409964
rect 258258 409952 258264 409964
rect 255556 409924 258264 409952
rect 255556 409912 255562 409924
rect 258258 409912 258264 409924
rect 258316 409912 258322 409964
rect 115842 409844 115848 409896
rect 115900 409884 115906 409896
rect 155218 409884 155224 409896
rect 115900 409856 155224 409884
rect 115900 409844 115906 409856
rect 155218 409844 155224 409856
rect 155276 409844 155282 409896
rect 187510 409844 187516 409896
rect 187568 409884 187574 409896
rect 190822 409884 190828 409896
rect 187568 409856 190828 409884
rect 187568 409844 187574 409856
rect 190822 409844 190828 409856
rect 190880 409844 190886 409896
rect 52454 409776 52460 409828
rect 52512 409816 52518 409828
rect 53650 409816 53656 409828
rect 52512 409788 53656 409816
rect 52512 409776 52518 409788
rect 53650 409776 53656 409788
rect 53708 409816 53714 409828
rect 66806 409816 66812 409828
rect 53708 409788 66812 409816
rect 53708 409776 53714 409788
rect 66806 409776 66812 409788
rect 66864 409776 66870 409828
rect 44082 409096 44088 409148
rect 44140 409136 44146 409148
rect 52454 409136 52460 409148
rect 44140 409108 52460 409136
rect 44140 409096 44146 409108
rect 52454 409096 52460 409108
rect 52512 409096 52518 409148
rect 115842 409096 115848 409148
rect 115900 409136 115906 409148
rect 124858 409136 124864 409148
rect 115900 409108 124864 409136
rect 115900 409096 115906 409108
rect 124858 409096 124864 409108
rect 124916 409096 124922 409148
rect 126882 408552 126888 408604
rect 126940 408592 126946 408604
rect 143534 408592 143540 408604
rect 126940 408564 143540 408592
rect 126940 408552 126946 408564
rect 143534 408552 143540 408564
rect 143592 408592 143598 408604
rect 144178 408592 144184 408604
rect 143592 408564 144184 408592
rect 143592 408552 143598 408564
rect 144178 408552 144184 408564
rect 144236 408552 144242 408604
rect 115842 408484 115848 408536
rect 115900 408524 115906 408536
rect 188338 408524 188344 408536
rect 115900 408496 188344 408524
rect 115900 408484 115906 408496
rect 188338 408484 188344 408496
rect 188396 408484 188402 408536
rect 255498 408484 255504 408536
rect 255556 408524 255562 408536
rect 276198 408524 276204 408536
rect 255556 408496 276204 408524
rect 255556 408484 255562 408496
rect 276198 408484 276204 408496
rect 276256 408484 276262 408536
rect 255498 407192 255504 407244
rect 255556 407232 255562 407244
rect 259546 407232 259552 407244
rect 255556 407204 259552 407232
rect 255556 407192 255562 407204
rect 259546 407192 259552 407204
rect 259604 407192 259610 407244
rect 52270 407124 52276 407176
rect 52328 407164 52334 407176
rect 66806 407164 66812 407176
rect 52328 407136 66812 407164
rect 52328 407124 52334 407136
rect 66806 407124 66812 407136
rect 66864 407124 66870 407176
rect 115842 407124 115848 407176
rect 115900 407164 115906 407176
rect 170398 407164 170404 407176
rect 115900 407136 170404 407164
rect 115900 407124 115906 407136
rect 170398 407124 170404 407136
rect 170456 407124 170462 407176
rect 162118 405764 162124 405816
rect 162176 405804 162182 405816
rect 191466 405804 191472 405816
rect 162176 405776 191472 405804
rect 162176 405764 162182 405776
rect 191466 405764 191472 405776
rect 191524 405764 191530 405816
rect 115750 405696 115756 405748
rect 115808 405736 115814 405748
rect 169018 405736 169024 405748
rect 115808 405708 169024 405736
rect 115808 405696 115814 405708
rect 169018 405696 169024 405708
rect 169076 405696 169082 405748
rect 255498 405696 255504 405748
rect 255556 405736 255562 405748
rect 274726 405736 274732 405748
rect 255556 405708 274732 405736
rect 255556 405696 255562 405708
rect 274726 405696 274732 405708
rect 274784 405696 274790 405748
rect 115842 405628 115848 405680
rect 115900 405668 115906 405680
rect 126882 405668 126888 405680
rect 115900 405640 126888 405668
rect 115900 405628 115906 405640
rect 126882 405628 126888 405640
rect 126940 405628 126946 405680
rect 62022 404336 62028 404388
rect 62080 404376 62086 404388
rect 66898 404376 66904 404388
rect 62080 404348 66904 404376
rect 62080 404336 62086 404348
rect 66898 404336 66904 404348
rect 66956 404336 66962 404388
rect 182910 404336 182916 404388
rect 182968 404376 182974 404388
rect 191374 404376 191380 404388
rect 182968 404348 191380 404376
rect 182968 404336 182974 404348
rect 191374 404336 191380 404348
rect 191432 404336 191438 404388
rect 255498 403384 255504 403436
rect 255556 403424 255562 403436
rect 257338 403424 257344 403436
rect 255556 403396 257344 403424
rect 255556 403384 255562 403396
rect 257338 403384 257344 403396
rect 257396 403384 257402 403436
rect 159358 403044 159364 403096
rect 159416 403084 159422 403096
rect 191466 403084 191472 403096
rect 159416 403056 191472 403084
rect 159416 403044 159422 403056
rect 191466 403044 191472 403056
rect 191524 403044 191530 403096
rect 54938 402976 54944 403028
rect 54996 403016 55002 403028
rect 66806 403016 66812 403028
rect 54996 402988 66812 403016
rect 54996 402976 55002 402988
rect 66806 402976 66812 402988
rect 66864 402976 66870 403028
rect 115842 402976 115848 403028
rect 115900 403016 115906 403028
rect 185762 403016 185768 403028
rect 115900 402988 185768 403016
rect 115900 402976 115906 402988
rect 185762 402976 185768 402988
rect 185820 402976 185826 403028
rect 114738 401344 114744 401396
rect 114796 401384 114802 401396
rect 116670 401384 116676 401396
rect 114796 401356 116676 401384
rect 114796 401344 114802 401356
rect 116670 401344 116676 401356
rect 116728 401344 116734 401396
rect 118786 400868 118792 400920
rect 118844 400908 118850 400920
rect 128354 400908 128360 400920
rect 118844 400880 128360 400908
rect 118844 400868 118850 400880
rect 128354 400868 128360 400880
rect 128412 400868 128418 400920
rect 187602 400732 187608 400784
rect 187660 400772 187666 400784
rect 191466 400772 191472 400784
rect 187660 400744 191472 400772
rect 187660 400732 187666 400744
rect 191466 400732 191472 400744
rect 191524 400732 191530 400784
rect 53650 400188 53656 400240
rect 53708 400228 53714 400240
rect 66714 400228 66720 400240
rect 53708 400200 66720 400228
rect 53708 400188 53714 400200
rect 66714 400188 66720 400200
rect 66772 400188 66778 400240
rect 115658 400188 115664 400240
rect 115716 400228 115722 400240
rect 152458 400228 152464 400240
rect 115716 400200 152464 400228
rect 115716 400188 115722 400200
rect 152458 400188 152464 400200
rect 152516 400188 152522 400240
rect 184382 400188 184388 400240
rect 184440 400228 184446 400240
rect 187602 400228 187608 400240
rect 184440 400200 187608 400228
rect 184440 400188 184446 400200
rect 187602 400188 187608 400200
rect 187660 400188 187666 400240
rect 255498 400188 255504 400240
rect 255556 400228 255562 400240
rect 277486 400228 277492 400240
rect 255556 400200 277492 400228
rect 255556 400188 255562 400200
rect 277486 400188 277492 400200
rect 277544 400188 277550 400240
rect 289722 399440 289728 399492
rect 289780 399480 289786 399492
rect 582742 399480 582748 399492
rect 289780 399452 582748 399480
rect 289780 399440 289786 399452
rect 582742 399440 582748 399452
rect 582800 399440 582806 399492
rect 115842 398828 115848 398880
rect 115900 398868 115906 398880
rect 151078 398868 151084 398880
rect 115900 398840 151084 398868
rect 115900 398828 115906 398840
rect 151078 398828 151084 398840
rect 151136 398828 151142 398880
rect 174538 398828 174544 398880
rect 174596 398868 174602 398880
rect 190822 398868 190828 398880
rect 174596 398840 190828 398868
rect 174596 398828 174602 398840
rect 190822 398828 190828 398840
rect 190880 398828 190886 398880
rect 255498 398828 255504 398880
rect 255556 398868 255562 398880
rect 258350 398868 258356 398880
rect 255556 398840 258356 398868
rect 255556 398828 255562 398840
rect 258350 398828 258356 398840
rect 258408 398868 258414 398880
rect 288710 398868 288716 398880
rect 258408 398840 288716 398868
rect 258408 398828 258414 398840
rect 288710 398828 288716 398840
rect 288768 398868 288774 398880
rect 289722 398868 289728 398880
rect 288768 398840 289728 398868
rect 288768 398828 288774 398840
rect 289722 398828 289728 398840
rect 289780 398828 289786 398880
rect 291102 398080 291108 398132
rect 291160 398120 291166 398132
rect 582466 398120 582472 398132
rect 291160 398092 582472 398120
rect 291160 398080 291166 398092
rect 582466 398080 582472 398092
rect 582524 398080 582530 398132
rect 115566 397536 115572 397588
rect 115624 397576 115630 397588
rect 117958 397576 117964 397588
rect 115624 397548 117964 397576
rect 115624 397536 115630 397548
rect 117958 397536 117964 397548
rect 118016 397576 118022 397588
rect 118786 397576 118792 397588
rect 118016 397548 118792 397576
rect 118016 397536 118022 397548
rect 118786 397536 118792 397548
rect 118844 397536 118850 397588
rect 180242 397536 180248 397588
rect 180300 397576 180306 397588
rect 191098 397576 191104 397588
rect 180300 397548 191104 397576
rect 180300 397536 180306 397548
rect 191098 397536 191104 397548
rect 191156 397536 191162 397588
rect 7558 397468 7564 397520
rect 7616 397508 7622 397520
rect 67726 397508 67732 397520
rect 7616 397480 67732 397508
rect 7616 397468 7622 397480
rect 67726 397468 67732 397480
rect 67784 397468 67790 397520
rect 113818 397468 113824 397520
rect 113876 397508 113882 397520
rect 188522 397508 188528 397520
rect 113876 397480 188528 397508
rect 113876 397468 113882 397480
rect 188522 397468 188528 397480
rect 188580 397468 188586 397520
rect 255498 397468 255504 397520
rect 255556 397508 255562 397520
rect 289814 397508 289820 397520
rect 255556 397480 289820 397508
rect 255556 397468 255562 397480
rect 289814 397468 289820 397480
rect 289872 397508 289878 397520
rect 291102 397508 291108 397520
rect 289872 397480 291108 397508
rect 289872 397468 289878 397480
rect 291102 397468 291108 397480
rect 291160 397468 291166 397520
rect 176746 397400 176752 397452
rect 176804 397440 176810 397452
rect 177942 397440 177948 397452
rect 176804 397412 177948 397440
rect 176804 397400 176810 397412
rect 177942 397400 177948 397412
rect 178000 397440 178006 397452
rect 191466 397440 191472 397452
rect 178000 397412 191472 397440
rect 178000 397400 178006 397412
rect 191466 397400 191472 397412
rect 191524 397400 191530 397452
rect 115842 396312 115848 396364
rect 115900 396352 115906 396364
rect 122098 396352 122104 396364
rect 115900 396324 122104 396352
rect 115900 396312 115906 396324
rect 122098 396312 122104 396324
rect 122156 396312 122162 396364
rect 127618 396040 127624 396092
rect 127676 396080 127682 396092
rect 191190 396080 191196 396092
rect 127676 396052 191196 396080
rect 127676 396040 127682 396052
rect 191190 396040 191196 396052
rect 191248 396080 191254 396092
rect 191374 396080 191380 396092
rect 191248 396052 191380 396080
rect 191248 396040 191254 396052
rect 191374 396040 191380 396052
rect 191432 396040 191438 396092
rect 64598 395428 64604 395480
rect 64656 395468 64662 395480
rect 67174 395468 67180 395480
rect 64656 395440 67180 395468
rect 64656 395428 64662 395440
rect 67174 395428 67180 395440
rect 67232 395428 67238 395480
rect 115842 394680 115848 394732
rect 115900 394720 115906 394732
rect 181530 394720 181536 394732
rect 115900 394692 181536 394720
rect 115900 394680 115906 394692
rect 181530 394680 181536 394692
rect 181588 394680 181594 394732
rect 60550 393388 60556 393440
rect 60608 393428 60614 393440
rect 65886 393428 65892 393440
rect 60608 393400 65892 393428
rect 60608 393388 60614 393400
rect 65886 393388 65892 393400
rect 65944 393388 65950 393440
rect 128998 393388 129004 393440
rect 129056 393428 129062 393440
rect 193398 393428 193404 393440
rect 129056 393400 193404 393428
rect 129056 393388 129062 393400
rect 193398 393388 193404 393400
rect 193456 393388 193462 393440
rect 59078 393320 59084 393372
rect 59136 393360 59142 393372
rect 66806 393360 66812 393372
rect 59136 393332 66812 393360
rect 59136 393320 59142 393332
rect 66806 393320 66812 393332
rect 66864 393320 66870 393372
rect 115842 393320 115848 393372
rect 115900 393360 115906 393372
rect 188430 393360 188436 393372
rect 115900 393332 188436 393360
rect 115900 393320 115906 393332
rect 188430 393320 188436 393332
rect 188488 393320 188494 393372
rect 255590 393320 255596 393372
rect 255648 393360 255654 393372
rect 271966 393360 271972 393372
rect 255648 393332 271972 393360
rect 255648 393320 255654 393332
rect 271966 393320 271972 393332
rect 272024 393320 272030 393372
rect 115842 392572 115848 392624
rect 115900 392612 115906 392624
rect 122834 392612 122840 392624
rect 115900 392584 122840 392612
rect 115900 392572 115906 392584
rect 122834 392572 122840 392584
rect 122892 392612 122898 392624
rect 123478 392612 123484 392624
rect 122892 392584 123484 392612
rect 122892 392572 122898 392584
rect 123478 392572 123484 392584
rect 123536 392572 123542 392624
rect 56410 391960 56416 392012
rect 56468 392000 56474 392012
rect 66254 392000 66260 392012
rect 56468 391972 66260 392000
rect 56468 391960 56474 391972
rect 66254 391960 66260 391972
rect 66312 391960 66318 392012
rect 188522 391892 188528 391944
rect 188580 391932 188586 391944
rect 191466 391932 191472 391944
rect 188580 391904 191472 391932
rect 188580 391892 188586 391904
rect 191466 391892 191472 391904
rect 191524 391892 191530 391944
rect 253566 391552 253572 391604
rect 253624 391592 253630 391604
rect 254026 391592 254032 391604
rect 253624 391564 254032 391592
rect 253624 391552 253630 391564
rect 254026 391552 254032 391564
rect 254084 391552 254090 391604
rect 250530 390940 250536 390992
rect 250588 390980 250594 390992
rect 258074 390980 258080 390992
rect 250588 390952 258080 390980
rect 250588 390940 250594 390952
rect 258074 390940 258080 390952
rect 258132 390940 258138 390992
rect 114830 390736 114836 390788
rect 114888 390776 114894 390788
rect 116578 390776 116584 390788
rect 114888 390748 116584 390776
rect 114888 390736 114894 390748
rect 116578 390736 116584 390748
rect 116636 390736 116642 390788
rect 67358 390600 67364 390652
rect 67416 390640 67422 390652
rect 73798 390640 73804 390652
rect 67416 390612 73804 390640
rect 67416 390600 67422 390612
rect 73798 390600 73804 390612
rect 73856 390600 73862 390652
rect 191006 390600 191012 390652
rect 191064 390640 191070 390652
rect 203518 390640 203524 390652
rect 191064 390612 203524 390640
rect 191064 390600 191070 390612
rect 203518 390600 203524 390612
rect 203576 390600 203582 390652
rect 69658 390532 69664 390584
rect 69716 390572 69722 390584
rect 163590 390572 163596 390584
rect 69716 390544 163596 390572
rect 69716 390532 69722 390544
rect 163590 390532 163596 390544
rect 163648 390572 163654 390584
rect 194134 390572 194140 390584
rect 163648 390544 194140 390572
rect 163648 390532 163654 390544
rect 194134 390532 194140 390544
rect 194192 390532 194198 390584
rect 96706 390464 96712 390516
rect 96764 390504 96770 390516
rect 97534 390504 97540 390516
rect 96764 390476 97540 390504
rect 96764 390464 96770 390476
rect 97534 390464 97540 390476
rect 97592 390464 97598 390516
rect 67634 390124 67640 390176
rect 67692 390164 67698 390176
rect 68784 390164 68790 390176
rect 67692 390136 68790 390164
rect 67692 390124 67698 390136
rect 68784 390124 68790 390136
rect 68842 390124 68848 390176
rect 56502 389784 56508 389836
rect 56560 389824 56566 389836
rect 86770 389824 86776 389836
rect 56560 389796 86776 389824
rect 56560 389784 56566 389796
rect 86770 389784 86776 389796
rect 86828 389824 86834 389836
rect 87782 389824 87788 389836
rect 86828 389796 87788 389824
rect 86828 389784 86834 389796
rect 87782 389784 87788 389796
rect 87840 389784 87846 389836
rect 242158 389784 242164 389836
rect 242216 389824 242222 389836
rect 254118 389824 254124 389836
rect 242216 389796 254124 389824
rect 242216 389784 242222 389796
rect 254118 389784 254124 389796
rect 254176 389784 254182 389836
rect 75086 389240 75092 389292
rect 75144 389280 75150 389292
rect 164970 389280 164976 389292
rect 75144 389252 164976 389280
rect 75144 389240 75150 389252
rect 164970 389240 164976 389252
rect 165028 389280 165034 389292
rect 202046 389280 202052 389292
rect 165028 389252 202052 389280
rect 165028 389240 165034 389252
rect 202046 389240 202052 389252
rect 202104 389240 202110 389292
rect 249242 389240 249248 389292
rect 249300 389280 249306 389292
rect 253658 389280 253664 389292
rect 249300 389252 253664 389280
rect 249300 389240 249306 389252
rect 253658 389240 253664 389252
rect 253716 389240 253722 389292
rect 94682 389172 94688 389224
rect 94740 389212 94746 389224
rect 227714 389212 227720 389224
rect 94740 389184 227720 389212
rect 94740 389172 94746 389184
rect 227714 389172 227720 389184
rect 227772 389212 227778 389224
rect 228542 389212 228548 389224
rect 227772 389184 228548 389212
rect 227772 389172 227778 389184
rect 228542 389172 228548 389184
rect 228600 389172 228606 389224
rect 234890 389172 234896 389224
rect 234948 389212 234954 389224
rect 249702 389212 249708 389224
rect 234948 389184 249708 389212
rect 234948 389172 234954 389184
rect 249702 389172 249708 389184
rect 249760 389172 249766 389224
rect 65978 389104 65984 389156
rect 66036 389144 66042 389156
rect 71682 389144 71688 389156
rect 66036 389116 71688 389144
rect 66036 389104 66042 389116
rect 71682 389104 71688 389116
rect 71740 389144 71746 389156
rect 72602 389144 72608 389156
rect 71740 389116 72608 389144
rect 71740 389104 71746 389116
rect 72602 389104 72608 389116
rect 72660 389104 72666 389156
rect 111886 389104 111892 389156
rect 111944 389144 111950 389156
rect 251818 389144 251824 389156
rect 111944 389116 251824 389144
rect 111944 389104 111950 389116
rect 251818 389104 251824 389116
rect 251876 389104 251882 389156
rect 241974 389036 241980 389088
rect 242032 389076 242038 389088
rect 273898 389076 273904 389088
rect 242032 389048 273904 389076
rect 242032 389036 242038 389048
rect 273898 389036 273904 389048
rect 273956 389036 273962 389088
rect 234062 388696 234068 388748
rect 234120 388736 234126 388748
rect 234522 388736 234528 388748
rect 234120 388708 234528 388736
rect 234120 388696 234126 388708
rect 234522 388696 234528 388708
rect 234580 388736 234586 388748
rect 239030 388736 239036 388748
rect 234580 388708 239036 388736
rect 234580 388696 234586 388708
rect 239030 388696 239036 388708
rect 239088 388696 239094 388748
rect 120718 388016 120724 388068
rect 120776 388056 120782 388068
rect 121546 388056 121552 388068
rect 120776 388028 121552 388056
rect 120776 388016 120782 388028
rect 121546 388016 121552 388028
rect 121604 388016 121610 388068
rect 57698 387812 57704 387864
rect 57756 387852 57762 387864
rect 66070 387852 66076 387864
rect 57756 387824 66076 387852
rect 57756 387812 57762 387824
rect 66070 387812 66076 387824
rect 66128 387812 66134 387864
rect 121454 387812 121460 387864
rect 121512 387812 121518 387864
rect 129090 387812 129096 387864
rect 129148 387852 129154 387864
rect 129734 387852 129740 387864
rect 129148 387824 129740 387852
rect 129148 387812 129154 387824
rect 129734 387812 129740 387824
rect 129792 387812 129798 387864
rect 214558 387812 214564 387864
rect 214616 387852 214622 387864
rect 216214 387852 216220 387864
rect 214616 387824 216220 387852
rect 214616 387812 214622 387824
rect 216214 387812 216220 387824
rect 216272 387812 216278 387864
rect 232498 387812 232504 387864
rect 232556 387852 232562 387864
rect 233326 387852 233332 387864
rect 232556 387824 233332 387852
rect 232556 387812 232562 387824
rect 233326 387812 233332 387824
rect 233384 387812 233390 387864
rect 241974 387812 241980 387864
rect 242032 387852 242038 387864
rect 242802 387852 242808 387864
rect 242032 387824 242808 387852
rect 242032 387812 242038 387824
rect 242802 387812 242808 387824
rect 242860 387812 242866 387864
rect 3418 387744 3424 387796
rect 3476 387784 3482 387796
rect 93946 387784 93952 387796
rect 3476 387756 93952 387784
rect 3476 387744 3482 387756
rect 93946 387744 93952 387756
rect 94004 387784 94010 387796
rect 94498 387784 94504 387796
rect 94004 387756 94504 387784
rect 94004 387744 94010 387756
rect 94498 387744 94504 387756
rect 94556 387744 94562 387796
rect 99466 387744 99472 387796
rect 99524 387784 99530 387796
rect 104158 387784 104164 387796
rect 99524 387756 104164 387784
rect 99524 387744 99530 387756
rect 104158 387744 104164 387756
rect 104216 387744 104222 387796
rect 108942 387744 108948 387796
rect 109000 387784 109006 387796
rect 114646 387784 114652 387796
rect 109000 387756 114652 387784
rect 109000 387744 109006 387756
rect 114646 387744 114652 387756
rect 114704 387744 114710 387796
rect 118786 387744 118792 387796
rect 118844 387784 118850 387796
rect 121472 387784 121500 387812
rect 218238 387784 218244 387796
rect 118844 387756 218244 387784
rect 118844 387744 118850 387756
rect 218238 387744 218244 387756
rect 218296 387784 218302 387796
rect 219250 387784 219256 387796
rect 218296 387756 219256 387784
rect 218296 387744 218302 387756
rect 219250 387744 219256 387756
rect 219308 387744 219314 387796
rect 101674 387676 101680 387728
rect 101732 387716 101738 387728
rect 125594 387716 125600 387728
rect 101732 387688 125600 387716
rect 101732 387676 101738 387688
rect 125594 387676 125600 387688
rect 125652 387716 125658 387728
rect 126238 387716 126244 387728
rect 125652 387688 126244 387716
rect 125652 387676 125658 387688
rect 126238 387676 126244 387688
rect 126296 387676 126302 387728
rect 180150 387676 180156 387728
rect 180208 387716 180214 387728
rect 255406 387716 255412 387728
rect 180208 387688 255412 387716
rect 180208 387676 180214 387688
rect 255406 387676 255412 387688
rect 255464 387676 255470 387728
rect 219250 387064 219256 387116
rect 219308 387104 219314 387116
rect 232590 387104 232596 387116
rect 219308 387076 232596 387104
rect 219308 387064 219314 387076
rect 232590 387064 232596 387076
rect 232648 387064 232654 387116
rect 253382 387064 253388 387116
rect 253440 387104 253446 387116
rect 267826 387104 267832 387116
rect 253440 387076 267832 387104
rect 253440 387064 253446 387076
rect 267826 387064 267832 387076
rect 267884 387064 267890 387116
rect 77294 386996 77300 387048
rect 77352 387036 77358 387048
rect 78030 387036 78036 387048
rect 77352 387008 78036 387036
rect 77352 386996 77358 387008
rect 78030 386996 78036 387008
rect 78088 386996 78094 387048
rect 84194 386996 84200 387048
rect 84252 387036 84258 387048
rect 85022 387036 85028 387048
rect 84252 387008 85028 387036
rect 84252 386996 84258 387008
rect 85022 386996 85028 387008
rect 85080 386996 85086 387048
rect 109034 386996 109040 387048
rect 109092 387036 109098 387048
rect 109494 387036 109500 387048
rect 109092 387008 109500 387036
rect 109092 386996 109098 387008
rect 109494 386996 109500 387008
rect 109552 386996 109558 387048
rect 223574 386996 223580 387048
rect 223632 387036 223638 387048
rect 224494 387036 224500 387048
rect 223632 387008 224500 387036
rect 223632 386996 223638 387008
rect 224494 386996 224500 387008
rect 224552 386996 224558 387048
rect 67818 386316 67824 386368
rect 67876 386356 67882 386368
rect 174538 386356 174544 386368
rect 67876 386328 174544 386356
rect 67876 386316 67882 386328
rect 174538 386316 174544 386328
rect 174596 386316 174602 386368
rect 186958 386316 186964 386368
rect 187016 386356 187022 386368
rect 208486 386356 208492 386368
rect 187016 386328 208492 386356
rect 187016 386316 187022 386328
rect 208486 386316 208492 386328
rect 208544 386316 208550 386368
rect 231118 386316 231124 386368
rect 231176 386356 231182 386368
rect 234246 386356 234252 386368
rect 231176 386328 234252 386356
rect 231176 386316 231182 386328
rect 234246 386316 234252 386328
rect 234304 386316 234310 386368
rect 103146 385636 103152 385688
rect 103204 385676 103210 385688
rect 187602 385676 187608 385688
rect 103204 385648 187608 385676
rect 103204 385636 103210 385648
rect 187602 385636 187608 385648
rect 187660 385636 187666 385688
rect 89622 385024 89628 385076
rect 89680 385064 89686 385076
rect 94314 385064 94320 385076
rect 89680 385036 94320 385064
rect 89680 385024 89686 385036
rect 94314 385024 94320 385036
rect 94372 385024 94378 385076
rect 231854 385024 231860 385076
rect 231912 385064 231918 385076
rect 281718 385064 281724 385076
rect 231912 385036 281724 385064
rect 231912 385024 231918 385036
rect 281718 385024 281724 385036
rect 281776 385024 281782 385076
rect 86862 384956 86868 385008
rect 86920 384996 86926 385008
rect 118786 384996 118792 385008
rect 86920 384968 118792 384996
rect 86920 384956 86926 384968
rect 118786 384956 118792 384968
rect 118844 384956 118850 385008
rect 190270 384956 190276 385008
rect 190328 384996 190334 385008
rect 216398 384996 216404 385008
rect 190328 384968 216404 384996
rect 190328 384956 190334 384968
rect 216398 384956 216404 384968
rect 216456 384956 216462 385008
rect 100386 384888 100392 384940
rect 100444 384928 100450 384940
rect 126882 384928 126888 384940
rect 100444 384900 126888 384928
rect 100444 384888 100450 384900
rect 126882 384888 126888 384900
rect 126940 384888 126946 384940
rect 119982 384276 119988 384328
rect 120040 384316 120046 384328
rect 186314 384316 186320 384328
rect 120040 384288 186320 384316
rect 120040 384276 120046 384288
rect 186314 384276 186320 384288
rect 186372 384316 186378 384328
rect 220998 384316 221004 384328
rect 186372 384288 221004 384316
rect 186372 384276 186378 384288
rect 220998 384276 221004 384288
rect 221056 384276 221062 384328
rect 244918 384276 244924 384328
rect 244976 384316 244982 384328
rect 259546 384316 259552 384328
rect 244976 384288 259552 384316
rect 244976 384276 244982 384288
rect 259546 384276 259552 384288
rect 259604 384276 259610 384328
rect 216398 383664 216404 383716
rect 216456 383704 216462 383716
rect 240226 383704 240232 383716
rect 216456 383676 240232 383704
rect 216456 383664 216462 383676
rect 240226 383664 240232 383676
rect 240284 383664 240290 383716
rect 242986 383664 242992 383716
rect 243044 383704 243050 383716
rect 243814 383704 243820 383716
rect 243044 383676 243820 383704
rect 243044 383664 243050 383676
rect 243814 383664 243820 383676
rect 243872 383664 243878 383716
rect 243998 383664 244004 383716
rect 244056 383704 244062 383716
rect 247678 383704 247684 383716
rect 244056 383676 247684 383704
rect 244056 383664 244062 383676
rect 247678 383664 247684 383676
rect 247736 383664 247742 383716
rect 97994 383596 98000 383648
rect 98052 383636 98058 383648
rect 120718 383636 120724 383648
rect 98052 383608 120724 383636
rect 98052 383596 98058 383608
rect 120718 383596 120724 383608
rect 120776 383596 120782 383648
rect 67726 382984 67732 383036
rect 67784 383024 67790 383036
rect 83458 383024 83464 383036
rect 67784 382996 83464 383024
rect 67784 382984 67790 382996
rect 83458 382984 83464 382996
rect 83516 382984 83522 383036
rect 80054 382916 80060 382968
rect 80112 382956 80118 382968
rect 106366 382956 106372 382968
rect 80112 382928 106372 382956
rect 80112 382916 80118 382928
rect 106366 382916 106372 382928
rect 106424 382956 106430 382968
rect 115934 382956 115940 382968
rect 106424 382928 115940 382956
rect 106424 382916 106430 382928
rect 115934 382916 115940 382928
rect 115992 382916 115998 382968
rect 125502 382916 125508 382968
rect 125560 382956 125566 382968
rect 231854 382956 231860 382968
rect 125560 382928 231860 382956
rect 125560 382916 125566 382928
rect 231854 382916 231860 382928
rect 231912 382916 231918 382968
rect 282914 382916 282920 382968
rect 282972 382956 282978 382968
rect 283098 382956 283104 382968
rect 282972 382928 283104 382956
rect 282972 382916 282978 382928
rect 283098 382916 283104 382928
rect 283156 382956 283162 382968
rect 582834 382956 582840 382968
rect 283156 382928 582840 382956
rect 283156 382916 283162 382928
rect 582834 382916 582840 382928
rect 582892 382916 582898 382968
rect 239398 382304 239404 382356
rect 239456 382344 239462 382356
rect 244274 382344 244280 382356
rect 239456 382316 244280 382344
rect 239456 382304 239462 382316
rect 244274 382304 244280 382316
rect 244332 382304 244338 382356
rect 226978 382236 226984 382288
rect 227036 382276 227042 382288
rect 273530 382276 273536 382288
rect 227036 382248 273536 382276
rect 227036 382236 227042 382248
rect 273530 382236 273536 382248
rect 273588 382236 273594 382288
rect 97718 382168 97724 382220
rect 97776 382208 97782 382220
rect 124214 382208 124220 382220
rect 97776 382180 124220 382208
rect 97776 382168 97782 382180
rect 124214 382168 124220 382180
rect 124272 382208 124278 382220
rect 125502 382208 125508 382220
rect 124272 382180 125508 382208
rect 124272 382168 124278 382180
rect 125502 382168 125508 382180
rect 125560 382168 125566 382220
rect 187602 382168 187608 382220
rect 187660 382208 187666 382220
rect 239122 382208 239128 382220
rect 187660 382180 239128 382208
rect 187660 382168 187666 382180
rect 239122 382168 239128 382180
rect 239180 382168 239186 382220
rect 111886 381692 111892 381744
rect 111944 381732 111950 381744
rect 112714 381732 112720 381744
rect 111944 381704 112720 381732
rect 111944 381692 111950 381704
rect 112714 381692 112720 381704
rect 112772 381692 112778 381744
rect 65978 381488 65984 381540
rect 66036 381528 66042 381540
rect 77386 381528 77392 381540
rect 66036 381500 77392 381528
rect 66036 381488 66042 381500
rect 77386 381488 77392 381500
rect 77444 381488 77450 381540
rect 188430 381488 188436 381540
rect 188488 381528 188494 381540
rect 223482 381528 223488 381540
rect 188488 381500 223488 381528
rect 188488 381488 188494 381500
rect 223482 381488 223488 381500
rect 223540 381488 223546 381540
rect 3418 380876 3424 380928
rect 3476 380916 3482 380928
rect 111886 380916 111892 380928
rect 3476 380888 111892 380916
rect 3476 380876 3482 380888
rect 111886 380876 111892 380888
rect 111944 380876 111950 380928
rect 230750 380876 230756 380928
rect 230808 380916 230814 380928
rect 273438 380916 273444 380928
rect 230808 380888 273444 380916
rect 230808 380876 230814 380888
rect 273438 380876 273444 380888
rect 273496 380876 273502 380928
rect 50982 380808 50988 380860
rect 51040 380848 51046 380860
rect 184290 380848 184296 380860
rect 51040 380820 184296 380848
rect 51040 380808 51046 380820
rect 184290 380808 184296 380820
rect 184348 380808 184354 380860
rect 189074 380808 189080 380860
rect 189132 380848 189138 380860
rect 189718 380848 189724 380860
rect 189132 380820 189724 380848
rect 189132 380808 189138 380820
rect 189718 380808 189724 380820
rect 189776 380848 189782 380860
rect 221274 380848 221280 380860
rect 189776 380820 221280 380848
rect 189776 380808 189782 380820
rect 221274 380808 221280 380820
rect 221332 380808 221338 380860
rect 223482 380808 223488 380860
rect 223540 380848 223546 380860
rect 251910 380848 251916 380860
rect 223540 380820 251916 380848
rect 223540 380808 223546 380820
rect 251910 380808 251916 380820
rect 251968 380808 251974 380860
rect 109126 380128 109132 380180
rect 109184 380168 109190 380180
rect 163498 380168 163504 380180
rect 109184 380140 163504 380168
rect 109184 380128 109190 380140
rect 163498 380128 163504 380140
rect 163556 380128 163562 380180
rect 246390 380128 246396 380180
rect 246448 380168 246454 380180
rect 254210 380168 254216 380180
rect 246448 380140 254216 380168
rect 246448 380128 246454 380140
rect 254210 380128 254216 380140
rect 254268 380128 254274 380180
rect 50706 379516 50712 379568
rect 50764 379556 50770 379568
rect 50982 379556 50988 379568
rect 50764 379528 50988 379556
rect 50764 379516 50770 379528
rect 50982 379516 50988 379528
rect 51040 379516 51046 379568
rect 52270 379448 52276 379500
rect 52328 379488 52334 379500
rect 130378 379488 130384 379500
rect 52328 379460 130384 379488
rect 52328 379448 52334 379460
rect 130378 379448 130384 379460
rect 130436 379448 130442 379500
rect 240226 379448 240232 379500
rect 240284 379488 240290 379500
rect 582926 379488 582932 379500
rect 240284 379460 582932 379488
rect 240284 379448 240290 379460
rect 582926 379448 582932 379460
rect 582984 379448 582990 379500
rect 92474 379380 92480 379432
rect 92532 379420 92538 379432
rect 125686 379420 125692 379432
rect 92532 379392 125692 379420
rect 92532 379380 92538 379392
rect 125686 379380 125692 379392
rect 125744 379420 125750 379432
rect 126422 379420 126428 379432
rect 125744 379392 126428 379420
rect 125744 379380 125750 379392
rect 126422 379380 126428 379392
rect 126480 379380 126486 379432
rect 129090 379380 129096 379432
rect 129148 379420 129154 379432
rect 204254 379420 204260 379432
rect 129148 379392 204260 379420
rect 129148 379380 129154 379392
rect 204254 379380 204260 379392
rect 204312 379380 204318 379432
rect 185762 379312 185768 379364
rect 185820 379352 185826 379364
rect 244918 379352 244924 379364
rect 185820 379324 244924 379352
rect 185820 379312 185826 379324
rect 244918 379312 244924 379324
rect 244976 379312 244982 379364
rect 245746 378156 245752 378208
rect 245804 378196 245810 378208
rect 246298 378196 246304 378208
rect 245804 378168 246304 378196
rect 245804 378156 245810 378168
rect 246298 378156 246304 378168
rect 246356 378196 246362 378208
rect 269298 378196 269304 378208
rect 246356 378168 269304 378196
rect 246356 378156 246362 378168
rect 269298 378156 269304 378168
rect 269356 378156 269362 378208
rect 67266 378088 67272 378140
rect 67324 378128 67330 378140
rect 162118 378128 162124 378140
rect 67324 378100 162124 378128
rect 67324 378088 67330 378100
rect 162118 378088 162124 378100
rect 162176 378088 162182 378140
rect 188338 378088 188344 378140
rect 188396 378128 188402 378140
rect 188890 378128 188896 378140
rect 188396 378100 188896 378128
rect 188396 378088 188402 378100
rect 188890 378088 188896 378100
rect 188948 378128 188954 378140
rect 256694 378128 256700 378140
rect 188948 378100 256700 378128
rect 188948 378088 188954 378100
rect 256694 378088 256700 378100
rect 256752 378088 256758 378140
rect 84286 377408 84292 377460
rect 84344 377448 84350 377460
rect 97258 377448 97264 377460
rect 84344 377420 97264 377448
rect 84344 377408 84350 377420
rect 97258 377408 97264 377420
rect 97316 377408 97322 377460
rect 97626 377408 97632 377460
rect 97684 377448 97690 377460
rect 118694 377448 118700 377460
rect 97684 377420 118700 377448
rect 97684 377408 97690 377420
rect 118694 377408 118700 377420
rect 118752 377448 118758 377460
rect 230750 377448 230756 377460
rect 118752 377420 230756 377448
rect 118752 377408 118758 377420
rect 230750 377408 230756 377420
rect 230808 377408 230814 377460
rect 256694 376728 256700 376780
rect 256752 376768 256758 376780
rect 257338 376768 257344 376780
rect 256752 376740 257344 376768
rect 256752 376728 256758 376740
rect 257338 376728 257344 376740
rect 257396 376768 257402 376780
rect 291286 376768 291292 376780
rect 257396 376740 291292 376768
rect 257396 376728 257402 376740
rect 291286 376728 291292 376740
rect 291344 376728 291350 376780
rect 73798 376592 73804 376644
rect 73856 376632 73862 376644
rect 159358 376632 159364 376644
rect 73856 376604 159364 376632
rect 73856 376592 73862 376604
rect 159358 376592 159364 376604
rect 159416 376592 159422 376644
rect 117958 376524 117964 376576
rect 118016 376564 118022 376576
rect 277486 376564 277492 376576
rect 118016 376536 277492 376564
rect 118016 376524 118022 376536
rect 277486 376524 277492 376536
rect 277544 376524 277550 376576
rect 58894 375980 58900 376032
rect 58952 376020 58958 376032
rect 76558 376020 76564 376032
rect 58952 375992 76564 376020
rect 58952 375980 58958 375992
rect 76558 375980 76564 375992
rect 76616 375980 76622 376032
rect 105538 375980 105544 376032
rect 105596 376020 105602 376032
rect 117958 376020 117964 376032
rect 105596 375992 117964 376020
rect 105596 375980 105602 375992
rect 117958 375980 117964 375992
rect 118016 375980 118022 376032
rect 88242 375300 88248 375352
rect 88300 375340 88306 375352
rect 91922 375340 91928 375352
rect 88300 375312 91928 375340
rect 88300 375300 88306 375312
rect 91922 375300 91928 375312
rect 91980 375340 91986 375352
rect 224954 375340 224960 375352
rect 91980 375312 224960 375340
rect 91980 375300 91986 375312
rect 224954 375300 224960 375312
rect 225012 375300 225018 375352
rect 72970 375232 72976 375284
rect 73028 375272 73034 375284
rect 168374 375272 168380 375284
rect 73028 375244 168380 375272
rect 73028 375232 73034 375244
rect 168374 375232 168380 375244
rect 168432 375232 168438 375284
rect 181530 375232 181536 375284
rect 181588 375272 181594 375284
rect 255498 375272 255504 375284
rect 181588 375244 255504 375272
rect 181588 375232 181594 375244
rect 255498 375232 255504 375244
rect 255556 375232 255562 375284
rect 170398 373940 170404 373992
rect 170456 373980 170462 373992
rect 242158 373980 242164 373992
rect 170456 373952 242164 373980
rect 170456 373940 170462 373952
rect 242158 373940 242164 373952
rect 242216 373940 242222 373992
rect 94498 373260 94504 373312
rect 94556 373300 94562 373312
rect 121454 373300 121460 373312
rect 94556 373272 121460 373300
rect 94556 373260 94562 373272
rect 121454 373260 121460 373272
rect 121512 373300 121518 373312
rect 226978 373300 226984 373312
rect 121512 373272 226984 373300
rect 121512 373260 121518 373272
rect 226978 373260 226984 373272
rect 227036 373260 227042 373312
rect 240778 373260 240784 373312
rect 240836 373300 240842 373312
rect 262214 373300 262220 373312
rect 240836 373272 262220 373300
rect 240836 373260 240842 373272
rect 262214 373260 262220 373272
rect 262272 373260 262278 373312
rect 106090 372512 106096 372564
rect 106148 372552 106154 372564
rect 242894 372552 242900 372564
rect 106148 372524 242900 372552
rect 106148 372512 106154 372524
rect 242894 372512 242900 372524
rect 242952 372512 242958 372564
rect 163498 372444 163504 372496
rect 163556 372484 163562 372496
rect 248414 372484 248420 372496
rect 163556 372456 248420 372484
rect 163556 372444 163562 372456
rect 248414 372444 248420 372456
rect 248472 372484 248478 372496
rect 250438 372484 250444 372496
rect 248472 372456 250444 372484
rect 248472 372444 248478 372456
rect 250438 372444 250444 372456
rect 250496 372444 250502 372496
rect 81434 371832 81440 371884
rect 81492 371872 81498 371884
rect 115934 371872 115940 371884
rect 81492 371844 115940 371872
rect 81492 371832 81498 371844
rect 115934 371832 115940 371844
rect 115992 371872 115998 371884
rect 117222 371872 117228 371884
rect 115992 371844 117228 371872
rect 115992 371832 115998 371844
rect 117222 371832 117228 371844
rect 117280 371832 117286 371884
rect 242894 371220 242900 371272
rect 242952 371260 242958 371272
rect 243538 371260 243544 371272
rect 242952 371232 243544 371260
rect 242952 371220 242958 371232
rect 243538 371220 243544 371232
rect 243596 371220 243602 371272
rect 102042 371152 102048 371204
rect 102100 371192 102106 371204
rect 235994 371192 236000 371204
rect 102100 371164 236000 371192
rect 102100 371152 102106 371164
rect 235994 371152 236000 371164
rect 236052 371152 236058 371204
rect 81250 370472 81256 370524
rect 81308 370512 81314 370524
rect 129090 370512 129096 370524
rect 81308 370484 129096 370512
rect 81308 370472 81314 370484
rect 129090 370472 129096 370484
rect 129148 370472 129154 370524
rect 187418 370472 187424 370524
rect 187476 370512 187482 370524
rect 197998 370512 198004 370524
rect 187476 370484 198004 370512
rect 187476 370472 187482 370484
rect 197998 370472 198004 370484
rect 198056 370472 198062 370524
rect 235994 369860 236000 369912
rect 236052 369900 236058 369912
rect 236638 369900 236644 369912
rect 236052 369872 236644 369900
rect 236052 369860 236058 369872
rect 236638 369860 236644 369872
rect 236696 369860 236702 369912
rect 111886 369792 111892 369844
rect 111944 369832 111950 369844
rect 274726 369832 274732 369844
rect 111944 369804 274732 369832
rect 111944 369792 111950 369804
rect 274726 369792 274732 369804
rect 274784 369792 274790 369844
rect 151078 369724 151084 369776
rect 151136 369764 151142 369776
rect 245838 369764 245844 369776
rect 151136 369736 245844 369764
rect 151136 369724 151142 369736
rect 245838 369724 245844 369736
rect 245896 369724 245902 369776
rect 245838 369316 245844 369368
rect 245896 369356 245902 369368
rect 246390 369356 246396 369368
rect 245896 369328 246396 369356
rect 245896 369316 245902 369328
rect 246390 369316 246396 369328
rect 246448 369316 246454 369368
rect 101398 369112 101404 369164
rect 101456 369152 101462 369164
rect 111886 369152 111892 369164
rect 101456 369124 111892 369152
rect 101456 369112 101462 369124
rect 111886 369112 111892 369124
rect 111944 369112 111950 369164
rect 126422 368432 126428 368484
rect 126480 368472 126486 368484
rect 226334 368472 226340 368484
rect 126480 368444 226340 368472
rect 126480 368432 126486 368444
rect 226334 368432 226340 368444
rect 226392 368472 226398 368484
rect 226978 368472 226984 368484
rect 226392 368444 226984 368472
rect 226392 368432 226398 368444
rect 226978 368432 226984 368444
rect 227036 368432 227042 368484
rect 67634 368364 67640 368416
rect 67692 368404 67698 368416
rect 128998 368404 129004 368416
rect 67692 368376 129004 368404
rect 67692 368364 67698 368376
rect 128998 368364 129004 368376
rect 129056 368364 129062 368416
rect 152458 368364 152464 368416
rect 152516 368404 152522 368416
rect 252554 368404 252560 368416
rect 152516 368376 252560 368404
rect 152516 368364 152522 368376
rect 252554 368364 252560 368376
rect 252612 368364 252618 368416
rect 59078 367004 59084 367056
rect 59136 367044 59142 367056
rect 59136 367016 183508 367044
rect 59136 367004 59142 367016
rect 88978 366936 88984 366988
rect 89036 366976 89042 366988
rect 183480 366976 183508 367016
rect 183554 367004 183560 367056
rect 183612 367044 183618 367056
rect 184382 367044 184388 367056
rect 183612 367016 184388 367044
rect 183612 367004 183618 367016
rect 184382 367004 184388 367016
rect 184440 367004 184446 367056
rect 189074 366976 189080 366988
rect 89036 366948 180794 366976
rect 183480 366948 189080 366976
rect 89036 366936 89042 366948
rect 180766 366840 180794 366948
rect 189074 366936 189080 366948
rect 189132 366936 189138 366988
rect 183554 366840 183560 366852
rect 180766 366812 183560 366840
rect 183554 366800 183560 366812
rect 183612 366800 183618 366852
rect 188798 366324 188804 366376
rect 188856 366364 188862 366376
rect 207106 366364 207112 366376
rect 188856 366336 207112 366364
rect 188856 366324 188862 366336
rect 207106 366324 207112 366336
rect 207164 366324 207170 366376
rect 108850 365644 108856 365696
rect 108908 365684 108914 365696
rect 246298 365684 246304 365696
rect 108908 365656 246304 365684
rect 108908 365644 108914 365656
rect 246298 365644 246304 365656
rect 246356 365644 246362 365696
rect 86770 364964 86776 365016
rect 86828 365004 86834 365016
rect 128998 365004 129004 365016
rect 86828 364976 129004 365004
rect 86828 364964 86834 364976
rect 128998 364964 129004 364976
rect 129056 364964 129062 365016
rect 170490 364352 170496 364404
rect 170548 364392 170554 364404
rect 213822 364392 213828 364404
rect 170548 364364 213828 364392
rect 170548 364352 170554 364364
rect 213822 364352 213828 364364
rect 213880 364352 213886 364404
rect 116578 364284 116584 364336
rect 116636 364324 116642 364336
rect 254026 364324 254032 364336
rect 116636 364296 254032 364324
rect 116636 364284 116642 364296
rect 254026 364284 254032 364296
rect 254084 364284 254090 364336
rect 71682 363604 71688 363656
rect 71740 363644 71746 363656
rect 195882 363644 195888 363656
rect 71740 363616 195888 363644
rect 71740 363604 71746 363616
rect 195882 363604 195888 363616
rect 195940 363604 195946 363656
rect 254026 362924 254032 362976
rect 254084 362964 254090 362976
rect 259546 362964 259552 362976
rect 254084 362936 259552 362964
rect 254084 362924 254090 362936
rect 259546 362924 259552 362936
rect 259604 362924 259610 362976
rect 77294 362856 77300 362908
rect 77352 362896 77358 362908
rect 205726 362896 205732 362908
rect 77352 362868 205732 362896
rect 77352 362856 77358 362868
rect 205726 362856 205732 362868
rect 205784 362856 205790 362908
rect 213822 362856 213828 362908
rect 213880 362896 213886 362908
rect 231118 362896 231124 362908
rect 213880 362868 231124 362896
rect 213880 362856 213886 362868
rect 231118 362856 231124 362868
rect 231176 362856 231182 362908
rect 195882 362788 195888 362840
rect 195940 362828 195946 362840
rect 198734 362828 198740 362840
rect 195940 362800 198740 362828
rect 195940 362788 195946 362800
rect 198734 362788 198740 362800
rect 198792 362788 198798 362840
rect 86862 362176 86868 362228
rect 86920 362216 86926 362228
rect 187694 362216 187700 362228
rect 86920 362188 187700 362216
rect 86920 362176 86926 362188
rect 187694 362176 187700 362188
rect 187752 362176 187758 362228
rect 198734 362176 198740 362228
rect 198792 362216 198798 362228
rect 293954 362216 293960 362228
rect 198792 362188 293960 362216
rect 198792 362176 198798 362188
rect 293954 362176 293960 362188
rect 294012 362176 294018 362228
rect 69014 361496 69020 361548
rect 69072 361536 69078 361548
rect 194594 361536 194600 361548
rect 69072 361508 194600 361536
rect 69072 361496 69078 361508
rect 194594 361496 194600 361508
rect 194652 361496 194658 361548
rect 123478 360816 123484 360868
rect 123536 360856 123542 360868
rect 271966 360856 271972 360868
rect 123536 360828 271972 360856
rect 123536 360816 123542 360828
rect 271966 360816 271972 360828
rect 272024 360816 272030 360868
rect 69014 360476 69020 360528
rect 69072 360516 69078 360528
rect 69750 360516 69756 360528
rect 69072 360488 69756 360516
rect 69072 360476 69078 360488
rect 69750 360476 69756 360488
rect 69808 360476 69814 360528
rect 124858 360136 124864 360188
rect 124916 360176 124922 360188
rect 245654 360176 245660 360188
rect 124916 360148 245660 360176
rect 124916 360136 124922 360148
rect 245654 360136 245660 360148
rect 245712 360136 245718 360188
rect 97258 360068 97264 360120
rect 97316 360108 97322 360120
rect 215386 360108 215392 360120
rect 97316 360080 215392 360108
rect 97316 360068 97322 360080
rect 215386 360068 215392 360080
rect 215444 360068 215450 360120
rect 215386 359660 215392 359712
rect 215444 359700 215450 359712
rect 215938 359700 215944 359712
rect 215444 359672 215944 359700
rect 215444 359660 215450 359672
rect 215938 359660 215944 359672
rect 215996 359660 216002 359712
rect 245654 359660 245660 359712
rect 245712 359700 245718 359712
rect 246298 359700 246304 359712
rect 245712 359672 246304 359700
rect 245712 359660 245718 359672
rect 246298 359660 246304 359672
rect 246356 359660 246362 359712
rect 82814 359456 82820 359508
rect 82872 359496 82878 359508
rect 103514 359496 103520 359508
rect 82872 359468 103520 359496
rect 82872 359456 82878 359468
rect 103514 359456 103520 359468
rect 103572 359456 103578 359508
rect 243538 359456 243544 359508
rect 243596 359496 243602 359508
rect 260926 359496 260932 359508
rect 243596 359468 260932 359496
rect 243596 359456 243602 359468
rect 260926 359456 260932 359468
rect 260984 359456 260990 359508
rect 104158 358708 104164 358760
rect 104216 358748 104222 358760
rect 234614 358748 234620 358760
rect 104216 358720 234620 358748
rect 104216 358708 104222 358720
rect 234614 358708 234620 358720
rect 234672 358748 234678 358760
rect 235258 358748 235264 358760
rect 234672 358720 235264 358748
rect 234672 358708 234678 358720
rect 235258 358708 235264 358720
rect 235316 358708 235322 358760
rect 3234 358640 3240 358692
rect 3292 358680 3298 358692
rect 7558 358680 7564 358692
rect 3292 358652 7564 358680
rect 3292 358640 3298 358652
rect 7558 358640 7564 358652
rect 7616 358640 7622 358692
rect 104710 357348 104716 357400
rect 104768 357388 104774 357400
rect 242802 357388 242808 357400
rect 104768 357360 242808 357388
rect 104768 357348 104774 357360
rect 242802 357348 242808 357360
rect 242860 357348 242866 357400
rect 242802 356668 242808 356720
rect 242860 356708 242866 356720
rect 254578 356708 254584 356720
rect 242860 356680 254584 356708
rect 242860 356668 242866 356680
rect 254578 356668 254584 356680
rect 254636 356668 254642 356720
rect 129090 355988 129096 356040
rect 129148 356028 129154 356040
rect 211154 356028 211160 356040
rect 129148 356000 211160 356028
rect 129148 355988 129154 356000
rect 211154 355988 211160 356000
rect 211212 356028 211218 356040
rect 211798 356028 211804 356040
rect 211212 356000 211804 356028
rect 211212 355988 211218 356000
rect 211798 355988 211804 356000
rect 211856 355988 211862 356040
rect 128998 354016 129004 354068
rect 129056 354056 129062 354068
rect 152550 354056 152556 354068
rect 129056 354028 152556 354056
rect 129056 354016 129062 354028
rect 152550 354016 152556 354028
rect 152608 354056 152614 354068
rect 216674 354056 216680 354068
rect 152608 354028 216680 354056
rect 152608 354016 152614 354028
rect 216674 354016 216680 354028
rect 216732 354016 216738 354068
rect 84194 353948 84200 354000
rect 84252 353988 84258 354000
rect 164878 353988 164884 354000
rect 84252 353960 164884 353988
rect 84252 353948 84258 353960
rect 164878 353948 164884 353960
rect 164936 353988 164942 354000
rect 214558 353988 214564 354000
rect 164936 353960 214564 353988
rect 164936 353948 164942 353960
rect 214558 353948 214564 353960
rect 214616 353948 214622 354000
rect 115382 353200 115388 353252
rect 115440 353240 115446 353252
rect 249242 353240 249248 353252
rect 115440 353212 249248 353240
rect 115440 353200 115446 353212
rect 249242 353200 249248 353212
rect 249300 353200 249306 353252
rect 218054 352520 218060 352572
rect 218112 352560 218118 352572
rect 249150 352560 249156 352572
rect 218112 352532 249156 352560
rect 218112 352520 218118 352532
rect 249150 352520 249156 352532
rect 249208 352520 249214 352572
rect 193030 351228 193036 351280
rect 193088 351268 193094 351280
rect 242986 351268 242992 351280
rect 193088 351240 242992 351268
rect 193088 351228 193094 351240
rect 242986 351228 242992 351240
rect 243044 351228 243050 351280
rect 169662 351160 169668 351212
rect 169720 351200 169726 351212
rect 178678 351200 178684 351212
rect 169720 351172 178684 351200
rect 169720 351160 169726 351172
rect 178678 351160 178684 351172
rect 178736 351160 178742 351212
rect 187418 351160 187424 351212
rect 187476 351200 187482 351212
rect 258166 351200 258172 351212
rect 187476 351172 258172 351200
rect 187476 351160 187482 351172
rect 258166 351160 258172 351172
rect 258224 351160 258230 351212
rect 169570 349800 169576 349852
rect 169628 349840 169634 349852
rect 253474 349840 253480 349852
rect 169628 349812 253480 349840
rect 169628 349800 169634 349812
rect 253474 349800 253480 349812
rect 253532 349800 253538 349852
rect 115198 349052 115204 349104
rect 115256 349092 115262 349104
rect 250530 349092 250536 349104
rect 115256 349064 250536 349092
rect 115256 349052 115262 349064
rect 250530 349052 250536 349064
rect 250588 349052 250594 349104
rect 202874 348372 202880 348424
rect 202932 348412 202938 348424
rect 252738 348412 252744 348424
rect 202932 348384 252744 348412
rect 202932 348372 202938 348384
rect 252738 348372 252744 348384
rect 252796 348372 252802 348424
rect 192846 347012 192852 347064
rect 192904 347052 192910 347064
rect 238110 347052 238116 347064
rect 192904 347024 238116 347052
rect 192904 347012 192910 347024
rect 238110 347012 238116 347024
rect 238168 347012 238174 347064
rect 177942 345652 177948 345704
rect 178000 345692 178006 345704
rect 239398 345692 239404 345704
rect 178000 345664 239404 345692
rect 178000 345652 178006 345664
rect 239398 345652 239404 345664
rect 239456 345652 239462 345704
rect 3418 345312 3424 345364
rect 3476 345352 3482 345364
rect 7558 345352 7564 345364
rect 3476 345324 7564 345352
rect 3476 345312 3482 345324
rect 7558 345312 7564 345324
rect 7616 345312 7622 345364
rect 198090 344292 198096 344344
rect 198148 344332 198154 344344
rect 250530 344332 250536 344344
rect 198148 344304 250536 344332
rect 198148 344292 198154 344304
rect 250530 344292 250536 344304
rect 250588 344292 250594 344344
rect 209774 342864 209780 342916
rect 209832 342904 209838 342916
rect 281810 342904 281816 342916
rect 209832 342876 281816 342904
rect 209832 342864 209838 342876
rect 281810 342864 281816 342876
rect 281868 342864 281874 342916
rect 247678 341572 247684 341624
rect 247736 341612 247742 341624
rect 258166 341612 258172 341624
rect 247736 341584 258172 341612
rect 247736 341572 247742 341584
rect 258166 341572 258172 341584
rect 258224 341572 258230 341624
rect 196618 341504 196624 341556
rect 196676 341544 196682 341556
rect 251910 341544 251916 341556
rect 196676 341516 251916 341544
rect 196676 341504 196682 341516
rect 251910 341504 251916 341516
rect 251968 341504 251974 341556
rect 173342 340892 173348 340944
rect 173400 340932 173406 340944
rect 244274 340932 244280 340944
rect 173400 340904 244280 340932
rect 173400 340892 173406 340904
rect 244274 340892 244280 340904
rect 244332 340892 244338 340944
rect 187510 340144 187516 340196
rect 187568 340184 187574 340196
rect 240870 340184 240876 340196
rect 187568 340156 240876 340184
rect 187568 340144 187574 340156
rect 240870 340144 240876 340156
rect 240928 340144 240934 340196
rect 92474 339464 92480 339516
rect 92532 339504 92538 339516
rect 266446 339504 266452 339516
rect 92532 339476 266452 339504
rect 92532 339464 92538 339476
rect 266446 339464 266452 339476
rect 266504 339464 266510 339516
rect 73062 338104 73068 338156
rect 73120 338144 73126 338156
rect 270678 338144 270684 338156
rect 73120 338116 270684 338144
rect 73120 338104 73126 338116
rect 270678 338104 270684 338116
rect 270736 338104 270742 338156
rect 236638 337356 236644 337408
rect 236696 337396 236702 337408
rect 262306 337396 262312 337408
rect 236696 337368 262312 337396
rect 236696 337356 236702 337368
rect 262306 337356 262312 337368
rect 262364 337356 262370 337408
rect 130470 336744 130476 336796
rect 130528 336784 130534 336796
rect 252554 336784 252560 336796
rect 130528 336756 252560 336784
rect 130528 336744 130534 336756
rect 252554 336744 252560 336756
rect 252612 336744 252618 336796
rect 169662 335996 169668 336048
rect 169720 336036 169726 336048
rect 205634 336036 205640 336048
rect 169720 336008 205640 336036
rect 169720 335996 169726 336008
rect 205634 335996 205640 336008
rect 205692 336036 205698 336048
rect 236638 336036 236644 336048
rect 205692 336008 236644 336036
rect 205692 335996 205698 336008
rect 236638 335996 236644 336008
rect 236696 335996 236702 336048
rect 137278 335316 137284 335368
rect 137336 335356 137342 335368
rect 253290 335356 253296 335368
rect 137336 335328 253296 335356
rect 137336 335316 137342 335328
rect 253290 335316 253296 335328
rect 253348 335316 253354 335368
rect 193398 334568 193404 334620
rect 193456 334608 193462 334620
rect 229094 334608 229100 334620
rect 193456 334580 229100 334608
rect 193456 334568 193462 334580
rect 229094 334568 229100 334580
rect 229152 334568 229158 334620
rect 252462 334568 252468 334620
rect 252520 334608 252526 334620
rect 260834 334608 260840 334620
rect 252520 334580 260840 334608
rect 252520 334568 252526 334580
rect 260834 334568 260840 334580
rect 260892 334568 260898 334620
rect 35802 333956 35808 334008
rect 35860 333996 35866 334008
rect 220078 333996 220084 334008
rect 35860 333968 220084 333996
rect 35860 333956 35866 333968
rect 220078 333956 220084 333968
rect 220136 333956 220142 334008
rect 223666 333208 223672 333260
rect 223724 333248 223730 333260
rect 238110 333248 238116 333260
rect 223724 333220 238116 333248
rect 223724 333208 223730 333220
rect 238110 333208 238116 333220
rect 238168 333208 238174 333260
rect 189902 332664 189908 332716
rect 189960 332704 189966 332716
rect 190362 332704 190368 332716
rect 189960 332676 190368 332704
rect 189960 332664 189966 332676
rect 190362 332664 190368 332676
rect 190420 332704 190426 332716
rect 274818 332704 274824 332716
rect 190420 332676 274824 332704
rect 190420 332664 190426 332676
rect 274818 332664 274824 332676
rect 274876 332664 274882 332716
rect 12342 332596 12348 332648
rect 12400 332636 12406 332648
rect 197354 332636 197360 332648
rect 12400 332608 197360 332636
rect 12400 332596 12406 332608
rect 197354 332596 197360 332608
rect 197412 332596 197418 332648
rect 193030 331848 193036 331900
rect 193088 331888 193094 331900
rect 233878 331888 233884 331900
rect 193088 331860 233884 331888
rect 193088 331848 193094 331860
rect 233878 331848 233884 331860
rect 233936 331848 233942 331900
rect 238018 331848 238024 331900
rect 238076 331888 238082 331900
rect 291378 331888 291384 331900
rect 238076 331860 291384 331888
rect 238076 331848 238082 331860
rect 291378 331848 291384 331860
rect 291436 331848 291442 331900
rect 138658 331236 138664 331288
rect 138716 331276 138722 331288
rect 211246 331276 211252 331288
rect 138716 331248 211252 331276
rect 138716 331236 138722 331248
rect 211246 331236 211252 331248
rect 211304 331236 211310 331288
rect 142798 329876 142804 329928
rect 142856 329916 142862 329928
rect 209038 329916 209044 329928
rect 142856 329888 209044 329916
rect 142856 329876 142862 329888
rect 209038 329876 209044 329888
rect 209096 329876 209102 329928
rect 223482 329876 223488 329928
rect 223540 329916 223546 329928
rect 259638 329916 259644 329928
rect 223540 329888 259644 329916
rect 223540 329876 223546 329888
rect 259638 329876 259644 329888
rect 259696 329876 259702 329928
rect 102870 329808 102876 329860
rect 102928 329848 102934 329860
rect 240226 329848 240232 329860
rect 102928 329820 240232 329848
rect 102928 329808 102934 329820
rect 240226 329808 240232 329820
rect 240284 329848 240290 329860
rect 240778 329848 240784 329860
rect 240284 329820 240784 329848
rect 240284 329808 240290 329820
rect 240778 329808 240784 329820
rect 240836 329808 240842 329860
rect 180150 329128 180156 329180
rect 180208 329168 180214 329180
rect 265158 329168 265164 329180
rect 180208 329140 265164 329168
rect 180208 329128 180214 329140
rect 265158 329128 265164 329140
rect 265216 329128 265222 329180
rect 128998 329060 129004 329112
rect 129056 329100 129062 329112
rect 255406 329100 255412 329112
rect 129056 329072 255412 329100
rect 129056 329060 129062 329072
rect 255406 329060 255412 329072
rect 255464 329100 255470 329112
rect 258258 329100 258264 329112
rect 255464 329072 258264 329100
rect 255464 329060 255470 329072
rect 258258 329060 258264 329072
rect 258316 329060 258322 329112
rect 226978 327700 226984 327752
rect 227036 327740 227042 327752
rect 254762 327740 254768 327752
rect 227036 327712 254768 327740
rect 227036 327700 227042 327712
rect 254762 327700 254768 327712
rect 254820 327700 254826 327752
rect 174538 327156 174544 327208
rect 174596 327196 174602 327208
rect 256694 327196 256700 327208
rect 174596 327168 256700 327196
rect 174596 327156 174602 327168
rect 256694 327156 256700 327168
rect 256752 327156 256758 327208
rect 37182 327088 37188 327140
rect 37240 327128 37246 327140
rect 204254 327128 204260 327140
rect 37240 327100 204260 327128
rect 37240 327088 37246 327100
rect 204254 327088 204260 327100
rect 204312 327088 204318 327140
rect 251818 326408 251824 326460
rect 251876 326448 251882 326460
rect 266446 326448 266452 326460
rect 251876 326420 266452 326448
rect 251876 326408 251882 326420
rect 266446 326408 266452 326420
rect 266504 326408 266510 326460
rect 68646 326340 68652 326392
rect 68704 326380 68710 326392
rect 167638 326380 167644 326392
rect 68704 326352 167644 326380
rect 68704 326340 68710 326352
rect 167638 326340 167644 326352
rect 167696 326340 167702 326392
rect 234522 326340 234528 326392
rect 234580 326380 234586 326392
rect 252002 326380 252008 326392
rect 234580 326352 252008 326380
rect 234580 326340 234586 326352
rect 252002 326340 252008 326352
rect 252060 326340 252066 326392
rect 126882 325660 126888 325712
rect 126940 325700 126946 325712
rect 250622 325700 250628 325712
rect 126940 325672 250628 325700
rect 126940 325660 126946 325672
rect 250622 325660 250628 325672
rect 250680 325660 250686 325712
rect 144270 324912 144276 324964
rect 144328 324952 144334 324964
rect 215938 324952 215944 324964
rect 144328 324924 215944 324952
rect 144328 324912 144334 324924
rect 215938 324912 215944 324924
rect 215996 324912 216002 324964
rect 228358 324912 228364 324964
rect 228416 324952 228422 324964
rect 278866 324952 278872 324964
rect 228416 324924 278872 324952
rect 228416 324912 228422 324924
rect 278866 324912 278872 324924
rect 278924 324912 278930 324964
rect 174630 324300 174636 324352
rect 174688 324340 174694 324352
rect 175182 324340 175188 324352
rect 174688 324312 175188 324340
rect 174688 324300 174694 324312
rect 175182 324300 175188 324312
rect 175240 324340 175246 324352
rect 280430 324340 280436 324352
rect 175240 324312 280436 324340
rect 175240 324300 175246 324312
rect 280430 324300 280436 324312
rect 280488 324300 280494 324352
rect 79318 323552 79324 323604
rect 79376 323592 79382 323604
rect 159358 323592 159364 323604
rect 79376 323564 159364 323592
rect 79376 323552 79382 323564
rect 159358 323552 159364 323564
rect 159416 323552 159422 323604
rect 198734 323552 198740 323604
rect 198792 323592 198798 323604
rect 255682 323592 255688 323604
rect 198792 323564 255688 323592
rect 198792 323552 198798 323564
rect 255682 323552 255688 323564
rect 255740 323552 255746 323604
rect 151170 323008 151176 323060
rect 151228 323048 151234 323060
rect 198734 323048 198740 323060
rect 151228 323020 198740 323048
rect 151228 323008 151234 323020
rect 198734 323008 198740 323020
rect 198792 323008 198798 323060
rect 161934 322940 161940 322992
rect 161992 322980 161998 322992
rect 162118 322980 162124 322992
rect 161992 322952 162124 322980
rect 161992 322940 161998 322952
rect 162118 322940 162124 322952
rect 162176 322980 162182 322992
rect 261018 322980 261024 322992
rect 162176 322952 261024 322980
rect 162176 322940 162182 322952
rect 261018 322940 261024 322952
rect 261076 322940 261082 322992
rect 116578 322192 116584 322244
rect 116636 322232 116642 322244
rect 158714 322232 158720 322244
rect 116636 322204 158720 322232
rect 116636 322192 116642 322204
rect 158714 322192 158720 322204
rect 158772 322232 158778 322244
rect 263870 322232 263876 322244
rect 158772 322204 263876 322232
rect 158772 322192 158778 322204
rect 263870 322192 263876 322204
rect 263928 322192 263934 322244
rect 107562 322124 107568 322176
rect 107620 322164 107626 322176
rect 115290 322164 115296 322176
rect 107620 322136 115296 322164
rect 107620 322124 107626 322136
rect 115290 322124 115296 322136
rect 115348 322124 115354 322176
rect 141510 321580 141516 321632
rect 141568 321620 141574 321632
rect 142062 321620 142068 321632
rect 141568 321592 142068 321620
rect 141568 321580 141574 321592
rect 142062 321580 142068 321592
rect 142120 321620 142126 321632
rect 265250 321620 265256 321632
rect 142120 321592 265256 321620
rect 142120 321580 142126 321592
rect 265250 321580 265256 321592
rect 265308 321580 265314 321632
rect 116026 321512 116032 321564
rect 116084 321552 116090 321564
rect 276106 321552 276112 321564
rect 116084 321524 276112 321552
rect 116084 321512 116090 321524
rect 276106 321512 276112 321524
rect 276164 321512 276170 321564
rect 104158 320832 104164 320884
rect 104216 320872 104222 320884
rect 137278 320872 137284 320884
rect 104216 320844 137284 320872
rect 104216 320832 104222 320844
rect 137278 320832 137284 320844
rect 137336 320832 137342 320884
rect 97994 320152 98000 320204
rect 98052 320192 98058 320204
rect 98052 320164 113174 320192
rect 98052 320152 98058 320164
rect 113146 320124 113174 320164
rect 180150 320152 180156 320204
rect 180208 320192 180214 320204
rect 270494 320192 270500 320204
rect 180208 320164 270500 320192
rect 180208 320152 180214 320164
rect 270494 320152 270500 320164
rect 270552 320152 270558 320204
rect 142890 320124 142896 320136
rect 113146 320096 142896 320124
rect 142890 320084 142896 320096
rect 142948 320124 142954 320136
rect 143442 320124 143448 320136
rect 142948 320096 143448 320124
rect 142948 320084 142954 320096
rect 143442 320084 143448 320096
rect 143500 320084 143506 320136
rect 100754 320016 100760 320068
rect 100812 320056 100818 320068
rect 102686 320056 102692 320068
rect 100812 320028 102692 320056
rect 100812 320016 100818 320028
rect 102686 320016 102692 320028
rect 102744 320056 102750 320068
rect 126882 320056 126888 320068
rect 102744 320028 126888 320056
rect 102744 320016 102750 320028
rect 126882 320016 126888 320028
rect 126940 320056 126946 320068
rect 127618 320056 127624 320068
rect 126940 320028 127624 320056
rect 126940 320016 126946 320028
rect 127618 320016 127624 320028
rect 127676 320016 127682 320068
rect 4062 319404 4068 319456
rect 4120 319444 4126 319456
rect 17218 319444 17224 319456
rect 4120 319416 17224 319444
rect 4120 319404 4126 319416
rect 17218 319404 17224 319416
rect 17276 319404 17282 319456
rect 143442 319404 143448 319456
rect 143500 319444 143506 319456
rect 211798 319444 211804 319456
rect 143500 319416 211804 319444
rect 143500 319404 143506 319416
rect 211798 319404 211804 319416
rect 211856 319404 211862 319456
rect 231118 319404 231124 319456
rect 231176 319444 231182 319456
rect 272518 319444 272524 319456
rect 231176 319416 272524 319444
rect 231176 319404 231182 319416
rect 272518 319404 272524 319416
rect 272576 319404 272582 319456
rect 178770 318792 178776 318844
rect 178828 318832 178834 318844
rect 179230 318832 179236 318844
rect 178828 318804 179236 318832
rect 178828 318792 178834 318804
rect 179230 318792 179236 318804
rect 179288 318832 179294 318844
rect 229738 318832 229744 318844
rect 179288 318804 229744 318832
rect 179288 318792 179294 318804
rect 229738 318792 229744 318804
rect 229796 318792 229802 318844
rect 265066 318724 265072 318776
rect 265124 318764 265130 318776
rect 265342 318764 265348 318776
rect 265124 318736 265348 318764
rect 265124 318724 265130 318736
rect 265342 318724 265348 318736
rect 265400 318724 265406 318776
rect 183002 317500 183008 317552
rect 183060 317540 183066 317552
rect 265342 317540 265348 317552
rect 183060 317512 265348 317540
rect 183060 317500 183066 317512
rect 265342 317500 265348 317512
rect 265400 317500 265406 317552
rect 82722 317432 82728 317484
rect 82780 317472 82786 317484
rect 233878 317472 233884 317484
rect 82780 317444 233884 317472
rect 82780 317432 82786 317444
rect 233878 317432 233884 317444
rect 233936 317432 233942 317484
rect 101582 316684 101588 316736
rect 101640 316724 101646 316736
rect 113266 316724 113272 316736
rect 101640 316696 113272 316724
rect 101640 316684 101646 316696
rect 113266 316684 113272 316696
rect 113324 316684 113330 316736
rect 135990 316684 135996 316736
rect 136048 316724 136054 316736
rect 259454 316724 259460 316736
rect 136048 316696 259460 316724
rect 136048 316684 136054 316696
rect 259454 316684 259460 316696
rect 259512 316684 259518 316736
rect 177850 316004 177856 316056
rect 177908 316044 177914 316056
rect 277578 316044 277584 316056
rect 177908 316016 277584 316044
rect 177908 316004 177914 316016
rect 277578 316004 277584 316016
rect 277636 316004 277642 316056
rect 229738 315256 229744 315308
rect 229796 315296 229802 315308
rect 256878 315296 256884 315308
rect 229796 315268 256884 315296
rect 229796 315256 229802 315268
rect 256878 315256 256884 315268
rect 256936 315256 256942 315308
rect 153838 314712 153844 314764
rect 153896 314752 153902 314764
rect 214282 314752 214288 314764
rect 153896 314724 214288 314752
rect 153896 314712 153902 314724
rect 214282 314712 214288 314724
rect 214340 314712 214346 314764
rect 67450 314644 67456 314696
rect 67508 314684 67514 314696
rect 268010 314684 268016 314696
rect 67508 314656 268016 314684
rect 67508 314644 67514 314656
rect 268010 314644 268016 314656
rect 268068 314644 268074 314696
rect 250530 314032 250536 314084
rect 250588 314072 250594 314084
rect 256970 314072 256976 314084
rect 250588 314044 256976 314072
rect 250588 314032 250594 314044
rect 256970 314032 256976 314044
rect 257028 314032 257034 314084
rect 171962 313352 171968 313404
rect 172020 313392 172026 313404
rect 174538 313392 174544 313404
rect 172020 313364 174544 313392
rect 172020 313352 172026 313364
rect 174538 313352 174544 313364
rect 174596 313352 174602 313404
rect 192478 313352 192484 313404
rect 192536 313392 192542 313404
rect 200114 313392 200120 313404
rect 192536 313364 200120 313392
rect 192536 313352 192542 313364
rect 200114 313352 200120 313364
rect 200172 313392 200178 313404
rect 201402 313392 201408 313404
rect 200172 313364 201408 313392
rect 200172 313352 200178 313364
rect 201402 313352 201408 313364
rect 201460 313352 201466 313404
rect 87598 313284 87604 313336
rect 87656 313324 87662 313336
rect 88242 313324 88248 313336
rect 87656 313296 88248 313324
rect 87656 313284 87662 313296
rect 88242 313284 88248 313296
rect 88300 313324 88306 313336
rect 266538 313324 266544 313336
rect 88300 313296 266544 313324
rect 88300 313284 88306 313296
rect 266538 313284 266544 313296
rect 266596 313284 266602 313336
rect 167730 311924 167736 311976
rect 167788 311964 167794 311976
rect 168282 311964 168288 311976
rect 167788 311936 168288 311964
rect 167788 311924 167794 311936
rect 168282 311924 168288 311936
rect 168340 311964 168346 311976
rect 226978 311964 226984 311976
rect 168340 311936 226984 311964
rect 168340 311924 168346 311936
rect 226978 311924 226984 311936
rect 227036 311924 227042 311976
rect 244550 311924 244556 311976
rect 244608 311964 244614 311976
rect 244918 311964 244924 311976
rect 244608 311936 244924 311964
rect 244608 311924 244614 311936
rect 244918 311924 244924 311936
rect 244976 311964 244982 311976
rect 262398 311964 262404 311976
rect 244976 311936 262404 311964
rect 244976 311924 244982 311936
rect 262398 311924 262404 311936
rect 262456 311924 262462 311976
rect 181530 311856 181536 311908
rect 181588 311896 181594 311908
rect 278958 311896 278964 311908
rect 181588 311868 278964 311896
rect 181588 311856 181594 311868
rect 278958 311856 278964 311868
rect 279016 311856 279022 311908
rect 193306 311108 193312 311160
rect 193364 311148 193370 311160
rect 205726 311148 205732 311160
rect 193364 311120 205732 311148
rect 193364 311108 193370 311120
rect 205726 311108 205732 311120
rect 205784 311108 205790 311160
rect 281442 311108 281448 311160
rect 281500 311148 281506 311160
rect 580258 311148 580264 311160
rect 281500 311120 580264 311148
rect 281500 311108 281506 311120
rect 580258 311108 580264 311120
rect 580316 311108 580322 311160
rect 266354 310972 266360 311024
rect 266412 311012 266418 311024
rect 266630 311012 266636 311024
rect 266412 310984 266636 311012
rect 266412 310972 266418 310984
rect 266630 310972 266636 310984
rect 266688 310972 266694 311024
rect 210418 310564 210424 310616
rect 210476 310604 210482 310616
rect 255406 310604 255412 310616
rect 210476 310576 255412 310604
rect 210476 310564 210482 310576
rect 255406 310564 255412 310576
rect 255464 310564 255470 310616
rect 174538 310496 174544 310548
rect 174596 310536 174602 310548
rect 266630 310536 266636 310548
rect 174596 310508 266636 310536
rect 174596 310496 174602 310508
rect 266630 310496 266636 310508
rect 266688 310496 266694 310548
rect 201402 309816 201408 309868
rect 201460 309856 201466 309868
rect 232498 309856 232504 309868
rect 201460 309828 232504 309856
rect 201460 309816 201466 309828
rect 232498 309816 232504 309828
rect 232556 309816 232562 309868
rect 41322 309748 41328 309800
rect 41380 309788 41386 309800
rect 172606 309788 172612 309800
rect 41380 309760 172612 309788
rect 41380 309748 41386 309760
rect 172606 309748 172612 309760
rect 172664 309788 172670 309800
rect 173158 309788 173164 309800
rect 172664 309760 173164 309788
rect 172664 309748 172670 309760
rect 173158 309748 173164 309760
rect 173216 309748 173222 309800
rect 223574 309748 223580 309800
rect 223632 309788 223638 309800
rect 255498 309788 255504 309800
rect 223632 309760 255504 309788
rect 223632 309748 223638 309760
rect 255498 309748 255504 309760
rect 255556 309748 255562 309800
rect 262858 309748 262864 309800
rect 262916 309788 262922 309800
rect 264974 309788 264980 309800
rect 262916 309760 264980 309788
rect 262916 309748 262922 309760
rect 264974 309748 264980 309760
rect 265032 309788 265038 309800
rect 287330 309788 287336 309800
rect 265032 309760 287336 309788
rect 265032 309748 265038 309760
rect 287330 309748 287336 309760
rect 287388 309748 287394 309800
rect 155218 309136 155224 309188
rect 155276 309176 155282 309188
rect 217410 309176 217416 309188
rect 155276 309148 217416 309176
rect 155276 309136 155282 309148
rect 217410 309136 217416 309148
rect 217468 309136 217474 309188
rect 240134 308456 240140 308508
rect 240192 308496 240198 308508
rect 258350 308496 258356 308508
rect 240192 308468 258356 308496
rect 240192 308456 240198 308468
rect 258350 308456 258356 308468
rect 258408 308456 258414 308508
rect 230474 308388 230480 308440
rect 230532 308428 230538 308440
rect 255590 308428 255596 308440
rect 230532 308400 255596 308428
rect 230532 308388 230538 308400
rect 255590 308388 255596 308400
rect 255648 308388 255654 308440
rect 171134 307844 171140 307896
rect 171192 307884 171198 307896
rect 215294 307884 215300 307896
rect 171192 307856 215300 307884
rect 171192 307844 171198 307856
rect 215294 307844 215300 307856
rect 215352 307844 215358 307896
rect 151078 307776 151084 307828
rect 151136 307816 151142 307828
rect 219710 307816 219716 307828
rect 151136 307788 219716 307816
rect 151136 307776 151142 307788
rect 219710 307776 219716 307788
rect 219768 307776 219774 307828
rect 220078 307708 220084 307760
rect 220136 307748 220142 307760
rect 224770 307748 224776 307760
rect 220136 307720 224776 307748
rect 220136 307708 220142 307720
rect 224770 307708 224776 307720
rect 224828 307708 224834 307760
rect 63402 307028 63408 307080
rect 63460 307068 63466 307080
rect 116578 307068 116584 307080
rect 63460 307040 116584 307068
rect 63460 307028 63466 307040
rect 116578 307028 116584 307040
rect 116636 307028 116642 307080
rect 236638 307028 236644 307080
rect 236696 307068 236702 307080
rect 241790 307068 241796 307080
rect 236696 307040 241796 307068
rect 236696 307028 236702 307040
rect 241790 307028 241796 307040
rect 241848 307028 241854 307080
rect 244458 307028 244464 307080
rect 244516 307068 244522 307080
rect 262214 307068 262220 307080
rect 244516 307040 262220 307068
rect 244516 307028 244522 307040
rect 262214 307028 262220 307040
rect 262272 307028 262278 307080
rect 148318 306416 148324 306468
rect 148376 306456 148382 306468
rect 215938 306456 215944 306468
rect 148376 306428 215944 306456
rect 148376 306416 148382 306428
rect 215938 306416 215944 306428
rect 215996 306416 216002 306468
rect 117222 306348 117228 306400
rect 117280 306388 117286 306400
rect 239306 306388 239312 306400
rect 117280 306360 239312 306388
rect 117280 306348 117286 306360
rect 239306 306348 239312 306360
rect 239364 306348 239370 306400
rect 242158 306348 242164 306400
rect 242216 306388 242222 306400
rect 276290 306388 276296 306400
rect 242216 306360 276296 306388
rect 242216 306348 242222 306360
rect 276290 306348 276296 306360
rect 276348 306348 276354 306400
rect 226978 305600 226984 305652
rect 227036 305640 227042 305652
rect 259454 305640 259460 305652
rect 227036 305612 259460 305640
rect 227036 305600 227042 305612
rect 259454 305600 259460 305612
rect 259512 305600 259518 305652
rect 141418 305056 141424 305108
rect 141476 305096 141482 305108
rect 216582 305096 216588 305108
rect 141476 305068 216588 305096
rect 141476 305056 141482 305068
rect 216582 305056 216588 305068
rect 216640 305056 216646 305108
rect 3234 304988 3240 305040
rect 3292 305028 3298 305040
rect 18598 305028 18604 305040
rect 3292 305000 18604 305028
rect 3292 304988 3298 305000
rect 18598 304988 18604 305000
rect 18656 304988 18662 305040
rect 77294 304988 77300 305040
rect 77352 305028 77358 305040
rect 86218 305028 86224 305040
rect 77352 305000 86224 305028
rect 77352 304988 77358 305000
rect 86218 304988 86224 305000
rect 86276 304988 86282 305040
rect 142890 304988 142896 305040
rect 142948 305028 142954 305040
rect 219066 305028 219072 305040
rect 142948 305000 219072 305028
rect 142948 304988 142954 305000
rect 219066 304988 219072 305000
rect 219124 304988 219130 305040
rect 250622 304988 250628 305040
rect 250680 305028 250686 305040
rect 252922 305028 252928 305040
rect 250680 305000 252928 305028
rect 250680 304988 250686 305000
rect 252922 304988 252928 305000
rect 252980 304988 252986 305040
rect 209038 304512 209044 304564
rect 209096 304552 209102 304564
rect 212166 304552 212172 304564
rect 209096 304524 212172 304552
rect 209096 304512 209102 304524
rect 212166 304512 212172 304524
rect 212224 304512 212230 304564
rect 86770 304308 86776 304360
rect 86828 304348 86834 304360
rect 95326 304348 95332 304360
rect 86828 304320 95332 304348
rect 86828 304308 86834 304320
rect 95326 304308 95332 304320
rect 95384 304308 95390 304360
rect 130378 304308 130384 304360
rect 130436 304348 130442 304360
rect 171134 304348 171140 304360
rect 130436 304320 171140 304348
rect 130436 304308 130442 304320
rect 171134 304308 171140 304320
rect 171192 304308 171198 304360
rect 232498 304308 232504 304360
rect 232556 304348 232562 304360
rect 252646 304348 252652 304360
rect 232556 304320 252652 304348
rect 232556 304308 232562 304320
rect 252646 304308 252652 304320
rect 252704 304308 252710 304360
rect 253198 304308 253204 304360
rect 253256 304348 253262 304360
rect 262858 304348 262864 304360
rect 253256 304320 262864 304348
rect 253256 304308 253262 304320
rect 262858 304308 262864 304320
rect 262916 304308 262922 304360
rect 60550 304240 60556 304292
rect 60608 304280 60614 304292
rect 181530 304280 181536 304292
rect 60608 304252 181536 304280
rect 60608 304240 60614 304252
rect 181530 304240 181536 304252
rect 181588 304240 181594 304292
rect 247494 304240 247500 304292
rect 247552 304280 247558 304292
rect 252462 304280 252468 304292
rect 247552 304252 252468 304280
rect 247552 304240 247558 304252
rect 252462 304240 252468 304252
rect 252520 304280 252526 304292
rect 295426 304280 295432 304292
rect 252520 304252 295432 304280
rect 252520 304240 252526 304252
rect 295426 304240 295432 304252
rect 295484 304240 295490 304292
rect 108850 303968 108856 304020
rect 108908 304008 108914 304020
rect 115382 304008 115388 304020
rect 108908 303980 115388 304008
rect 108908 303968 108914 303980
rect 115382 303968 115388 303980
rect 115440 303968 115446 304020
rect 182818 303764 182824 303816
rect 182876 303804 182882 303816
rect 231026 303804 231032 303816
rect 182876 303776 231032 303804
rect 182876 303764 182882 303776
rect 231026 303764 231032 303776
rect 231084 303764 231090 303816
rect 189810 303696 189816 303748
rect 189868 303736 189874 303748
rect 196342 303736 196348 303748
rect 189868 303708 196348 303736
rect 189868 303696 189874 303708
rect 196342 303696 196348 303708
rect 196400 303696 196406 303748
rect 197354 303628 197360 303680
rect 197412 303668 197418 303680
rect 197998 303668 198004 303680
rect 197412 303640 198004 303668
rect 197412 303628 197418 303640
rect 197998 303628 198004 303640
rect 198056 303628 198062 303680
rect 200206 303628 200212 303680
rect 200264 303668 200270 303680
rect 201126 303668 201132 303680
rect 200264 303640 201132 303668
rect 200264 303628 200270 303640
rect 201126 303628 201132 303640
rect 201184 303628 201190 303680
rect 230106 303628 230112 303680
rect 230164 303668 230170 303680
rect 238662 303668 238668 303680
rect 230164 303640 238668 303668
rect 230164 303628 230170 303640
rect 238662 303628 238668 303640
rect 238720 303628 238726 303680
rect 244274 303628 244280 303680
rect 244332 303668 244338 303680
rect 244550 303668 244556 303680
rect 244332 303640 244556 303668
rect 244332 303628 244338 303640
rect 244550 303628 244556 303640
rect 244608 303628 244614 303680
rect 201402 303560 201408 303612
rect 201460 303600 201466 303612
rect 210418 303600 210424 303612
rect 201460 303572 210424 303600
rect 201460 303560 201466 303572
rect 210418 303560 210424 303572
rect 210476 303560 210482 303612
rect 153102 302880 153108 302932
rect 153160 302920 153166 302932
rect 192478 302920 192484 302932
rect 153160 302892 192484 302920
rect 153160 302880 153166 302892
rect 192478 302880 192484 302892
rect 192536 302880 192542 302932
rect 192754 302268 192760 302320
rect 192812 302308 192818 302320
rect 198826 302308 198832 302320
rect 192812 302280 198832 302308
rect 192812 302268 192818 302280
rect 198826 302268 198832 302280
rect 198884 302268 198890 302320
rect 250622 302268 250628 302320
rect 250680 302308 250686 302320
rect 260834 302308 260840 302320
rect 250680 302280 260840 302308
rect 250680 302268 250686 302280
rect 260834 302268 260840 302280
rect 260892 302268 260898 302320
rect 115290 302200 115296 302252
rect 115348 302240 115354 302252
rect 118786 302240 118792 302252
rect 115348 302212 118792 302240
rect 115348 302200 115354 302212
rect 118786 302200 118792 302212
rect 118844 302200 118850 302252
rect 180242 302200 180248 302252
rect 180300 302240 180306 302252
rect 218422 302240 218428 302252
rect 180300 302212 218428 302240
rect 180300 302200 180306 302212
rect 218422 302200 218428 302212
rect 218480 302200 218486 302252
rect 252002 302200 252008 302252
rect 252060 302240 252066 302252
rect 253014 302240 253020 302252
rect 252060 302212 253020 302240
rect 252060 302200 252066 302212
rect 253014 302200 253020 302212
rect 253072 302200 253078 302252
rect 241054 302132 241060 302184
rect 241112 302172 241118 302184
rect 253658 302172 253664 302184
rect 241112 302144 253664 302172
rect 241112 302132 241118 302144
rect 253658 302132 253664 302144
rect 253716 302132 253722 302184
rect 253290 301520 253296 301572
rect 253348 301560 253354 301572
rect 254118 301560 254124 301572
rect 253348 301532 254124 301560
rect 253348 301520 253354 301532
rect 254118 301520 254124 301532
rect 254176 301520 254182 301572
rect 91186 301452 91192 301504
rect 91244 301492 91250 301504
rect 135990 301492 135996 301504
rect 91244 301464 135996 301492
rect 91244 301452 91250 301464
rect 135990 301452 135996 301464
rect 136048 301452 136054 301504
rect 191466 301452 191472 301504
rect 191524 301492 191530 301504
rect 191742 301492 191748 301504
rect 191524 301464 191748 301492
rect 191524 301452 191530 301464
rect 191742 301452 191748 301464
rect 191800 301452 191806 301504
rect 191742 301316 191748 301368
rect 191800 301356 191806 301368
rect 196710 301356 196716 301368
rect 191800 301328 196716 301356
rect 191800 301316 191806 301328
rect 196710 301316 196716 301328
rect 196768 301316 196774 301368
rect 240134 301356 240140 301368
rect 219406 301328 240140 301356
rect 191098 301016 191104 301028
rect 180766 300988 191104 301016
rect 175918 300908 175924 300960
rect 175976 300948 175982 300960
rect 180766 300948 180794 300988
rect 191098 300976 191104 300988
rect 191156 300976 191162 301028
rect 175976 300920 180794 300948
rect 175976 300908 175982 300920
rect 159450 300840 159456 300892
rect 159508 300880 159514 300892
rect 219406 300880 219434 301328
rect 240134 301316 240140 301328
rect 240192 301316 240198 301368
rect 246482 301316 246488 301368
rect 246540 301316 246546 301368
rect 249150 301316 249156 301368
rect 249208 301356 249214 301368
rect 253106 301356 253112 301368
rect 249208 301328 253112 301356
rect 249208 301316 249214 301328
rect 253106 301316 253112 301328
rect 253164 301316 253170 301368
rect 159508 300852 219434 300880
rect 159508 300840 159514 300852
rect 178034 300772 178040 300824
rect 178092 300812 178098 300824
rect 178770 300812 178776 300824
rect 178092 300784 178776 300812
rect 178092 300772 178098 300784
rect 178770 300772 178776 300784
rect 178828 300772 178834 300824
rect 192202 300772 192208 300824
rect 192260 300812 192266 300824
rect 195054 300812 195060 300824
rect 192260 300784 195060 300812
rect 192260 300772 192266 300784
rect 195054 300772 195060 300784
rect 195112 300772 195118 300824
rect 206462 300812 206468 300824
rect 200086 300784 206468 300812
rect 93946 300160 93952 300212
rect 94004 300200 94010 300212
rect 95050 300200 95056 300212
rect 94004 300172 95056 300200
rect 94004 300160 94010 300172
rect 95050 300160 95056 300172
rect 95108 300160 95114 300212
rect 186958 299888 186964 299940
rect 187016 299928 187022 299940
rect 187602 299928 187608 299940
rect 187016 299900 187608 299928
rect 187016 299888 187022 299900
rect 187602 299888 187608 299900
rect 187660 299928 187666 299940
rect 191742 299928 191748 299940
rect 187660 299900 191748 299928
rect 187660 299888 187666 299900
rect 191742 299888 191748 299900
rect 191800 299888 191806 299940
rect 77938 299548 77944 299600
rect 77996 299588 78002 299600
rect 178034 299588 178040 299600
rect 77996 299560 178040 299588
rect 77996 299548 78002 299560
rect 178034 299548 178040 299560
rect 178092 299548 178098 299600
rect 95050 299480 95056 299532
rect 95108 299520 95114 299532
rect 147030 299520 147036 299532
rect 95108 299492 147036 299520
rect 95108 299480 95114 299492
rect 147030 299480 147036 299492
rect 147088 299480 147094 299532
rect 149790 299480 149796 299532
rect 149848 299520 149854 299532
rect 200086 299520 200114 300784
rect 206462 300772 206468 300784
rect 206520 300772 206526 300824
rect 246500 300812 246528 301316
rect 252830 300812 252836 300824
rect 246500 300784 252836 300812
rect 252830 300772 252836 300784
rect 252888 300772 252894 300824
rect 256602 299548 256608 299600
rect 256660 299588 256666 299600
rect 288526 299588 288532 299600
rect 256660 299560 288532 299588
rect 256660 299548 256666 299560
rect 288526 299548 288532 299560
rect 288584 299548 288590 299600
rect 149848 299492 200114 299520
rect 149848 299480 149854 299492
rect 256510 299480 256516 299532
rect 256568 299520 256574 299532
rect 289814 299520 289820 299532
rect 256568 299492 289820 299520
rect 256568 299480 256574 299492
rect 289814 299480 289820 299492
rect 289872 299480 289878 299532
rect 105630 299412 105636 299464
rect 105688 299452 105694 299464
rect 107562 299452 107568 299464
rect 105688 299424 107568 299452
rect 105688 299412 105694 299424
rect 107562 299412 107568 299424
rect 107620 299452 107626 299464
rect 190638 299452 190644 299464
rect 107620 299424 190644 299452
rect 107620 299412 107626 299424
rect 190638 299412 190644 299424
rect 190696 299412 190702 299464
rect 272518 299412 272524 299464
rect 272576 299452 272582 299464
rect 580166 299452 580172 299464
rect 272576 299424 580172 299452
rect 272576 299412 272582 299424
rect 580166 299412 580172 299424
rect 580224 299412 580230 299464
rect 67542 298732 67548 298784
rect 67600 298772 67606 298784
rect 167638 298772 167644 298784
rect 67600 298744 167644 298772
rect 67600 298732 67606 298744
rect 167638 298732 167644 298744
rect 167696 298732 167702 298784
rect 253106 298188 253112 298240
rect 253164 298228 253170 298240
rect 262398 298228 262404 298240
rect 253164 298200 262404 298228
rect 253164 298188 253170 298200
rect 262398 298188 262404 298200
rect 262456 298188 262462 298240
rect 256602 298120 256608 298172
rect 256660 298160 256666 298172
rect 285766 298160 285772 298172
rect 256660 298132 285772 298160
rect 256660 298120 256666 298132
rect 285766 298120 285772 298132
rect 285824 298120 285830 298172
rect 255866 297440 255872 297492
rect 255924 297480 255930 297492
rect 266354 297480 266360 297492
rect 255924 297452 266360 297480
rect 255924 297440 255930 297452
rect 266354 297440 266360 297452
rect 266412 297440 266418 297492
rect 256510 297372 256516 297424
rect 256568 297412 256574 297424
rect 259546 297412 259552 297424
rect 256568 297384 259552 297412
rect 256568 297372 256574 297384
rect 259546 297372 259552 297384
rect 259604 297412 259610 297424
rect 287238 297412 287244 297424
rect 259604 297384 287244 297412
rect 259604 297372 259610 297384
rect 287238 297372 287244 297384
rect 287296 297372 287302 297424
rect 119338 296692 119344 296744
rect 119396 296732 119402 296744
rect 191742 296732 191748 296744
rect 119396 296704 191748 296732
rect 119396 296692 119402 296704
rect 191742 296692 191748 296704
rect 191800 296692 191806 296744
rect 259362 296624 259368 296676
rect 259420 296664 259426 296676
rect 262490 296664 262496 296676
rect 259420 296636 262496 296664
rect 259420 296624 259426 296636
rect 262490 296624 262496 296636
rect 262548 296624 262554 296676
rect 76006 295944 76012 295996
rect 76064 295984 76070 295996
rect 174630 295984 174636 295996
rect 76064 295956 174636 295984
rect 76064 295944 76070 295956
rect 174630 295944 174636 295956
rect 174688 295944 174694 295996
rect 256602 295944 256608 295996
rect 256660 295984 256666 295996
rect 258258 295984 258264 295996
rect 256660 295956 258264 295984
rect 256660 295944 256666 295956
rect 258258 295944 258264 295956
rect 258316 295984 258322 295996
rect 276382 295984 276388 295996
rect 258316 295956 276388 295984
rect 258316 295944 258322 295956
rect 276382 295944 276388 295956
rect 276440 295944 276446 295996
rect 128354 295332 128360 295384
rect 128412 295372 128418 295384
rect 187602 295372 187608 295384
rect 128412 295344 187608 295372
rect 128412 295332 128418 295344
rect 187602 295332 187608 295344
rect 187660 295372 187666 295384
rect 193030 295372 193036 295384
rect 187660 295344 193036 295372
rect 187660 295332 187666 295344
rect 193030 295332 193036 295344
rect 193088 295332 193094 295384
rect 256602 294992 256608 295044
rect 256660 295032 256666 295044
rect 262490 295032 262496 295044
rect 256660 295004 262496 295032
rect 256660 294992 256666 295004
rect 262490 294992 262496 295004
rect 262548 294992 262554 295044
rect 96614 294584 96620 294636
rect 96672 294624 96678 294636
rect 129090 294624 129096 294636
rect 96672 294596 129096 294624
rect 96672 294584 96678 294596
rect 129090 294584 129096 294596
rect 129148 294584 129154 294636
rect 140130 294584 140136 294636
rect 140188 294624 140194 294636
rect 186958 294624 186964 294636
rect 140188 294596 186964 294624
rect 140188 294584 140194 294596
rect 186958 294584 186964 294596
rect 187016 294584 187022 294636
rect 258074 294584 258080 294636
rect 258132 294624 258138 294636
rect 258258 294624 258264 294636
rect 258132 294596 258264 294624
rect 258132 294584 258138 294596
rect 258258 294584 258264 294596
rect 258316 294584 258322 294636
rect 184842 294108 184848 294160
rect 184900 294148 184906 294160
rect 191742 294148 191748 294160
rect 184900 294120 191748 294148
rect 184900 294108 184906 294120
rect 191742 294108 191748 294120
rect 191800 294108 191806 294160
rect 102962 294040 102968 294092
rect 103020 294080 103026 294092
rect 104158 294080 104164 294092
rect 103020 294052 104164 294080
rect 103020 294040 103026 294052
rect 104158 294040 104164 294052
rect 104216 294040 104222 294092
rect 256602 293972 256608 294024
rect 256660 294012 256666 294024
rect 269114 294012 269120 294024
rect 256660 293984 269120 294012
rect 256660 293972 256666 293984
rect 269114 293972 269120 293984
rect 269172 293972 269178 294024
rect 102134 293904 102140 293956
rect 102192 293944 102198 293956
rect 102778 293944 102784 293956
rect 102192 293916 102784 293944
rect 102192 293904 102198 293916
rect 102778 293904 102784 293916
rect 102836 293944 102842 293956
rect 128354 293944 128360 293956
rect 102836 293916 128360 293944
rect 102836 293904 102842 293916
rect 128354 293904 128360 293916
rect 128412 293904 128418 293956
rect 93118 293292 93124 293344
rect 93176 293332 93182 293344
rect 102134 293332 102140 293344
rect 93176 293304 102140 293332
rect 93176 293292 93182 293304
rect 102134 293292 102140 293304
rect 102192 293292 102198 293344
rect 84194 293224 84200 293276
rect 84252 293264 84258 293276
rect 177298 293264 177304 293276
rect 84252 293236 177304 293264
rect 84252 293224 84258 293236
rect 177298 293224 177304 293236
rect 177356 293224 177362 293276
rect 262398 293224 262404 293276
rect 262456 293264 262462 293276
rect 281534 293264 281540 293276
rect 262456 293236 281540 293264
rect 262456 293224 262462 293236
rect 281534 293224 281540 293236
rect 281592 293224 281598 293276
rect 256602 292884 256608 292936
rect 256660 292924 256666 292936
rect 259638 292924 259644 292936
rect 256660 292896 259644 292924
rect 256660 292884 256666 292896
rect 259638 292884 259644 292896
rect 259696 292924 259702 292936
rect 260742 292924 260748 292936
rect 259696 292896 260748 292924
rect 259696 292884 259702 292896
rect 260742 292884 260748 292896
rect 260800 292884 260806 292936
rect 187418 292584 187424 292596
rect 186332 292556 187424 292584
rect 99282 292476 99288 292528
rect 99340 292516 99346 292528
rect 186332 292516 186360 292556
rect 187418 292544 187424 292556
rect 187476 292584 187482 292596
rect 191742 292584 191748 292596
rect 187476 292556 191748 292584
rect 187476 292544 187482 292556
rect 191742 292544 191748 292556
rect 191800 292544 191806 292596
rect 99340 292488 186360 292516
rect 99340 292476 99346 292488
rect 255406 292204 255412 292256
rect 255464 292244 255470 292256
rect 259362 292244 259368 292256
rect 255464 292216 259368 292244
rect 255464 292204 255470 292216
rect 259362 292204 259368 292216
rect 259420 292204 259426 292256
rect 264882 291864 264888 291916
rect 264940 291904 264946 291916
rect 280798 291904 280804 291916
rect 264940 291876 280804 291904
rect 264940 291864 264946 291876
rect 280798 291864 280804 291876
rect 280856 291904 280862 291916
rect 291194 291904 291200 291916
rect 280856 291876 291200 291904
rect 280856 291864 280862 291876
rect 291194 291864 291200 291876
rect 291252 291864 291258 291916
rect 53650 291796 53656 291848
rect 53708 291836 53714 291848
rect 53708 291808 161474 291836
rect 53708 291796 53714 291808
rect 161446 291768 161474 291808
rect 183462 291796 183468 291848
rect 183520 291836 183526 291848
rect 191742 291836 191748 291848
rect 183520 291808 191748 291836
rect 183520 291796 183526 291808
rect 191742 291796 191748 291808
rect 191800 291796 191806 291848
rect 260742 291796 260748 291848
rect 260800 291836 260806 291848
rect 291470 291836 291476 291848
rect 260800 291808 291476 291836
rect 260800 291796 260806 291808
rect 291470 291796 291476 291808
rect 291528 291796 291534 291848
rect 182910 291768 182916 291780
rect 161446 291740 182916 291768
rect 182910 291728 182916 291740
rect 182968 291728 182974 291780
rect 72418 291184 72424 291236
rect 72476 291224 72482 291236
rect 76006 291224 76012 291236
rect 72476 291196 76012 291224
rect 72476 291184 72482 291196
rect 76006 291184 76012 291196
rect 76064 291184 76070 291236
rect 98454 291184 98460 291236
rect 98512 291224 98518 291236
rect 99282 291224 99288 291236
rect 98512 291196 99288 291224
rect 98512 291184 98518 291196
rect 99282 291184 99288 291196
rect 99340 291184 99346 291236
rect 255406 290504 255412 290556
rect 255464 290544 255470 290556
rect 258442 290544 258448 290556
rect 255464 290516 258448 290544
rect 255464 290504 255470 290516
rect 258442 290504 258448 290516
rect 258500 290544 258506 290556
rect 262582 290544 262588 290556
rect 258500 290516 262588 290544
rect 258500 290504 258506 290516
rect 262582 290504 262588 290516
rect 262640 290504 262646 290556
rect 39850 290436 39856 290488
rect 39908 290476 39914 290488
rect 61746 290476 61752 290488
rect 39908 290448 61752 290476
rect 39908 290436 39914 290448
rect 61746 290436 61752 290448
rect 61804 290476 61810 290488
rect 73246 290476 73252 290488
rect 61804 290448 73252 290476
rect 61804 290436 61810 290448
rect 73246 290436 73252 290448
rect 73304 290436 73310 290488
rect 77018 290436 77024 290488
rect 77076 290476 77082 290488
rect 84838 290476 84844 290488
rect 77076 290448 84844 290476
rect 77076 290436 77082 290448
rect 84838 290436 84844 290448
rect 84896 290436 84902 290488
rect 88610 290436 88616 290488
rect 88668 290476 88674 290488
rect 99558 290476 99564 290488
rect 88668 290448 99564 290476
rect 88668 290436 88674 290448
rect 99558 290436 99564 290448
rect 99616 290436 99622 290488
rect 258718 290436 258724 290488
rect 258776 290476 258782 290488
rect 274818 290476 274824 290488
rect 258776 290448 274824 290476
rect 258776 290436 258782 290448
rect 274818 290436 274824 290448
rect 274876 290436 274882 290488
rect 184842 290300 184848 290352
rect 184900 290340 184906 290352
rect 188890 290340 188896 290352
rect 184900 290312 188896 290340
rect 184900 290300 184906 290312
rect 188890 290300 188896 290312
rect 188948 290340 188954 290352
rect 191742 290340 191748 290352
rect 188948 290312 191748 290340
rect 188948 290300 188954 290312
rect 191742 290300 191748 290312
rect 191800 290300 191806 290352
rect 61838 290096 61844 290148
rect 61896 290136 61902 290148
rect 62758 290136 62764 290148
rect 61896 290108 62764 290136
rect 61896 290096 61902 290108
rect 62758 290096 62764 290108
rect 62816 290096 62822 290148
rect 108390 289824 108396 289876
rect 108448 289864 108454 289876
rect 184842 289864 184848 289876
rect 108448 289836 184848 289864
rect 108448 289824 108454 289836
rect 184842 289824 184848 289836
rect 184900 289824 184906 289876
rect 169754 289756 169760 289808
rect 169812 289796 169818 289808
rect 171042 289796 171048 289808
rect 169812 289768 171048 289796
rect 169812 289756 169818 289768
rect 171042 289756 171048 289768
rect 171100 289796 171106 289808
rect 191558 289796 191564 289808
rect 171100 289768 191564 289796
rect 171100 289756 171106 289768
rect 191558 289756 191564 289768
rect 191616 289756 191622 289808
rect 255498 289756 255504 289808
rect 255556 289796 255562 289808
rect 267826 289796 267832 289808
rect 255556 289768 267832 289796
rect 255556 289756 255562 289768
rect 267826 289756 267832 289768
rect 267884 289796 267890 289808
rect 274818 289796 274824 289808
rect 267884 289768 274824 289796
rect 267884 289756 267890 289768
rect 274818 289756 274824 289768
rect 274876 289756 274882 289808
rect 118970 289144 118976 289196
rect 119028 289184 119034 289196
rect 151170 289184 151176 289196
rect 119028 289156 151176 289184
rect 119028 289144 119034 289156
rect 151170 289144 151176 289156
rect 151228 289144 151234 289196
rect 91002 289076 91008 289128
rect 91060 289116 91066 289128
rect 185578 289116 185584 289128
rect 91060 289088 185584 289116
rect 91060 289076 91066 289088
rect 185578 289076 185584 289088
rect 185636 289076 185642 289128
rect 253658 288736 253664 288788
rect 253716 288776 253722 288788
rect 254118 288776 254124 288788
rect 253716 288748 254124 288776
rect 253716 288736 253722 288748
rect 254118 288736 254124 288748
rect 254176 288736 254182 288788
rect 56318 288464 56324 288516
rect 56376 288504 56382 288516
rect 72510 288504 72516 288516
rect 56376 288476 72516 288504
rect 56376 288464 56382 288476
rect 72510 288464 72516 288476
rect 72568 288464 72574 288516
rect 90266 288464 90272 288516
rect 90324 288504 90330 288516
rect 91002 288504 91008 288516
rect 90324 288476 91008 288504
rect 90324 288464 90330 288476
rect 91002 288464 91008 288476
rect 91060 288464 91066 288516
rect 67358 288396 67364 288448
rect 67416 288436 67422 288448
rect 118050 288436 118056 288448
rect 67416 288408 118056 288436
rect 67416 288396 67422 288408
rect 118050 288396 118056 288408
rect 118108 288396 118114 288448
rect 253842 288396 253848 288448
rect 253900 288436 253906 288448
rect 269206 288436 269212 288448
rect 253900 288408 269212 288436
rect 253900 288396 253906 288408
rect 269206 288396 269212 288408
rect 269264 288396 269270 288448
rect 7558 288328 7564 288380
rect 7616 288368 7622 288380
rect 37090 288368 37096 288380
rect 7616 288340 37096 288368
rect 7616 288328 7622 288340
rect 37090 288328 37096 288340
rect 37148 288328 37154 288380
rect 166534 288328 166540 288380
rect 166592 288368 166598 288380
rect 166902 288368 166908 288380
rect 166592 288340 166908 288368
rect 166592 288328 166598 288340
rect 166902 288328 166908 288340
rect 166960 288368 166966 288380
rect 191742 288368 191748 288380
rect 166960 288340 191748 288368
rect 166960 288328 166966 288340
rect 191742 288328 191748 288340
rect 191800 288328 191806 288380
rect 255314 288328 255320 288380
rect 255372 288368 255378 288380
rect 265250 288368 265256 288380
rect 255372 288340 265256 288368
rect 255372 288328 255378 288340
rect 265250 288328 265256 288340
rect 265308 288328 265314 288380
rect 171870 288260 171876 288312
rect 171928 288300 171934 288312
rect 172422 288300 172428 288312
rect 171928 288272 172428 288300
rect 171928 288260 171934 288272
rect 172422 288260 172428 288272
rect 172480 288300 172486 288312
rect 190638 288300 190644 288312
rect 172480 288272 190644 288300
rect 172480 288260 172486 288272
rect 190638 288260 190644 288272
rect 190696 288260 190702 288312
rect 255498 288260 255504 288312
rect 255556 288300 255562 288312
rect 261018 288300 261024 288312
rect 255556 288272 261024 288300
rect 255556 288260 255562 288272
rect 261018 288260 261024 288272
rect 261076 288260 261082 288312
rect 68646 287716 68652 287768
rect 68704 287756 68710 287768
rect 78674 287756 78680 287768
rect 68704 287728 78680 287756
rect 68704 287716 68710 287728
rect 78674 287716 78680 287728
rect 78732 287716 78738 287768
rect 157978 287716 157984 287768
rect 158036 287756 158042 287768
rect 166534 287756 166540 287768
rect 158036 287728 166540 287756
rect 158036 287716 158042 287728
rect 166534 287716 166540 287728
rect 166592 287716 166598 287768
rect 37090 287648 37096 287700
rect 37148 287688 37154 287700
rect 70486 287688 70492 287700
rect 37148 287660 70492 287688
rect 37148 287648 37154 287660
rect 70486 287648 70492 287660
rect 70544 287648 70550 287700
rect 159358 287648 159364 287700
rect 159416 287688 159422 287700
rect 171870 287688 171876 287700
rect 159416 287660 171876 287688
rect 159416 287648 159422 287660
rect 171870 287648 171876 287660
rect 171928 287648 171934 287700
rect 88058 287104 88064 287156
rect 88116 287144 88122 287156
rect 93762 287144 93768 287156
rect 88116 287116 93768 287144
rect 88116 287104 88122 287116
rect 93762 287104 93768 287116
rect 93820 287144 93826 287156
rect 157978 287144 157984 287156
rect 93820 287116 157984 287144
rect 93820 287104 93826 287116
rect 157978 287104 157984 287116
rect 158036 287104 158042 287156
rect 159358 287076 159364 287088
rect 82786 287048 159364 287076
rect 75822 286968 75828 287020
rect 75880 287008 75886 287020
rect 77938 287008 77944 287020
rect 75880 286980 77944 287008
rect 75880 286968 75886 286980
rect 77938 286968 77944 286980
rect 77996 286968 78002 287020
rect 79226 286968 79232 287020
rect 79284 287008 79290 287020
rect 79962 287008 79968 287020
rect 79284 286980 79968 287008
rect 79284 286968 79290 286980
rect 79962 286968 79968 286980
rect 80020 287008 80026 287020
rect 82786 287008 82814 287048
rect 159358 287036 159364 287048
rect 159416 287036 159422 287088
rect 80020 286980 82814 287008
rect 80020 286968 80026 286980
rect 255498 286968 255504 287020
rect 255556 287008 255562 287020
rect 276106 287008 276112 287020
rect 255556 286980 276112 287008
rect 255556 286968 255562 286980
rect 276106 286968 276112 286980
rect 276164 286968 276170 287020
rect 255406 286900 255412 286952
rect 255464 286940 255470 286952
rect 262214 286940 262220 286952
rect 255464 286912 262220 286940
rect 255464 286900 255470 286912
rect 262214 286900 262220 286912
rect 262272 286900 262278 286952
rect 97442 286560 97448 286612
rect 97500 286600 97506 286612
rect 97902 286600 97908 286612
rect 97500 286572 97908 286600
rect 97500 286560 97506 286572
rect 97902 286560 97908 286572
rect 97960 286560 97966 286612
rect 81986 286424 81992 286476
rect 82044 286464 82050 286476
rect 83458 286464 83464 286476
rect 82044 286436 83464 286464
rect 82044 286424 82050 286436
rect 83458 286424 83464 286436
rect 83516 286424 83522 286476
rect 86862 286288 86868 286340
rect 86920 286328 86926 286340
rect 88978 286328 88984 286340
rect 86920 286300 88984 286328
rect 86920 286288 86926 286300
rect 88978 286288 88984 286300
rect 89036 286288 89042 286340
rect 169754 286288 169760 286340
rect 169812 286328 169818 286340
rect 170582 286328 170588 286340
rect 169812 286300 170588 286328
rect 169812 286288 169818 286300
rect 170582 286288 170588 286300
rect 170640 286328 170646 286340
rect 180150 286328 180156 286340
rect 170640 286300 180156 286328
rect 170640 286288 170646 286300
rect 180150 286288 180156 286300
rect 180208 286288 180214 286340
rect 50982 285744 50988 285796
rect 51040 285784 51046 285796
rect 69106 285784 69112 285796
rect 51040 285756 69112 285784
rect 51040 285744 51046 285756
rect 69106 285744 69112 285756
rect 69164 285784 69170 285796
rect 69658 285784 69664 285796
rect 69164 285756 69664 285784
rect 69164 285744 69170 285756
rect 69658 285744 69664 285756
rect 69716 285744 69722 285796
rect 70302 285744 70308 285796
rect 70360 285784 70366 285796
rect 76006 285784 76012 285796
rect 70360 285756 76012 285784
rect 70360 285744 70366 285756
rect 76006 285744 76012 285756
rect 76064 285744 76070 285796
rect 78582 285744 78588 285796
rect 78640 285784 78646 285796
rect 78640 285756 80054 285784
rect 78640 285744 78646 285756
rect 73614 285716 73620 285728
rect 52380 285688 73620 285716
rect 45462 285540 45468 285592
rect 45520 285580 45526 285592
rect 51718 285580 51724 285592
rect 45520 285552 51724 285580
rect 45520 285540 45526 285552
rect 51718 285540 51724 285552
rect 51776 285580 51782 285592
rect 52380 285580 52408 285688
rect 73614 285676 73620 285688
rect 73672 285676 73678 285728
rect 80026 285716 80054 285756
rect 90818 285744 90824 285796
rect 90876 285784 90882 285796
rect 112438 285784 112444 285796
rect 90876 285756 112444 285784
rect 90876 285744 90882 285756
rect 112438 285744 112444 285756
rect 112496 285744 112502 285796
rect 160922 285744 160928 285796
rect 160980 285784 160986 285796
rect 191006 285784 191012 285796
rect 160980 285756 191012 285784
rect 160980 285744 160986 285756
rect 191006 285744 191012 285756
rect 191064 285744 191070 285796
rect 169754 285716 169760 285728
rect 80026 285688 169760 285716
rect 169754 285676 169760 285688
rect 169812 285676 169818 285728
rect 80146 285648 80152 285660
rect 51776 285552 52408 285580
rect 55186 285620 80152 285648
rect 51776 285540 51782 285552
rect 48130 285472 48136 285524
rect 48188 285512 48194 285524
rect 55186 285512 55214 285620
rect 80146 285608 80152 285620
rect 80204 285608 80210 285660
rect 48188 285484 55214 285512
rect 48188 285472 48194 285484
rect 177298 284928 177304 284980
rect 177356 284968 177362 284980
rect 191742 284968 191748 284980
rect 177356 284940 191748 284968
rect 177356 284928 177362 284940
rect 191742 284928 191748 284940
rect 191800 284928 191806 284980
rect 96430 284384 96436 284436
rect 96488 284424 96494 284436
rect 96488 284396 99374 284424
rect 96488 284384 96494 284396
rect 92382 284316 92388 284368
rect 92440 284356 92446 284368
rect 99006 284356 99012 284368
rect 92440 284328 99012 284356
rect 92440 284316 92446 284328
rect 99006 284316 99012 284328
rect 99064 284316 99070 284368
rect 99346 284356 99374 284396
rect 115842 284356 115848 284368
rect 99346 284328 115848 284356
rect 115842 284316 115848 284328
rect 115900 284316 115906 284368
rect 176562 284316 176568 284368
rect 176620 284356 176626 284368
rect 178034 284356 178040 284368
rect 176620 284328 178040 284356
rect 176620 284316 176626 284328
rect 178034 284316 178040 284328
rect 178092 284316 178098 284368
rect 263686 284316 263692 284368
rect 263744 284356 263750 284368
rect 264882 284356 264888 284368
rect 263744 284328 264888 284356
rect 263744 284316 263750 284328
rect 264882 284316 264888 284328
rect 264940 284316 264946 284368
rect 152642 284248 152648 284300
rect 152700 284288 152706 284300
rect 193030 284288 193036 284300
rect 152700 284260 193036 284288
rect 152700 284248 152706 284260
rect 193030 284248 193036 284260
rect 193088 284248 193094 284300
rect 255498 284248 255504 284300
rect 255556 284288 255562 284300
rect 266446 284288 266452 284300
rect 255556 284260 266452 284288
rect 255556 284248 255562 284260
rect 266446 284248 266452 284260
rect 266504 284288 266510 284300
rect 267826 284288 267832 284300
rect 266504 284260 267832 284288
rect 266504 284248 266510 284260
rect 267826 284248 267832 284260
rect 267884 284248 267890 284300
rect 259086 284180 259092 284232
rect 259144 284220 259150 284232
rect 266538 284220 266544 284232
rect 259144 284192 266544 284220
rect 259144 284180 259150 284192
rect 266538 284180 266544 284192
rect 266596 284180 266602 284232
rect 130562 283568 130568 283620
rect 130620 283608 130626 283620
rect 152642 283608 152648 283620
rect 130620 283580 152648 283608
rect 130620 283568 130626 283580
rect 152642 283568 152648 283580
rect 152700 283568 152706 283620
rect 73246 283432 73252 283484
rect 73304 283432 73310 283484
rect 73264 283404 73292 283432
rect 74718 283404 74724 283416
rect 73264 283376 74724 283404
rect 74718 283364 74724 283376
rect 74776 283364 74782 283416
rect 92474 283364 92480 283416
rect 92532 283404 92538 283416
rect 92934 283404 92940 283416
rect 92532 283376 92940 283404
rect 92532 283364 92538 283376
rect 92934 283364 92940 283376
rect 92992 283364 92998 283416
rect 99098 283268 99104 283280
rect 70366 283240 99104 283268
rect 67542 283024 67548 283076
rect 67600 283064 67606 283076
rect 70366 283064 70394 283240
rect 99098 283228 99104 283240
rect 99156 283228 99162 283280
rect 67600 283036 70394 283064
rect 67600 283024 67606 283036
rect 70946 283024 70952 283076
rect 71004 283064 71010 283076
rect 98822 283064 98828 283076
rect 71004 283036 98828 283064
rect 71004 283024 71010 283036
rect 98822 283024 98828 283036
rect 98880 283024 98886 283076
rect 64690 282956 64696 283008
rect 64748 282996 64754 283008
rect 66806 282996 66812 283008
rect 64748 282968 66812 282996
rect 64748 282956 64754 282968
rect 66806 282956 66812 282968
rect 66864 282956 66870 283008
rect 75362 282956 75368 283008
rect 75420 282956 75426 283008
rect 81250 282956 81256 283008
rect 81308 282956 81314 283008
rect 89530 282956 89536 283008
rect 89588 282956 89594 283008
rect 65886 282208 65892 282260
rect 65944 282248 65950 282260
rect 66162 282248 66168 282260
rect 65944 282220 66168 282248
rect 65944 282208 65950 282220
rect 66162 282208 66168 282220
rect 66220 282208 66226 282260
rect 57790 282140 57796 282192
rect 57848 282180 57854 282192
rect 67082 282180 67088 282192
rect 57848 282152 67088 282180
rect 57848 282140 57854 282152
rect 67082 282140 67088 282152
rect 67140 282140 67146 282192
rect 67266 282140 67272 282192
rect 67324 282180 67330 282192
rect 75380 282180 75408 282956
rect 81268 282860 81296 282956
rect 89548 282860 89576 282956
rect 97994 282860 98000 282872
rect 81268 282832 84194 282860
rect 89548 282832 98000 282860
rect 67324 282152 75408 282180
rect 67324 282140 67330 282152
rect 84166 281636 84194 282832
rect 97994 282820 98000 282832
rect 98052 282820 98058 282872
rect 168466 282820 168472 282872
rect 168524 282860 168530 282872
rect 169570 282860 169576 282872
rect 168524 282832 169576 282860
rect 168524 282820 168530 282832
rect 169570 282820 169576 282832
rect 169628 282860 169634 282872
rect 191558 282860 191564 282872
rect 169628 282832 191564 282860
rect 169628 282820 169634 282832
rect 191558 282820 191564 282832
rect 191616 282820 191622 282872
rect 255498 282820 255504 282872
rect 255556 282860 255562 282872
rect 268010 282860 268016 282872
rect 255556 282832 268016 282860
rect 255556 282820 255562 282832
rect 268010 282820 268016 282832
rect 268068 282820 268074 282872
rect 100754 282684 100760 282736
rect 100812 282724 100818 282736
rect 102870 282724 102876 282736
rect 100812 282696 102876 282724
rect 100812 282684 100818 282696
rect 102870 282684 102876 282696
rect 102928 282684 102934 282736
rect 115842 282140 115848 282192
rect 115900 282180 115906 282192
rect 149698 282180 149704 282192
rect 115900 282152 149704 282180
rect 115900 282140 115906 282152
rect 149698 282140 149704 282152
rect 149756 282180 149762 282192
rect 168466 282180 168472 282192
rect 149756 282152 168472 282180
rect 149756 282140 149762 282152
rect 168466 282140 168472 282152
rect 168524 282140 168530 282192
rect 255406 281868 255412 281920
rect 255464 281908 255470 281920
rect 259454 281908 259460 281920
rect 255464 281880 259460 281908
rect 255464 281868 255470 281880
rect 259454 281868 259460 281880
rect 259512 281868 259518 281920
rect 98914 281636 98920 281648
rect 84166 281608 98920 281636
rect 98914 281596 98920 281608
rect 98972 281596 98978 281648
rect 97994 281528 98000 281580
rect 98052 281568 98058 281580
rect 173802 281568 173808 281580
rect 98052 281540 173808 281568
rect 98052 281528 98058 281540
rect 173802 281528 173808 281540
rect 173860 281528 173866 281580
rect 184290 281528 184296 281580
rect 184348 281568 184354 281580
rect 191742 281568 191748 281580
rect 184348 281540 191748 281568
rect 184348 281528 184354 281540
rect 191742 281528 191748 281540
rect 191800 281528 191806 281580
rect 100754 281460 100760 281512
rect 100812 281500 100818 281512
rect 118970 281500 118976 281512
rect 100812 281472 118976 281500
rect 100812 281460 100818 281472
rect 118970 281460 118976 281472
rect 119028 281460 119034 281512
rect 168282 281460 168288 281512
rect 168340 281500 168346 281512
rect 171870 281500 171876 281512
rect 168340 281472 171876 281500
rect 168340 281460 168346 281472
rect 171870 281460 171876 281472
rect 171928 281460 171934 281512
rect 255406 281324 255412 281376
rect 255464 281364 255470 281376
rect 259086 281364 259092 281376
rect 255464 281336 259092 281364
rect 255464 281324 255470 281336
rect 259086 281324 259092 281336
rect 259144 281324 259150 281376
rect 255406 281188 255412 281240
rect 255464 281228 255470 281240
rect 259730 281228 259736 281240
rect 255464 281200 259736 281228
rect 255464 281188 255470 281200
rect 259730 281188 259736 281200
rect 259788 281188 259794 281240
rect 167730 280780 167736 280832
rect 167788 280820 167794 280832
rect 175918 280820 175924 280832
rect 167788 280792 175924 280820
rect 167788 280780 167794 280792
rect 175918 280780 175924 280792
rect 175976 280780 175982 280832
rect 61746 280236 61752 280288
rect 61804 280276 61810 280288
rect 66898 280276 66904 280288
rect 61804 280248 66904 280276
rect 61804 280236 61810 280248
rect 66898 280236 66904 280248
rect 66956 280236 66962 280288
rect 14458 280168 14464 280220
rect 14516 280208 14522 280220
rect 66530 280208 66536 280220
rect 14516 280180 66536 280208
rect 14516 280168 14522 280180
rect 66530 280168 66536 280180
rect 66588 280208 66594 280220
rect 67174 280208 67180 280220
rect 66588 280180 67180 280208
rect 66588 280168 66594 280180
rect 67174 280168 67180 280180
rect 67232 280168 67238 280220
rect 100846 280168 100852 280220
rect 100904 280208 100910 280220
rect 156690 280208 156696 280220
rect 100904 280180 156696 280208
rect 100904 280168 100910 280180
rect 156690 280168 156696 280180
rect 156748 280168 156754 280220
rect 100754 280100 100760 280152
rect 100812 280140 100818 280152
rect 159542 280140 159548 280152
rect 100812 280112 159548 280140
rect 100812 280100 100818 280112
rect 159542 280100 159548 280112
rect 159600 280100 159606 280152
rect 168466 280100 168472 280152
rect 168524 280140 168530 280152
rect 191558 280140 191564 280152
rect 168524 280112 191564 280140
rect 168524 280100 168530 280112
rect 191558 280100 191564 280112
rect 191616 280100 191622 280152
rect 255406 280100 255412 280152
rect 255464 280140 255470 280152
rect 278958 280140 278964 280152
rect 255464 280112 278964 280140
rect 255464 280100 255470 280112
rect 278958 280100 278964 280112
rect 279016 280100 279022 280152
rect 255498 280032 255504 280084
rect 255556 280072 255562 280084
rect 274726 280072 274732 280084
rect 255556 280044 274732 280072
rect 255556 280032 255562 280044
rect 274726 280032 274732 280044
rect 274784 280032 274790 280084
rect 4062 279420 4068 279472
rect 4120 279460 4126 279472
rect 45370 279460 45376 279472
rect 4120 279432 45376 279460
rect 4120 279420 4126 279432
rect 45370 279420 45376 279432
rect 45428 279460 45434 279472
rect 60550 279460 60556 279472
rect 45428 279432 60556 279460
rect 45428 279420 45434 279432
rect 60550 279420 60556 279432
rect 60608 279460 60614 279472
rect 66622 279460 66628 279472
rect 60608 279432 66628 279460
rect 60608 279420 60614 279432
rect 66622 279420 66628 279432
rect 66680 279420 66686 279472
rect 98822 279420 98828 279472
rect 98880 279460 98886 279472
rect 165522 279460 165528 279472
rect 98880 279432 165528 279460
rect 98880 279420 98886 279432
rect 165522 279420 165528 279432
rect 165580 279460 165586 279472
rect 189902 279460 189908 279472
rect 165580 279432 189908 279460
rect 165580 279420 165586 279432
rect 189902 279420 189908 279432
rect 189960 279420 189966 279472
rect 53558 278672 53564 278724
rect 53616 278712 53622 278724
rect 53742 278712 53748 278724
rect 53616 278684 53748 278712
rect 53616 278672 53622 278684
rect 53742 278672 53748 278684
rect 53800 278672 53806 278724
rect 99098 278672 99104 278724
rect 99156 278712 99162 278724
rect 157334 278712 157340 278724
rect 99156 278684 157340 278712
rect 99156 278672 99162 278684
rect 157334 278672 157340 278684
rect 157392 278672 157398 278724
rect 173802 278672 173808 278724
rect 173860 278712 173866 278724
rect 174630 278712 174636 278724
rect 173860 278684 174636 278712
rect 173860 278672 173866 278684
rect 174630 278672 174636 278684
rect 174688 278672 174694 278724
rect 255406 278672 255412 278724
rect 255464 278712 255470 278724
rect 261110 278712 261116 278724
rect 255464 278684 261116 278712
rect 255464 278672 255470 278684
rect 261110 278672 261116 278684
rect 261168 278672 261174 278724
rect 100754 278604 100760 278656
rect 100812 278644 100818 278656
rect 130470 278644 130476 278656
rect 100812 278616 130476 278644
rect 100812 278604 100818 278616
rect 130470 278604 130476 278616
rect 130528 278604 130534 278656
rect 53558 277992 53564 278044
rect 53616 278032 53622 278044
rect 66806 278032 66812 278044
rect 53616 278004 66812 278032
rect 53616 277992 53622 278004
rect 66806 277992 66812 278004
rect 66864 277992 66870 278044
rect 133230 277992 133236 278044
rect 133288 278032 133294 278044
rect 174538 278032 174544 278044
rect 133288 278004 174544 278032
rect 133288 277992 133294 278004
rect 174538 277992 174544 278004
rect 174596 277992 174602 278044
rect 263686 277516 263692 277568
rect 263744 277556 263750 277568
rect 269298 277556 269304 277568
rect 263744 277528 269304 277556
rect 263744 277516 263750 277528
rect 269298 277516 269304 277528
rect 269356 277516 269362 277568
rect 174630 277380 174636 277432
rect 174688 277420 174694 277432
rect 192846 277420 192852 277432
rect 174688 277392 192852 277420
rect 174688 277380 174694 277392
rect 192846 277380 192852 277392
rect 192904 277380 192910 277432
rect 61654 277312 61660 277364
rect 61712 277352 61718 277364
rect 66898 277352 66904 277364
rect 61712 277324 66904 277352
rect 61712 277312 61718 277324
rect 66898 277312 66904 277324
rect 66956 277312 66962 277364
rect 118050 277312 118056 277364
rect 118108 277352 118114 277364
rect 118108 277324 180794 277352
rect 118108 277312 118114 277324
rect 100754 277244 100760 277296
rect 100812 277284 100818 277296
rect 163498 277284 163504 277296
rect 100812 277256 163504 277284
rect 100812 277244 100818 277256
rect 163498 277244 163504 277256
rect 163556 277244 163562 277296
rect 180766 277284 180794 277324
rect 185486 277312 185492 277364
rect 185544 277352 185550 277364
rect 193214 277352 193220 277364
rect 185544 277324 193220 277352
rect 185544 277312 185550 277324
rect 193214 277312 193220 277324
rect 193272 277312 193278 277364
rect 255406 277312 255412 277364
rect 255464 277352 255470 277364
rect 273530 277352 273536 277364
rect 255464 277324 273536 277352
rect 255464 277312 255470 277324
rect 273530 277312 273536 277324
rect 273588 277312 273594 277364
rect 190454 277284 190460 277296
rect 180766 277256 190460 277284
rect 190454 277244 190460 277256
rect 190512 277284 190518 277296
rect 191282 277284 191288 277296
rect 190512 277256 191288 277284
rect 190512 277244 190518 277256
rect 191282 277244 191288 277256
rect 191340 277244 191346 277296
rect 255498 277244 255504 277296
rect 255556 277284 255562 277296
rect 269390 277284 269396 277296
rect 255556 277256 269396 277284
rect 255556 277244 255562 277256
rect 269390 277244 269396 277256
rect 269448 277244 269454 277296
rect 269390 276020 269396 276072
rect 269448 276060 269454 276072
rect 271874 276060 271880 276072
rect 269448 276032 271880 276060
rect 269448 276020 269454 276032
rect 271874 276020 271880 276032
rect 271932 276020 271938 276072
rect 99006 275952 99012 276004
rect 99064 275992 99070 276004
rect 185578 275992 185584 276004
rect 99064 275964 185584 275992
rect 99064 275952 99070 275964
rect 185578 275952 185584 275964
rect 185636 275952 185642 276004
rect 255406 275952 255412 276004
rect 255464 275992 255470 276004
rect 271966 275992 271972 276004
rect 255464 275964 271972 275992
rect 255464 275952 255470 275964
rect 271966 275952 271972 275964
rect 272024 275952 272030 276004
rect 108298 274660 108304 274712
rect 108356 274700 108362 274712
rect 110414 274700 110420 274712
rect 108356 274672 110420 274700
rect 108356 274660 108362 274672
rect 110414 274660 110420 274672
rect 110472 274660 110478 274712
rect 255406 274660 255412 274712
rect 255464 274700 255470 274712
rect 255464 274672 273944 274700
rect 255464 274660 255470 274672
rect 100754 274592 100760 274644
rect 100812 274632 100818 274644
rect 100812 274604 161474 274632
rect 100812 274592 100818 274604
rect 161446 274564 161474 274604
rect 177850 274592 177856 274644
rect 177908 274632 177914 274644
rect 182174 274632 182180 274644
rect 177908 274604 182180 274632
rect 177908 274592 177914 274604
rect 182174 274592 182180 274604
rect 182232 274592 182238 274644
rect 255498 274592 255504 274644
rect 255556 274632 255562 274644
rect 273438 274632 273444 274644
rect 255556 274604 273444 274632
rect 255556 274592 255562 274604
rect 273438 274592 273444 274604
rect 273496 274592 273502 274644
rect 273916 274576 273944 274672
rect 183002 274564 183008 274576
rect 161446 274536 183008 274564
rect 183002 274524 183008 274536
rect 183060 274524 183066 274576
rect 255406 274524 255412 274576
rect 255464 274564 255470 274576
rect 265158 274564 265164 274576
rect 255464 274536 265164 274564
rect 255464 274524 255470 274536
rect 265158 274524 265164 274536
rect 265216 274564 265222 274576
rect 269298 274564 269304 274576
rect 265216 274536 269304 274564
rect 265216 274524 265222 274536
rect 269298 274524 269304 274536
rect 269356 274524 269362 274576
rect 273898 274524 273904 274576
rect 273956 274564 273962 274576
rect 274634 274564 274640 274576
rect 273956 274536 274640 274564
rect 273956 274524 273962 274536
rect 274634 274524 274640 274536
rect 274692 274524 274698 274576
rect 53742 273912 53748 273964
rect 53800 273952 53806 273964
rect 65886 273952 65892 273964
rect 53800 273924 65892 273952
rect 53800 273912 53806 273924
rect 65886 273912 65892 273924
rect 65944 273952 65950 273964
rect 66530 273952 66536 273964
rect 65944 273924 66536 273952
rect 65944 273912 65950 273924
rect 66530 273912 66536 273924
rect 66588 273912 66594 273964
rect 100754 273164 100760 273216
rect 100812 273204 100818 273216
rect 108942 273204 108948 273216
rect 100812 273176 108948 273204
rect 100812 273164 100818 273176
rect 108942 273164 108948 273176
rect 109000 273164 109006 273216
rect 255498 273164 255504 273216
rect 255556 273204 255562 273216
rect 281718 273204 281724 273216
rect 255556 273176 281724 273204
rect 255556 273164 255562 273176
rect 281718 273164 281724 273176
rect 281776 273164 281782 273216
rect 255406 273096 255412 273148
rect 255464 273136 255470 273148
rect 259454 273136 259460 273148
rect 255464 273108 259460 273136
rect 255464 273096 255470 273108
rect 259454 273096 259460 273108
rect 259512 273096 259518 273148
rect 157334 272552 157340 272604
rect 157392 272592 157398 272604
rect 172514 272592 172520 272604
rect 157392 272564 172520 272592
rect 157392 272552 157398 272564
rect 172514 272552 172520 272564
rect 172572 272592 172578 272604
rect 173802 272592 173808 272604
rect 172572 272564 173808 272592
rect 172572 272552 172578 272564
rect 173802 272552 173808 272564
rect 173860 272552 173866 272604
rect 50890 272484 50896 272536
rect 50948 272524 50954 272536
rect 60458 272524 60464 272536
rect 50948 272496 60464 272524
rect 50948 272484 50954 272496
rect 60458 272484 60464 272496
rect 60516 272484 60522 272536
rect 108942 272484 108948 272536
rect 109000 272524 109006 272536
rect 135990 272524 135996 272536
rect 109000 272496 135996 272524
rect 109000 272484 109006 272496
rect 135990 272484 135996 272496
rect 136048 272484 136054 272536
rect 162210 272484 162216 272536
rect 162268 272524 162274 272536
rect 177298 272524 177304 272536
rect 162268 272496 177304 272524
rect 162268 272484 162274 272496
rect 177298 272484 177304 272496
rect 177356 272484 177362 272536
rect 177390 271940 177396 271992
rect 177448 271980 177454 271992
rect 191742 271980 191748 271992
rect 177448 271952 191748 271980
rect 177448 271940 177454 271952
rect 191742 271940 191748 271952
rect 191800 271940 191806 271992
rect 43990 271872 43996 271924
rect 44048 271912 44054 271924
rect 66622 271912 66628 271924
rect 44048 271884 66628 271912
rect 44048 271872 44054 271884
rect 66622 271872 66628 271884
rect 66680 271872 66686 271924
rect 173802 271872 173808 271924
rect 173860 271912 173866 271924
rect 191650 271912 191656 271924
rect 173860 271884 191656 271912
rect 173860 271872 173866 271884
rect 191650 271872 191656 271884
rect 191708 271872 191714 271924
rect 100754 271804 100760 271856
rect 100812 271844 100818 271856
rect 105630 271844 105636 271856
rect 100812 271816 105636 271844
rect 100812 271804 100818 271816
rect 105630 271804 105636 271816
rect 105688 271804 105694 271856
rect 164142 271804 164148 271856
rect 164200 271844 164206 271856
rect 164878 271844 164884 271856
rect 164200 271816 164884 271844
rect 164200 271804 164206 271816
rect 164878 271804 164884 271816
rect 164936 271844 164942 271856
rect 184290 271844 184296 271856
rect 164936 271816 184296 271844
rect 164936 271804 164942 271816
rect 184290 271804 184296 271816
rect 184348 271804 184354 271856
rect 255406 271804 255412 271856
rect 255464 271844 255470 271856
rect 270678 271844 270684 271856
rect 255464 271816 270684 271844
rect 255464 271804 255470 271816
rect 270678 271804 270684 271816
rect 270736 271804 270742 271856
rect 46842 271124 46848 271176
rect 46900 271164 46906 271176
rect 60550 271164 60556 271176
rect 46900 271136 60556 271164
rect 46900 271124 46906 271136
rect 60550 271124 60556 271136
rect 60608 271124 60614 271176
rect 106182 271124 106188 271176
rect 106240 271164 106246 271176
rect 115198 271164 115204 271176
rect 106240 271136 115204 271164
rect 106240 271124 106246 271136
rect 115198 271124 115204 271136
rect 115256 271124 115262 271176
rect 60550 270512 60556 270564
rect 60608 270552 60614 270564
rect 66254 270552 66260 270564
rect 60608 270524 66260 270552
rect 60608 270512 60614 270524
rect 66254 270512 66260 270524
rect 66312 270512 66318 270564
rect 175918 270512 175924 270564
rect 175976 270552 175982 270564
rect 191742 270552 191748 270564
rect 175976 270524 191748 270552
rect 175976 270512 175982 270524
rect 191742 270512 191748 270524
rect 191800 270512 191806 270564
rect 255406 270512 255412 270564
rect 255464 270552 255470 270564
rect 258258 270552 258264 270564
rect 255464 270524 258264 270552
rect 255464 270512 255470 270524
rect 258258 270512 258264 270524
rect 258316 270552 258322 270564
rect 261018 270552 261024 270564
rect 258316 270524 261024 270552
rect 258316 270512 258322 270524
rect 261018 270512 261024 270524
rect 261076 270512 261082 270564
rect 59170 270444 59176 270496
rect 59228 270484 59234 270496
rect 60642 270484 60648 270496
rect 59228 270456 60648 270484
rect 59228 270444 59234 270456
rect 60642 270444 60648 270456
rect 60700 270444 60706 270496
rect 100754 270444 100760 270496
rect 100812 270484 100818 270496
rect 106090 270484 106096 270496
rect 100812 270456 106096 270484
rect 100812 270444 100818 270456
rect 106090 270444 106096 270456
rect 106148 270444 106154 270496
rect 255498 270444 255504 270496
rect 255556 270484 255562 270496
rect 265066 270484 265072 270496
rect 255556 270456 265072 270484
rect 255556 270444 255562 270456
rect 265066 270444 265072 270456
rect 265124 270444 265130 270496
rect 291286 270444 291292 270496
rect 291344 270484 291350 270496
rect 291654 270484 291660 270496
rect 291344 270456 291660 270484
rect 291344 270444 291350 270456
rect 291654 270444 291660 270456
rect 291712 270484 291718 270496
rect 580166 270484 580172 270496
rect 291712 270456 580172 270484
rect 291712 270444 291718 270456
rect 580166 270444 580172 270456
rect 580224 270444 580230 270496
rect 145650 269832 145656 269884
rect 145708 269872 145714 269884
rect 162118 269872 162124 269884
rect 145708 269844 162124 269872
rect 145708 269832 145714 269844
rect 162118 269832 162124 269844
rect 162176 269832 162182 269884
rect 144822 269764 144828 269816
rect 144880 269804 144886 269816
rect 188430 269804 188436 269816
rect 144880 269776 188436 269804
rect 144880 269764 144886 269776
rect 188430 269764 188436 269776
rect 188488 269764 188494 269816
rect 259362 269764 259368 269816
rect 259420 269804 259426 269816
rect 277486 269804 277492 269816
rect 259420 269776 277492 269804
rect 259420 269764 259426 269776
rect 277486 269764 277492 269776
rect 277544 269764 277550 269816
rect 104250 269084 104256 269136
rect 104308 269124 104314 269136
rect 123478 269124 123484 269136
rect 104308 269096 123484 269124
rect 104308 269084 104314 269096
rect 123478 269084 123484 269096
rect 123536 269084 123542 269136
rect 185762 269084 185768 269136
rect 185820 269124 185826 269136
rect 190822 269124 190828 269136
rect 185820 269096 190828 269124
rect 185820 269084 185826 269096
rect 190822 269084 190828 269096
rect 190880 269084 190886 269136
rect 255406 269084 255412 269136
rect 255464 269124 255470 269136
rect 255464 269096 258074 269124
rect 255464 269084 255470 269096
rect 57882 269016 57888 269068
rect 57940 269056 57946 269068
rect 60642 269056 60648 269068
rect 57940 269028 60648 269056
rect 57940 269016 57946 269028
rect 60642 269016 60648 269028
rect 60700 269016 60706 269068
rect 100754 269016 100760 269068
rect 100812 269056 100818 269068
rect 133230 269056 133236 269068
rect 100812 269028 133236 269056
rect 100812 269016 100818 269028
rect 133230 269016 133236 269028
rect 133288 269016 133294 269068
rect 258046 269056 258074 269096
rect 258718 269056 258724 269068
rect 258046 269028 258724 269056
rect 258718 269016 258724 269028
rect 258776 269056 258782 269068
rect 293954 269056 293960 269068
rect 258776 269028 293960 269056
rect 258776 269016 258782 269028
rect 293954 269016 293960 269028
rect 294012 269016 294018 269068
rect 255406 268948 255412 269000
rect 255464 268988 255470 269000
rect 259362 268988 259368 269000
rect 255464 268960 259368 268988
rect 255464 268948 255470 268960
rect 259362 268948 259368 268960
rect 259420 268948 259426 269000
rect 255498 268880 255504 268932
rect 255556 268920 255562 268932
rect 258810 268920 258816 268932
rect 255556 268892 258816 268920
rect 255556 268880 255562 268892
rect 258810 268880 258816 268892
rect 258868 268880 258874 268932
rect 60642 268404 60648 268456
rect 60700 268444 60706 268456
rect 66898 268444 66904 268456
rect 60700 268416 66904 268444
rect 60700 268404 60706 268416
rect 66898 268404 66904 268416
rect 66956 268404 66962 268456
rect 54846 268336 54852 268388
rect 54904 268376 54910 268388
rect 55030 268376 55036 268388
rect 54904 268348 55036 268376
rect 54904 268336 54910 268348
rect 55030 268336 55036 268348
rect 55088 268376 55094 268388
rect 66806 268376 66812 268388
rect 55088 268348 66812 268376
rect 55088 268336 55094 268348
rect 66806 268336 66812 268348
rect 66864 268336 66870 268388
rect 100754 268336 100760 268388
rect 100812 268376 100818 268388
rect 111058 268376 111064 268388
rect 100812 268348 111064 268376
rect 100812 268336 100818 268348
rect 111058 268336 111064 268348
rect 111116 268336 111122 268388
rect 188430 267792 188436 267844
rect 188488 267832 188494 267844
rect 191742 267832 191748 267844
rect 188488 267804 191748 267832
rect 188488 267792 188494 267804
rect 191742 267792 191748 267804
rect 191800 267792 191806 267844
rect 180150 267724 180156 267776
rect 180208 267764 180214 267776
rect 191466 267764 191472 267776
rect 180208 267736 191472 267764
rect 180208 267724 180214 267736
rect 191466 267724 191472 267736
rect 191524 267724 191530 267776
rect 52362 266976 52368 267028
rect 52420 267016 52426 267028
rect 63218 267016 63224 267028
rect 52420 266988 63224 267016
rect 52420 266976 52426 266988
rect 63218 266976 63224 266988
rect 63276 267016 63282 267028
rect 66622 267016 66628 267028
rect 63276 266988 66628 267016
rect 63276 266976 63282 266988
rect 66622 266976 66628 266988
rect 66680 266976 66686 267028
rect 100754 266976 100760 267028
rect 100812 267016 100818 267028
rect 104802 267016 104808 267028
rect 100812 266988 104808 267016
rect 100812 266976 100818 266988
rect 104802 266976 104808 266988
rect 104860 266976 104866 267028
rect 156414 266976 156420 267028
rect 156472 267016 156478 267028
rect 176010 267016 176016 267028
rect 156472 266988 176016 267016
rect 156472 266976 156478 266988
rect 176010 266976 176016 266988
rect 176068 266976 176074 267028
rect 255406 266976 255412 267028
rect 255464 267016 255470 267028
rect 266814 267016 266820 267028
rect 255464 266988 266820 267016
rect 255464 266976 255470 266988
rect 266814 266976 266820 266988
rect 266872 267016 266878 267028
rect 267642 267016 267648 267028
rect 266872 266988 267648 267016
rect 266872 266976 266878 266988
rect 267642 266976 267648 266988
rect 267700 266976 267706 267028
rect 63310 266364 63316 266416
rect 63368 266404 63374 266416
rect 66438 266404 66444 266416
rect 63368 266376 66444 266404
rect 63368 266364 63374 266376
rect 66438 266364 66444 266376
rect 66496 266364 66502 266416
rect 104802 266364 104808 266416
rect 104860 266404 104866 266416
rect 109770 266404 109776 266416
rect 104860 266376 109776 266404
rect 104860 266364 104866 266376
rect 109770 266364 109776 266376
rect 109828 266364 109834 266416
rect 186958 266364 186964 266416
rect 187016 266404 187022 266416
rect 191742 266404 191748 266416
rect 187016 266376 191748 266404
rect 187016 266364 187022 266376
rect 191742 266364 191748 266376
rect 191800 266364 191806 266416
rect 255498 266364 255504 266416
rect 255556 266404 255562 266416
rect 260926 266404 260932 266416
rect 255556 266376 260932 266404
rect 255556 266364 255562 266376
rect 260926 266364 260932 266376
rect 260984 266364 260990 266416
rect 255406 266296 255412 266348
rect 255464 266336 255470 266348
rect 291378 266336 291384 266348
rect 255464 266308 291384 266336
rect 255464 266296 255470 266308
rect 291378 266296 291384 266308
rect 291436 266296 291442 266348
rect 119430 265684 119436 265736
rect 119488 265724 119494 265736
rect 144270 265724 144276 265736
rect 119488 265696 144276 265724
rect 119488 265684 119494 265696
rect 144270 265684 144276 265696
rect 144328 265684 144334 265736
rect 48038 265616 48044 265668
rect 48096 265656 48102 265668
rect 57238 265656 57244 265668
rect 48096 265628 57244 265656
rect 48096 265616 48102 265628
rect 57238 265616 57244 265628
rect 57296 265616 57302 265668
rect 101490 265616 101496 265668
rect 101548 265656 101554 265668
rect 151262 265656 151268 265668
rect 101548 265628 151268 265656
rect 101548 265616 101554 265628
rect 151262 265616 151268 265628
rect 151320 265616 151326 265668
rect 168282 265616 168288 265668
rect 168340 265656 168346 265668
rect 184934 265656 184940 265668
rect 168340 265628 184940 265656
rect 168340 265616 168346 265628
rect 184934 265616 184940 265628
rect 184992 265616 184998 265668
rect 57238 264936 57244 264988
rect 57296 264976 57302 264988
rect 57882 264976 57888 264988
rect 57296 264948 57888 264976
rect 57296 264936 57302 264948
rect 57882 264936 57888 264948
rect 57940 264976 57946 264988
rect 66806 264976 66812 264988
rect 57940 264948 66812 264976
rect 57940 264936 57946 264948
rect 66806 264936 66812 264948
rect 66864 264936 66870 264988
rect 100754 264936 100760 264988
rect 100812 264976 100818 264988
rect 115198 264976 115204 264988
rect 100812 264948 115204 264976
rect 100812 264936 100818 264948
rect 115198 264936 115204 264948
rect 115256 264936 115262 264988
rect 184198 264936 184204 264988
rect 184256 264976 184262 264988
rect 190822 264976 190828 264988
rect 184256 264948 190828 264976
rect 184256 264936 184262 264948
rect 190822 264936 190828 264948
rect 190880 264936 190886 264988
rect 255498 264936 255504 264988
rect 255556 264976 255562 264988
rect 262490 264976 262496 264988
rect 255556 264948 262496 264976
rect 255556 264936 255562 264948
rect 262490 264936 262496 264948
rect 262548 264936 262554 264988
rect 39942 264188 39948 264240
rect 40000 264228 40006 264240
rect 66254 264228 66260 264240
rect 40000 264200 66260 264228
rect 40000 264188 40006 264200
rect 66254 264188 66260 264200
rect 66312 264188 66318 264240
rect 255406 264188 255412 264240
rect 255464 264228 255470 264240
rect 269850 264228 269856 264240
rect 255464 264200 269856 264228
rect 255464 264188 255470 264200
rect 269850 264188 269856 264200
rect 269908 264188 269914 264240
rect 100846 263644 100852 263696
rect 100904 263684 100910 263696
rect 148502 263684 148508 263696
rect 100904 263656 148508 263684
rect 100904 263644 100910 263656
rect 148502 263644 148508 263656
rect 148560 263644 148566 263696
rect 173158 263644 173164 263696
rect 173216 263684 173222 263696
rect 191742 263684 191748 263696
rect 173216 263656 191748 263684
rect 173216 263644 173222 263656
rect 191742 263644 191748 263656
rect 191800 263644 191806 263696
rect 59078 263576 59084 263628
rect 59136 263616 59142 263628
rect 66806 263616 66812 263628
rect 59136 263588 66812 263616
rect 59136 263576 59142 263588
rect 66806 263576 66812 263588
rect 66864 263576 66870 263628
rect 100754 263576 100760 263628
rect 100812 263616 100818 263628
rect 184290 263616 184296 263628
rect 100812 263588 184296 263616
rect 100812 263576 100818 263588
rect 184290 263576 184296 263588
rect 184348 263576 184354 263628
rect 255406 263576 255412 263628
rect 255464 263616 255470 263628
rect 266538 263616 266544 263628
rect 255464 263588 266544 263616
rect 255464 263576 255470 263588
rect 266538 263576 266544 263588
rect 266596 263616 266602 263628
rect 267182 263616 267188 263628
rect 266596 263588 267188 263616
rect 266596 263576 266602 263588
rect 267182 263576 267188 263588
rect 267240 263576 267246 263628
rect 255038 263236 255044 263288
rect 255096 263276 255102 263288
rect 259270 263276 259276 263288
rect 255096 263248 259276 263276
rect 255096 263236 255102 263248
rect 259270 263236 259276 263248
rect 259328 263236 259334 263288
rect 39298 262828 39304 262880
rect 39356 262868 39362 262880
rect 67082 262868 67088 262880
rect 39356 262840 67088 262868
rect 39356 262828 39362 262840
rect 67082 262828 67088 262840
rect 67140 262828 67146 262880
rect 100754 262828 100760 262880
rect 100812 262868 100818 262880
rect 108390 262868 108396 262880
rect 100812 262840 108396 262868
rect 100812 262828 100818 262840
rect 108390 262828 108396 262840
rect 108448 262828 108454 262880
rect 255590 262828 255596 262880
rect 255648 262868 255654 262880
rect 265158 262868 265164 262880
rect 255648 262840 265164 262868
rect 255648 262828 255654 262840
rect 265158 262828 265164 262840
rect 265216 262868 265222 262880
rect 276014 262868 276020 262880
rect 265216 262840 276020 262868
rect 265216 262828 265222 262840
rect 276014 262828 276020 262840
rect 276072 262828 276078 262880
rect 169018 262284 169024 262336
rect 169076 262324 169082 262336
rect 191006 262324 191012 262336
rect 169076 262296 191012 262324
rect 169076 262284 169082 262296
rect 191006 262284 191012 262296
rect 191064 262284 191070 262336
rect 100754 262216 100760 262268
rect 100812 262256 100818 262268
rect 124858 262256 124864 262268
rect 100812 262228 124864 262256
rect 100812 262216 100818 262228
rect 124858 262216 124864 262228
rect 124916 262216 124922 262268
rect 163498 262216 163504 262268
rect 163556 262256 163562 262268
rect 191742 262256 191748 262268
rect 163556 262228 191748 262256
rect 163556 262216 163562 262228
rect 191742 262216 191748 262228
rect 191800 262216 191806 262268
rect 278130 262216 278136 262268
rect 278188 262256 278194 262268
rect 284386 262256 284392 262268
rect 278188 262228 284392 262256
rect 278188 262216 278194 262228
rect 284386 262216 284392 262228
rect 284444 262216 284450 262268
rect 100846 262148 100852 262200
rect 100904 262188 100910 262200
rect 106182 262188 106188 262200
rect 100904 262160 106188 262188
rect 100904 262148 100910 262160
rect 106182 262148 106188 262160
rect 106240 262188 106246 262200
rect 126238 262188 126244 262200
rect 106240 262160 126244 262188
rect 106240 262148 106246 262160
rect 126238 262148 126244 262160
rect 126296 262148 126302 262200
rect 284662 262148 284668 262200
rect 284720 262188 284726 262200
rect 288710 262188 288716 262200
rect 284720 262160 288716 262188
rect 284720 262148 284726 262160
rect 288710 262148 288716 262160
rect 288768 262148 288774 262200
rect 14550 260856 14556 260908
rect 14608 260896 14614 260908
rect 66898 260896 66904 260908
rect 14608 260868 66904 260896
rect 14608 260856 14614 260868
rect 66898 260856 66904 260868
rect 66956 260856 66962 260908
rect 164878 260856 164884 260908
rect 164936 260896 164942 260908
rect 191558 260896 191564 260908
rect 164936 260868 191564 260896
rect 164936 260856 164942 260868
rect 191558 260856 191564 260868
rect 191616 260856 191622 260908
rect 258810 260856 258816 260908
rect 258868 260896 258874 260908
rect 284662 260896 284668 260908
rect 258868 260868 284668 260896
rect 258868 260856 258874 260868
rect 284662 260856 284668 260868
rect 284720 260856 284726 260908
rect 255406 260788 255412 260840
rect 255464 260828 255470 260840
rect 280338 260828 280344 260840
rect 255464 260800 280344 260828
rect 255464 260788 255470 260800
rect 280338 260788 280344 260800
rect 280396 260788 280402 260840
rect 271782 260720 271788 260772
rect 271840 260760 271846 260772
rect 289906 260760 289912 260772
rect 271840 260732 289912 260760
rect 271840 260720 271846 260732
rect 289906 260720 289912 260732
rect 289964 260720 289970 260772
rect 56502 260108 56508 260160
rect 56560 260148 56566 260160
rect 66254 260148 66260 260160
rect 56560 260120 66260 260148
rect 56560 260108 56566 260120
rect 66254 260108 66260 260120
rect 66312 260108 66318 260160
rect 169110 259632 169116 259684
rect 169168 259672 169174 259684
rect 170674 259672 170680 259684
rect 169168 259644 170680 259672
rect 169168 259632 169174 259644
rect 170674 259632 170680 259644
rect 170732 259632 170738 259684
rect 100754 259496 100760 259548
rect 100812 259536 100818 259548
rect 133230 259536 133236 259548
rect 100812 259508 133236 259536
rect 100812 259496 100818 259508
rect 133230 259496 133236 259508
rect 133288 259496 133294 259548
rect 100846 259428 100852 259480
rect 100904 259468 100910 259480
rect 145742 259468 145748 259480
rect 100904 259440 145748 259468
rect 100904 259428 100910 259440
rect 145742 259428 145748 259440
rect 145800 259428 145806 259480
rect 170398 259428 170404 259480
rect 170456 259468 170462 259480
rect 191742 259468 191748 259480
rect 170456 259440 191748 259468
rect 170456 259428 170462 259440
rect 191742 259428 191748 259440
rect 191800 259428 191806 259480
rect 255498 259428 255504 259480
rect 255556 259468 255562 259480
rect 270678 259468 270684 259480
rect 255556 259440 270684 259468
rect 255556 259428 255562 259440
rect 270678 259428 270684 259440
rect 270736 259468 270742 259480
rect 271782 259468 271788 259480
rect 270736 259440 271788 259468
rect 270736 259428 270742 259440
rect 271782 259428 271788 259440
rect 271840 259428 271846 259480
rect 255406 259360 255412 259412
rect 255464 259400 255470 259412
rect 260742 259400 260748 259412
rect 255464 259372 260748 259400
rect 255464 259360 255470 259372
rect 260742 259360 260748 259372
rect 260800 259360 260806 259412
rect 278038 259360 278044 259412
rect 278096 259400 278102 259412
rect 281626 259400 281632 259412
rect 278096 259372 281632 259400
rect 278096 259360 278102 259372
rect 281626 259360 281632 259372
rect 281684 259400 281690 259412
rect 580166 259400 580172 259412
rect 281684 259372 580172 259400
rect 281684 259360 281690 259372
rect 580166 259360 580172 259372
rect 580224 259360 580230 259412
rect 49602 258680 49608 258732
rect 49660 258720 49666 258732
rect 64782 258720 64788 258732
rect 49660 258692 64788 258720
rect 49660 258680 49666 258692
rect 64782 258680 64788 258692
rect 64840 258720 64846 258732
rect 66438 258720 66444 258732
rect 64840 258692 66444 258720
rect 64840 258680 64846 258692
rect 66438 258680 66444 258692
rect 66496 258680 66502 258732
rect 101674 258680 101680 258732
rect 101732 258720 101738 258732
rect 155402 258720 155408 258732
rect 101732 258692 155408 258720
rect 101732 258680 101738 258692
rect 155402 258680 155408 258692
rect 155460 258680 155466 258732
rect 167638 258136 167644 258188
rect 167696 258176 167702 258188
rect 191742 258176 191748 258188
rect 167696 258148 191748 258176
rect 167696 258136 167702 258148
rect 191742 258136 191748 258148
rect 191800 258136 191806 258188
rect 126238 258068 126244 258120
rect 126296 258108 126302 258120
rect 190638 258108 190644 258120
rect 126296 258080 190644 258108
rect 126296 258068 126302 258080
rect 190638 258068 190644 258080
rect 190696 258068 190702 258120
rect 258166 258068 258172 258120
rect 258224 258108 258230 258120
rect 285950 258108 285956 258120
rect 258224 258080 285956 258108
rect 258224 258068 258230 258080
rect 285950 258068 285956 258080
rect 286008 258108 286014 258120
rect 287054 258108 287060 258120
rect 286008 258080 287060 258108
rect 286008 258068 286014 258080
rect 287054 258068 287060 258080
rect 287112 258068 287118 258120
rect 50706 258000 50712 258052
rect 50764 258040 50770 258052
rect 66254 258040 66260 258052
rect 50764 258012 66260 258040
rect 50764 258000 50770 258012
rect 66254 258000 66260 258012
rect 66312 258000 66318 258052
rect 66438 258000 66444 258052
rect 66496 258040 66502 258052
rect 68186 258040 68192 258052
rect 66496 258012 68192 258040
rect 66496 258000 66502 258012
rect 68186 258000 68192 258012
rect 68244 258000 68250 258052
rect 190730 258000 190736 258052
rect 190788 258040 190794 258052
rect 193398 258040 193404 258052
rect 190788 258012 193404 258040
rect 190788 258000 190794 258012
rect 193398 258000 193404 258012
rect 193456 258000 193462 258052
rect 255406 257388 255412 257440
rect 255464 257428 255470 257440
rect 258810 257428 258816 257440
rect 255464 257400 258816 257428
rect 255464 257388 255470 257400
rect 258810 257388 258816 257400
rect 258868 257388 258874 257440
rect 111150 257320 111156 257372
rect 111208 257360 111214 257372
rect 171962 257360 171968 257372
rect 111208 257332 171968 257360
rect 111208 257320 111214 257332
rect 171962 257320 171968 257332
rect 172020 257320 172026 257372
rect 180610 257320 180616 257372
rect 180668 257360 180674 257372
rect 183554 257360 183560 257372
rect 180668 257332 183560 257360
rect 180668 257320 180674 257332
rect 183554 257320 183560 257332
rect 183612 257320 183618 257372
rect 263778 257320 263784 257372
rect 263836 257360 263842 257372
rect 285858 257360 285864 257372
rect 263836 257332 285864 257360
rect 263836 257320 263842 257332
rect 285858 257320 285864 257332
rect 285916 257320 285922 257372
rect 63402 256844 63408 256896
rect 63460 256884 63466 256896
rect 66622 256884 66628 256896
rect 63460 256856 66628 256884
rect 63460 256844 63466 256856
rect 66622 256844 66628 256856
rect 66680 256844 66686 256896
rect 171778 256708 171784 256760
rect 171836 256748 171842 256760
rect 191650 256748 191656 256760
rect 171836 256720 191656 256748
rect 171836 256708 171842 256720
rect 191650 256708 191656 256720
rect 191708 256708 191714 256760
rect 255406 256708 255412 256760
rect 255464 256748 255470 256760
rect 261110 256748 261116 256760
rect 255464 256720 261116 256748
rect 255464 256708 255470 256720
rect 261110 256708 261116 256720
rect 261168 256708 261174 256760
rect 255498 256028 255504 256080
rect 255556 256068 255562 256080
rect 263778 256068 263784 256080
rect 255556 256040 263784 256068
rect 255556 256028 255562 256040
rect 263778 256028 263784 256040
rect 263836 256028 263842 256080
rect 124122 255960 124128 256012
rect 124180 256000 124186 256012
rect 159450 256000 159456 256012
rect 124180 255972 159456 256000
rect 124180 255960 124186 255972
rect 159450 255960 159456 255972
rect 159508 255960 159514 256012
rect 255406 255960 255412 256012
rect 255464 256000 255470 256012
rect 287698 256000 287704 256012
rect 255464 255972 287704 256000
rect 255464 255960 255470 255972
rect 287698 255960 287704 255972
rect 287756 256000 287762 256012
rect 288618 256000 288624 256012
rect 287756 255972 288624 256000
rect 287756 255960 287762 255972
rect 288618 255960 288624 255972
rect 288676 255960 288682 256012
rect 100846 255348 100852 255400
rect 100904 255388 100910 255400
rect 174814 255388 174820 255400
rect 100904 255360 174820 255388
rect 100904 255348 100910 255360
rect 174814 255348 174820 255360
rect 174872 255348 174878 255400
rect 177298 255348 177304 255400
rect 177356 255388 177362 255400
rect 191006 255388 191012 255400
rect 177356 255360 191012 255388
rect 177356 255348 177362 255360
rect 191006 255348 191012 255360
rect 191064 255348 191070 255400
rect 174538 255280 174544 255332
rect 174596 255320 174602 255332
rect 190822 255320 190828 255332
rect 174596 255292 190828 255320
rect 174596 255280 174602 255292
rect 190822 255280 190828 255292
rect 190880 255280 190886 255332
rect 3142 255212 3148 255264
rect 3200 255252 3206 255264
rect 14458 255252 14464 255264
rect 3200 255224 14464 255252
rect 3200 255212 3206 255224
rect 14458 255212 14464 255224
rect 14516 255212 14522 255264
rect 255498 255212 255504 255264
rect 255556 255252 255562 255264
rect 258166 255252 258172 255264
rect 255556 255224 258172 255252
rect 255556 255212 255562 255224
rect 258166 255212 258172 255224
rect 258224 255212 258230 255264
rect 100846 254940 100852 254992
rect 100904 254980 100910 254992
rect 105538 254980 105544 254992
rect 100904 254952 105544 254980
rect 100904 254940 100910 254952
rect 105538 254940 105544 254952
rect 105596 254940 105602 254992
rect 53466 254532 53472 254584
rect 53524 254572 53530 254584
rect 59262 254572 59268 254584
rect 53524 254544 59268 254572
rect 53524 254532 53530 254544
rect 59262 254532 59268 254544
rect 59320 254572 59326 254584
rect 66806 254572 66812 254584
rect 59320 254544 66812 254572
rect 59320 254532 59326 254544
rect 66806 254532 66812 254544
rect 66864 254532 66870 254584
rect 100846 253920 100852 253972
rect 100904 253960 100910 253972
rect 153930 253960 153936 253972
rect 100904 253932 153936 253960
rect 100904 253920 100910 253932
rect 153930 253920 153936 253932
rect 153988 253920 153994 253972
rect 160738 253920 160744 253972
rect 160796 253960 160802 253972
rect 191650 253960 191656 253972
rect 160796 253932 191656 253960
rect 160796 253920 160802 253932
rect 191650 253920 191656 253932
rect 191708 253920 191714 253972
rect 255406 253920 255412 253972
rect 255464 253960 255470 253972
rect 266630 253960 266636 253972
rect 255464 253932 266636 253960
rect 255464 253920 255470 253932
rect 266630 253920 266636 253932
rect 266688 253960 266694 253972
rect 266906 253960 266912 253972
rect 266688 253932 266912 253960
rect 266688 253920 266694 253932
rect 266906 253920 266912 253932
rect 266964 253920 266970 253972
rect 270402 253852 270408 253904
rect 270460 253892 270466 253904
rect 287146 253892 287152 253904
rect 270460 253864 287152 253892
rect 270460 253852 270466 253864
rect 287146 253852 287152 253864
rect 287204 253852 287210 253904
rect 255406 253240 255412 253292
rect 255464 253280 255470 253292
rect 269390 253280 269396 253292
rect 255464 253252 269396 253280
rect 255464 253240 255470 253252
rect 269390 253240 269396 253252
rect 269448 253280 269454 253292
rect 270402 253280 270408 253292
rect 269448 253252 270408 253280
rect 269448 253240 269454 253252
rect 270402 253240 270408 253252
rect 270460 253240 270466 253292
rect 18598 253172 18604 253224
rect 18656 253212 18662 253224
rect 66990 253212 66996 253224
rect 18656 253184 66996 253212
rect 18656 253172 18662 253184
rect 66990 253172 66996 253184
rect 67048 253212 67054 253224
rect 67266 253212 67272 253224
rect 67048 253184 67272 253212
rect 67048 253172 67054 253184
rect 67266 253172 67272 253184
rect 67324 253172 67330 253224
rect 108390 253172 108396 253224
rect 108448 253212 108454 253224
rect 145650 253212 145656 253224
rect 108448 253184 145656 253212
rect 108448 253172 108454 253184
rect 145650 253172 145656 253184
rect 145708 253172 145714 253224
rect 161014 253172 161020 253224
rect 161072 253212 161078 253224
rect 174722 253212 174728 253224
rect 161072 253184 174728 253212
rect 161072 253172 161078 253184
rect 174722 253172 174728 253184
rect 174780 253172 174786 253224
rect 258534 253172 258540 253224
rect 258592 253212 258598 253224
rect 258592 253184 277394 253212
rect 258592 253172 258598 253184
rect 277366 253144 277394 253184
rect 277578 253172 277584 253224
rect 277636 253212 277642 253224
rect 278130 253212 278136 253224
rect 277636 253184 278136 253212
rect 277636 253172 277642 253184
rect 278130 253172 278136 253184
rect 278188 253172 278194 253224
rect 279418 253144 279424 253156
rect 277366 253116 279424 253144
rect 279418 253104 279424 253116
rect 279476 253144 279482 253156
rect 281626 253144 281632 253156
rect 279476 253116 281632 253144
rect 279476 253104 279482 253116
rect 281626 253104 281632 253116
rect 281684 253104 281690 253156
rect 185670 252628 185676 252680
rect 185728 252668 185734 252680
rect 191650 252668 191656 252680
rect 185728 252640 191656 252668
rect 185728 252628 185734 252640
rect 191650 252628 191656 252640
rect 191708 252628 191714 252680
rect 100846 252560 100852 252612
rect 100904 252600 100910 252612
rect 105538 252600 105544 252612
rect 100904 252572 105544 252600
rect 100904 252560 100910 252572
rect 105538 252560 105544 252572
rect 105596 252560 105602 252612
rect 181438 252560 181444 252612
rect 181496 252600 181502 252612
rect 191558 252600 191564 252612
rect 181496 252572 191564 252600
rect 181496 252560 181502 252572
rect 191558 252560 191564 252572
rect 191616 252560 191622 252612
rect 66898 252492 66904 252544
rect 66956 252532 66962 252544
rect 68278 252532 68284 252544
rect 66956 252504 68284 252532
rect 66956 252492 66962 252504
rect 68278 252492 68284 252504
rect 68336 252492 68342 252544
rect 108482 252492 108488 252544
rect 108540 252532 108546 252544
rect 108850 252532 108856 252544
rect 108540 252504 108856 252532
rect 108540 252492 108546 252504
rect 108850 252492 108856 252504
rect 108908 252532 108914 252544
rect 119338 252532 119344 252544
rect 108908 252504 119344 252532
rect 108908 252492 108914 252504
rect 119338 252492 119344 252504
rect 119396 252492 119402 252544
rect 176470 251880 176476 251932
rect 176528 251920 176534 251932
rect 179414 251920 179420 251932
rect 176528 251892 179420 251920
rect 176528 251880 176534 251892
rect 179414 251880 179420 251892
rect 179472 251880 179478 251932
rect 54938 251812 54944 251864
rect 54996 251852 55002 251864
rect 66806 251852 66812 251864
rect 54996 251824 66812 251852
rect 54996 251812 55002 251824
rect 66806 251812 66812 251824
rect 66864 251812 66870 251864
rect 106918 251812 106924 251864
rect 106976 251852 106982 251864
rect 168374 251852 168380 251864
rect 106976 251824 168380 251852
rect 106976 251812 106982 251824
rect 168374 251812 168380 251824
rect 168432 251852 168438 251864
rect 177482 251852 177488 251864
rect 168432 251824 177488 251852
rect 168432 251812 168438 251824
rect 177482 251812 177488 251824
rect 177540 251812 177546 251864
rect 255406 251812 255412 251864
rect 255464 251852 255470 251864
rect 258258 251852 258264 251864
rect 255464 251824 258264 251852
rect 255464 251812 255470 251824
rect 258258 251812 258264 251824
rect 258316 251812 258322 251864
rect 270402 251812 270408 251864
rect 270460 251852 270466 251864
rect 582374 251852 582380 251864
rect 270460 251824 582380 251852
rect 270460 251812 270466 251824
rect 582374 251812 582380 251824
rect 582432 251812 582438 251864
rect 255498 251200 255504 251252
rect 255556 251240 255562 251252
rect 269390 251240 269396 251252
rect 255556 251212 269396 251240
rect 255556 251200 255562 251212
rect 269390 251200 269396 251212
rect 269448 251240 269454 251252
rect 270402 251240 270408 251252
rect 269448 251212 270408 251240
rect 269448 251200 269454 251212
rect 270402 251200 270408 251212
rect 270460 251200 270466 251252
rect 53650 251132 53656 251184
rect 53708 251172 53714 251184
rect 66806 251172 66812 251184
rect 53708 251144 66812 251172
rect 53708 251132 53714 251144
rect 66806 251132 66812 251144
rect 66864 251132 66870 251184
rect 107838 251132 107844 251184
rect 107896 251172 107902 251184
rect 109678 251172 109684 251184
rect 107896 251144 109684 251172
rect 107896 251132 107902 251144
rect 109678 251132 109684 251144
rect 109736 251132 109742 251184
rect 160002 251132 160008 251184
rect 160060 251172 160066 251184
rect 161106 251172 161112 251184
rect 160060 251144 161112 251172
rect 160060 251132 160066 251144
rect 161106 251132 161112 251144
rect 161164 251132 161170 251184
rect 100846 250996 100852 251048
rect 100904 251036 100910 251048
rect 104250 251036 104256 251048
rect 100904 251008 104256 251036
rect 100904 250996 100910 251008
rect 104250 250996 104256 251008
rect 104308 250996 104314 251048
rect 101950 250452 101956 250504
rect 102008 250492 102014 250504
rect 108482 250492 108488 250504
rect 102008 250464 108488 250492
rect 102008 250452 102014 250464
rect 108482 250452 108488 250464
rect 108540 250452 108546 250504
rect 262306 250452 262312 250504
rect 262364 250492 262370 250504
rect 280246 250492 280252 250504
rect 262364 250464 280252 250492
rect 262364 250452 262370 250464
rect 280246 250452 280252 250464
rect 280304 250452 280310 250504
rect 255866 249908 255872 249960
rect 255924 249948 255930 249960
rect 257338 249948 257344 249960
rect 255924 249920 257344 249948
rect 255924 249908 255930 249920
rect 257338 249908 257344 249920
rect 257396 249908 257402 249960
rect 41230 249772 41236 249824
rect 41288 249812 41294 249824
rect 66438 249812 66444 249824
rect 41288 249784 66444 249812
rect 41288 249772 41294 249784
rect 66438 249772 66444 249784
rect 66496 249772 66502 249824
rect 112530 249772 112536 249824
rect 112588 249812 112594 249824
rect 160002 249812 160008 249824
rect 112588 249784 160008 249812
rect 112588 249772 112594 249784
rect 160002 249772 160008 249784
rect 160060 249772 160066 249824
rect 160830 249772 160836 249824
rect 160888 249812 160894 249824
rect 190638 249812 190644 249824
rect 160888 249784 190644 249812
rect 160888 249772 160894 249784
rect 190638 249772 190644 249784
rect 190696 249772 190702 249824
rect 255498 249772 255504 249824
rect 255556 249812 255562 249824
rect 262306 249812 262312 249824
rect 255556 249784 262312 249812
rect 255556 249772 255562 249784
rect 262306 249772 262312 249784
rect 262364 249772 262370 249824
rect 99190 249704 99196 249756
rect 99248 249744 99254 249756
rect 111794 249744 111800 249756
rect 99248 249716 111800 249744
rect 99248 249704 99254 249716
rect 111794 249704 111800 249716
rect 111852 249704 111858 249756
rect 254946 249704 254952 249756
rect 255004 249744 255010 249756
rect 278038 249744 278044 249756
rect 255004 249716 278044 249744
rect 255004 249704 255010 249716
rect 278038 249704 278044 249716
rect 278096 249704 278102 249756
rect 55122 249024 55128 249076
rect 55180 249064 55186 249076
rect 55858 249064 55864 249076
rect 55180 249036 55864 249064
rect 55180 249024 55186 249036
rect 55858 249024 55864 249036
rect 55916 249064 55922 249076
rect 66622 249064 66628 249076
rect 55916 249036 66628 249064
rect 55916 249024 55922 249036
rect 66622 249024 66628 249036
rect 66680 249024 66686 249076
rect 100846 249024 100852 249076
rect 100904 249064 100910 249076
rect 103606 249064 103612 249076
rect 100904 249036 103612 249064
rect 100904 249024 100910 249036
rect 103606 249024 103612 249036
rect 103664 249024 103670 249076
rect 255406 249024 255412 249076
rect 255464 249064 255470 249076
rect 269022 249064 269028 249076
rect 255464 249036 269028 249064
rect 255464 249024 255470 249036
rect 269022 249024 269028 249036
rect 269080 249024 269086 249076
rect 104802 248548 104808 248600
rect 104860 248588 104866 248600
rect 106274 248588 106280 248600
rect 104860 248560 106280 248588
rect 104860 248548 104866 248560
rect 106274 248548 106280 248560
rect 106332 248548 106338 248600
rect 166258 248480 166264 248532
rect 166316 248520 166322 248532
rect 190822 248520 190828 248532
rect 166316 248492 190828 248520
rect 166316 248480 166322 248492
rect 190822 248480 190828 248492
rect 190880 248480 190886 248532
rect 116670 248412 116676 248464
rect 116728 248452 116734 248464
rect 192478 248452 192484 248464
rect 116728 248424 192484 248452
rect 116728 248412 116734 248424
rect 192478 248412 192484 248424
rect 192536 248412 192542 248464
rect 269022 248412 269028 248464
rect 269080 248452 269086 248464
rect 582374 248452 582380 248464
rect 269080 248424 582380 248452
rect 269080 248412 269086 248424
rect 582374 248412 582380 248424
rect 582432 248412 582438 248464
rect 110966 247664 110972 247716
rect 111024 247704 111030 247716
rect 115934 247704 115940 247716
rect 111024 247676 115940 247704
rect 111024 247664 111030 247676
rect 115934 247664 115940 247676
rect 115992 247664 115998 247716
rect 142982 247664 142988 247716
rect 143040 247704 143046 247716
rect 189902 247704 189908 247716
rect 143040 247676 189908 247704
rect 143040 247664 143046 247676
rect 189902 247664 189908 247676
rect 189960 247664 189966 247716
rect 255498 247664 255504 247716
rect 255556 247704 255562 247716
rect 262674 247704 262680 247716
rect 255556 247676 262680 247704
rect 255556 247664 255562 247676
rect 262674 247664 262680 247676
rect 262732 247664 262738 247716
rect 102778 247052 102784 247104
rect 102836 247092 102842 247104
rect 110414 247092 110420 247104
rect 102836 247064 110420 247092
rect 102836 247052 102842 247064
rect 110414 247052 110420 247064
rect 110472 247092 110478 247104
rect 110966 247092 110972 247104
rect 110472 247064 110972 247092
rect 110472 247052 110478 247064
rect 110966 247052 110972 247064
rect 111024 247052 111030 247104
rect 183002 247052 183008 247104
rect 183060 247092 183066 247104
rect 191650 247092 191656 247104
rect 183060 247064 191656 247092
rect 183060 247052 183066 247064
rect 191650 247052 191656 247064
rect 191708 247052 191714 247104
rect 252922 247052 252928 247104
rect 252980 247092 252986 247104
rect 254026 247092 254032 247104
rect 252980 247064 254032 247092
rect 252980 247052 252986 247064
rect 254026 247052 254032 247064
rect 254084 247052 254090 247104
rect 254210 247052 254216 247104
rect 254268 247092 254274 247104
rect 258166 247092 258172 247104
rect 254268 247064 258172 247092
rect 254268 247052 254274 247064
rect 258166 247052 258172 247064
rect 258224 247052 258230 247104
rect 100846 246304 100852 246356
rect 100904 246344 100910 246356
rect 108298 246344 108304 246356
rect 100904 246316 108304 246344
rect 100904 246304 100910 246316
rect 108298 246304 108304 246316
rect 108356 246304 108362 246356
rect 184842 246304 184848 246356
rect 184900 246344 184906 246356
rect 193674 246344 193680 246356
rect 184900 246316 193680 246344
rect 184900 246304 184906 246316
rect 193674 246304 193680 246316
rect 193732 246304 193738 246356
rect 255406 246304 255412 246356
rect 255464 246344 255470 246356
rect 280154 246344 280160 246356
rect 255464 246316 280160 246344
rect 255464 246304 255470 246316
rect 280154 246304 280160 246316
rect 280212 246304 280218 246356
rect 255406 245760 255412 245812
rect 255464 245800 255470 245812
rect 259638 245800 259644 245812
rect 255464 245772 259644 245800
rect 255464 245760 255470 245772
rect 259638 245760 259644 245772
rect 259696 245760 259702 245812
rect 100846 245624 100852 245676
rect 100904 245664 100910 245676
rect 147122 245664 147128 245676
rect 100904 245636 147128 245664
rect 100904 245624 100910 245636
rect 147122 245624 147128 245636
rect 147180 245624 147186 245676
rect 58986 245556 58992 245608
rect 59044 245596 59050 245608
rect 66806 245596 66812 245608
rect 59044 245568 66812 245596
rect 59044 245556 59050 245568
rect 66806 245556 66812 245568
rect 66864 245556 66870 245608
rect 255406 245556 255412 245608
rect 255464 245596 255470 245608
rect 273346 245596 273352 245608
rect 255464 245568 273352 245596
rect 255464 245556 255470 245568
rect 273346 245556 273352 245568
rect 273404 245556 273410 245608
rect 100846 244944 100852 244996
rect 100904 244984 100910 244996
rect 107746 244984 107752 244996
rect 100904 244956 107752 244984
rect 100904 244944 100910 244956
rect 107746 244944 107752 244956
rect 107804 244944 107810 244996
rect 151354 244944 151360 244996
rect 151412 244984 151418 244996
rect 166350 244984 166356 244996
rect 151412 244956 166356 244984
rect 151412 244944 151418 244956
rect 166350 244944 166356 244956
rect 166408 244984 166414 244996
rect 184474 244984 184480 244996
rect 166408 244956 184480 244984
rect 166408 244944 166414 244956
rect 184474 244944 184480 244956
rect 184532 244944 184538 244996
rect 103606 244876 103612 244928
rect 103664 244916 103670 244928
rect 129734 244916 129740 244928
rect 103664 244888 129740 244916
rect 103664 244876 103670 244888
rect 129734 244876 129740 244888
rect 129792 244876 129798 244928
rect 147030 244876 147036 244928
rect 147088 244916 147094 244928
rect 192938 244916 192944 244928
rect 147088 244888 192944 244916
rect 147088 244876 147094 244888
rect 192938 244876 192944 244888
rect 192996 244876 193002 244928
rect 273346 244876 273352 244928
rect 273404 244916 273410 244928
rect 291286 244916 291292 244928
rect 273404 244888 291292 244916
rect 273404 244876 273410 244888
rect 291286 244876 291292 244888
rect 291344 244876 291350 244928
rect 187142 244264 187148 244316
rect 187200 244304 187206 244316
rect 191650 244304 191656 244316
rect 187200 244276 191656 244304
rect 187200 244264 187206 244276
rect 191650 244264 191656 244276
rect 191708 244264 191714 244316
rect 255498 244264 255504 244316
rect 255556 244304 255562 244316
rect 273346 244304 273352 244316
rect 255556 244276 273352 244304
rect 255556 244264 255562 244276
rect 273346 244264 273352 244276
rect 273404 244264 273410 244316
rect 56410 244196 56416 244248
rect 56468 244236 56474 244248
rect 66806 244236 66812 244248
rect 56468 244208 66812 244236
rect 56468 244196 56474 244208
rect 66806 244196 66812 244208
rect 66864 244196 66870 244248
rect 255406 244196 255412 244248
rect 255464 244236 255470 244248
rect 281810 244236 281816 244248
rect 255464 244208 281816 244236
rect 255464 244196 255470 244208
rect 281810 244196 281816 244208
rect 281868 244236 281874 244248
rect 288618 244236 288624 244248
rect 281868 244208 288624 244236
rect 281868 244196 281874 244208
rect 288618 244196 288624 244208
rect 288676 244196 288682 244248
rect 97994 243516 98000 243568
rect 98052 243556 98058 243568
rect 98270 243556 98276 243568
rect 98052 243528 98276 243556
rect 98052 243516 98058 243528
rect 98270 243516 98276 243528
rect 98328 243516 98334 243568
rect 140130 243556 140136 243568
rect 103486 243528 140136 243556
rect 103486 243012 103514 243528
rect 140130 243516 140136 243528
rect 140188 243516 140194 243568
rect 145742 243516 145748 243568
rect 145800 243556 145806 243568
rect 184382 243556 184388 243568
rect 145800 243528 184388 243556
rect 145800 243516 145806 243528
rect 184382 243516 184388 243528
rect 184440 243516 184446 243568
rect 253198 243516 253204 243568
rect 253256 243556 253262 243568
rect 262398 243556 262404 243568
rect 253256 243528 262404 243556
rect 253256 243516 253262 243528
rect 262398 243516 262404 243528
rect 262456 243516 262462 243568
rect 95988 242984 103514 243012
rect 59262 242904 59268 242956
rect 59320 242944 59326 242956
rect 66622 242944 66628 242956
rect 59320 242916 66628 242944
rect 59320 242904 59326 242916
rect 66622 242904 66628 242916
rect 66680 242904 66686 242956
rect 67634 242904 67640 242956
rect 67692 242944 67698 242956
rect 68646 242944 68652 242956
rect 67692 242916 68652 242944
rect 67692 242904 67698 242916
rect 68646 242904 68652 242916
rect 68704 242904 68710 242956
rect 61746 242156 61752 242208
rect 61804 242196 61810 242208
rect 61804 242168 64874 242196
rect 61804 242156 61810 242168
rect 64846 241788 64874 242168
rect 95988 241800 96016 242984
rect 100846 242904 100852 242956
rect 100904 242944 100910 242956
rect 107010 242944 107016 242956
rect 100904 242916 107016 242944
rect 100904 242904 100910 242916
rect 107010 242904 107016 242916
rect 107068 242904 107074 242956
rect 178678 242904 178684 242956
rect 178736 242944 178742 242956
rect 191650 242944 191656 242956
rect 178736 242916 191656 242944
rect 178736 242904 178742 242916
rect 191650 242904 191656 242916
rect 191708 242904 191714 242956
rect 75362 241788 75368 241800
rect 64846 241760 75368 241788
rect 75362 241748 75368 241760
rect 75420 241748 75426 241800
rect 95970 241748 95976 241800
rect 96028 241748 96034 241800
rect 82630 241612 82636 241664
rect 82688 241652 82694 241664
rect 130562 241652 130568 241664
rect 82688 241624 130568 241652
rect 82688 241612 82694 241624
rect 130562 241612 130568 241624
rect 130620 241612 130626 241664
rect 93210 241544 93216 241596
rect 93268 241584 93274 241596
rect 97718 241584 97724 241596
rect 93268 241556 97724 241584
rect 93268 241544 93274 241556
rect 97718 241544 97724 241556
rect 97776 241544 97782 241596
rect 102226 241544 102232 241596
rect 102284 241584 102290 241596
rect 257062 241584 257068 241596
rect 102284 241556 219434 241584
rect 102284 241544 102290 241556
rect 81434 241476 81440 241528
rect 81492 241516 81498 241528
rect 82400 241516 82406 241528
rect 81492 241488 82406 241516
rect 81492 241476 81498 241488
rect 82400 241476 82406 241488
rect 82458 241476 82464 241528
rect 135990 241476 135996 241528
rect 136048 241516 136054 241528
rect 214006 241516 214012 241528
rect 136048 241488 214012 241516
rect 136048 241476 136054 241488
rect 214006 241476 214012 241488
rect 214064 241516 214070 241528
rect 215202 241516 215208 241528
rect 214064 241488 215208 241516
rect 214064 241476 214070 241488
rect 215202 241476 215208 241488
rect 215260 241476 215266 241528
rect 219406 241516 219434 241556
rect 249076 241556 257068 241584
rect 249076 241528 249104 241556
rect 257062 241544 257068 241556
rect 257120 241544 257126 241596
rect 220078 241516 220084 241528
rect 219406 241488 220084 241516
rect 220078 241476 220084 241488
rect 220136 241476 220142 241528
rect 249058 241476 249064 241528
rect 249116 241476 249122 241528
rect 251910 241476 251916 241528
rect 251968 241516 251974 241528
rect 252922 241516 252928 241528
rect 251968 241488 252928 241516
rect 251968 241476 251974 241488
rect 252922 241476 252928 241488
rect 252980 241476 252986 241528
rect 3510 241408 3516 241460
rect 3568 241448 3574 241460
rect 14550 241448 14556 241460
rect 3568 241420 14556 241448
rect 3568 241408 3574 241420
rect 14550 241408 14556 241420
rect 14608 241408 14614 241460
rect 58526 241408 58532 241460
rect 58584 241448 58590 241460
rect 58894 241448 58900 241460
rect 58584 241420 58900 241448
rect 58584 241408 58590 241420
rect 58894 241408 58900 241420
rect 58952 241448 58958 241460
rect 74672 241448 74678 241460
rect 58952 241420 74678 241448
rect 58952 241408 58958 241420
rect 74672 241408 74678 241420
rect 74730 241408 74736 241460
rect 151262 241408 151268 241460
rect 151320 241448 151326 241460
rect 273438 241448 273444 241460
rect 151320 241420 273444 241448
rect 151320 241408 151326 241420
rect 273438 241408 273444 241420
rect 273496 241448 273502 241460
rect 273898 241448 273904 241460
rect 273496 241420 273904 241448
rect 273496 241408 273502 241420
rect 273898 241408 273904 241420
rect 273956 241408 273962 241460
rect 68922 241340 68928 241392
rect 68980 241380 68986 241392
rect 77478 241380 77484 241392
rect 68980 241352 77484 241380
rect 68980 241340 68986 241352
rect 77478 241340 77484 241352
rect 77536 241340 77542 241392
rect 192938 241340 192944 241392
rect 192996 241380 193002 241392
rect 205174 241380 205180 241392
rect 192996 241352 205180 241380
rect 192996 241340 193002 241352
rect 205174 241340 205180 241352
rect 205232 241340 205238 241392
rect 244274 240796 244280 240848
rect 244332 240836 244338 240848
rect 255406 240836 255412 240848
rect 244332 240808 255412 240836
rect 244332 240796 244338 240808
rect 255406 240796 255412 240808
rect 255464 240796 255470 240848
rect 50890 240728 50896 240780
rect 50948 240768 50954 240780
rect 58526 240768 58532 240780
rect 50948 240740 58532 240768
rect 50948 240728 50954 240740
rect 58526 240728 58532 240740
rect 58584 240728 58590 240780
rect 180242 240728 180248 240780
rect 180300 240768 180306 240780
rect 186314 240768 186320 240780
rect 180300 240740 186320 240768
rect 180300 240728 180306 240740
rect 186314 240728 186320 240740
rect 186372 240728 186378 240780
rect 255590 240728 255596 240780
rect 255648 240768 255654 240780
rect 582558 240768 582564 240780
rect 255648 240740 582564 240768
rect 255648 240728 255654 240740
rect 582558 240728 582564 240740
rect 582616 240728 582622 240780
rect 75914 240116 75920 240168
rect 75972 240156 75978 240168
rect 76558 240156 76564 240168
rect 75972 240128 76564 240156
rect 75972 240116 75978 240128
rect 76558 240116 76564 240128
rect 76616 240116 76622 240168
rect 80054 240116 80060 240168
rect 80112 240156 80118 240168
rect 80974 240156 80980 240168
rect 80112 240128 80980 240156
rect 80112 240116 80118 240128
rect 80974 240116 80980 240128
rect 81032 240116 81038 240168
rect 91094 240116 91100 240168
rect 91152 240156 91158 240168
rect 92290 240156 92296 240168
rect 91152 240128 92296 240156
rect 91152 240116 91158 240128
rect 92290 240116 92296 240128
rect 92348 240116 92354 240168
rect 95234 240116 95240 240168
rect 95292 240156 95298 240168
rect 95878 240156 95884 240168
rect 95292 240128 95884 240156
rect 95292 240116 95298 240128
rect 95878 240116 95884 240128
rect 95936 240116 95942 240168
rect 101398 240116 101404 240168
rect 101456 240156 101462 240168
rect 172606 240156 172612 240168
rect 101456 240128 172612 240156
rect 101456 240116 101462 240128
rect 172606 240116 172612 240128
rect 172664 240116 172670 240168
rect 209038 240116 209044 240168
rect 209096 240156 209102 240168
rect 209096 240128 226380 240156
rect 209096 240116 209102 240128
rect 69474 240048 69480 240100
rect 69532 240088 69538 240100
rect 163590 240088 163596 240100
rect 69532 240060 163596 240088
rect 69532 240048 69538 240060
rect 163590 240048 163596 240060
rect 163648 240088 163654 240100
rect 164050 240088 164056 240100
rect 163648 240060 164056 240088
rect 163648 240048 163654 240060
rect 164050 240048 164056 240060
rect 164108 240048 164114 240100
rect 195238 240088 195244 240100
rect 171106 240060 195244 240088
rect 73890 239980 73896 240032
rect 73948 240020 73954 240032
rect 164970 240020 164976 240032
rect 73948 239992 164976 240020
rect 73948 239980 73954 239992
rect 164970 239980 164976 239992
rect 165028 240020 165034 240032
rect 171106 240020 171134 240060
rect 195238 240048 195244 240060
rect 195296 240048 195302 240100
rect 226352 240088 226380 240128
rect 226352 240060 238754 240088
rect 165028 239992 171134 240020
rect 238726 240020 238754 240060
rect 251818 240048 251824 240100
rect 251876 240088 251882 240100
rect 254026 240088 254032 240100
rect 251876 240060 254032 240088
rect 251876 240048 251882 240060
rect 254026 240048 254032 240060
rect 254084 240048 254090 240100
rect 256878 240020 256884 240032
rect 238726 239992 256884 240020
rect 165028 239980 165034 239992
rect 256878 239980 256884 239992
rect 256936 239980 256942 240032
rect 77478 239912 77484 239964
rect 77536 239952 77542 239964
rect 77938 239952 77944 239964
rect 77536 239924 77944 239952
rect 77536 239912 77542 239924
rect 77938 239912 77944 239924
rect 77996 239912 78002 239964
rect 197354 239436 197360 239488
rect 197412 239476 197418 239488
rect 231854 239476 231860 239488
rect 197412 239448 231860 239476
rect 197412 239436 197418 239448
rect 231854 239436 231860 239448
rect 231912 239436 231918 239488
rect 164050 239368 164056 239420
rect 164108 239408 164114 239420
rect 171134 239408 171140 239420
rect 164108 239380 171140 239408
rect 164108 239368 164114 239380
rect 171134 239368 171140 239380
rect 171192 239408 171198 239420
rect 211890 239408 211896 239420
rect 171192 239380 211896 239408
rect 171192 239368 171198 239380
rect 211890 239368 211896 239380
rect 211948 239368 211954 239420
rect 284294 239408 284300 239420
rect 258046 239380 284300 239408
rect 256050 239232 256056 239284
rect 256108 239272 256114 239284
rect 256786 239272 256792 239284
rect 256108 239244 256792 239272
rect 256108 239232 256114 239244
rect 256786 239232 256792 239244
rect 256844 239272 256850 239284
rect 258046 239272 258074 239380
rect 284294 239368 284300 239380
rect 284352 239368 284358 239420
rect 256844 239244 258074 239272
rect 256844 239232 256850 239244
rect 52362 238756 52368 238808
rect 52420 238796 52426 238808
rect 69198 238796 69204 238808
rect 52420 238768 69204 238796
rect 52420 238756 52426 238768
rect 69198 238756 69204 238768
rect 69256 238756 69262 238808
rect 243538 238756 243544 238808
rect 243596 238796 243602 238808
rect 248506 238796 248512 238808
rect 243596 238768 248512 238796
rect 243596 238756 243602 238768
rect 248506 238756 248512 238768
rect 248564 238756 248570 238808
rect 64598 238688 64604 238740
rect 64656 238728 64662 238740
rect 77662 238728 77668 238740
rect 64656 238700 77668 238728
rect 64656 238688 64662 238700
rect 77662 238688 77668 238700
rect 77720 238688 77726 238740
rect 84286 238688 84292 238740
rect 84344 238728 84350 238740
rect 111886 238728 111892 238740
rect 84344 238700 111892 238728
rect 84344 238688 84350 238700
rect 111886 238688 111892 238700
rect 111944 238728 111950 238740
rect 112530 238728 112536 238740
rect 111944 238700 112536 238728
rect 111944 238688 111950 238700
rect 112530 238688 112536 238700
rect 112588 238688 112594 238740
rect 82814 238620 82820 238672
rect 82872 238660 82878 238672
rect 95142 238660 95148 238672
rect 82872 238632 95148 238660
rect 82872 238620 82878 238632
rect 95142 238620 95148 238632
rect 95200 238620 95206 238672
rect 125502 238076 125508 238128
rect 125560 238116 125566 238128
rect 177390 238116 177396 238128
rect 125560 238088 177396 238116
rect 125560 238076 125566 238088
rect 177390 238076 177396 238088
rect 177448 238076 177454 238128
rect 246298 238076 246304 238128
rect 246356 238116 246362 238128
rect 261110 238116 261116 238128
rect 246356 238088 261116 238116
rect 246356 238076 246362 238088
rect 261110 238076 261116 238088
rect 261168 238076 261174 238128
rect 174814 238008 174820 238060
rect 174872 238048 174878 238060
rect 238846 238048 238852 238060
rect 174872 238020 238852 238048
rect 174872 238008 174878 238020
rect 238846 238008 238852 238020
rect 238904 238048 238910 238060
rect 248414 238048 248420 238060
rect 238904 238020 248420 238048
rect 238904 238008 238910 238020
rect 248414 238008 248420 238020
rect 248472 238008 248478 238060
rect 250346 238008 250352 238060
rect 250404 238048 250410 238060
rect 270678 238048 270684 238060
rect 250404 238020 270684 238048
rect 250404 238008 250410 238020
rect 270678 238008 270684 238020
rect 270736 238008 270742 238060
rect 77662 237396 77668 237448
rect 77720 237436 77726 237448
rect 78030 237436 78036 237448
rect 77720 237408 78036 237436
rect 77720 237396 77726 237408
rect 78030 237396 78036 237408
rect 78088 237396 78094 237448
rect 79962 237396 79968 237448
rect 80020 237436 80026 237448
rect 80146 237436 80152 237448
rect 80020 237408 80152 237436
rect 80020 237396 80026 237408
rect 80146 237396 80152 237408
rect 80204 237396 80210 237448
rect 94682 237396 94688 237448
rect 94740 237436 94746 237448
rect 95326 237436 95332 237448
rect 94740 237408 95332 237436
rect 94740 237396 94746 237408
rect 95326 237396 95332 237408
rect 95384 237396 95390 237448
rect 193214 237396 193220 237448
rect 193272 237436 193278 237448
rect 195974 237436 195980 237448
rect 193272 237408 195980 237436
rect 193272 237396 193278 237408
rect 195974 237396 195980 237408
rect 196032 237396 196038 237448
rect 84194 237328 84200 237380
rect 84252 237368 84258 237380
rect 180242 237368 180248 237380
rect 84252 237340 180248 237368
rect 84252 237328 84258 237340
rect 180242 237328 180248 237340
rect 180300 237328 180306 237380
rect 168282 237260 168288 237312
rect 168340 237300 168346 237312
rect 262490 237300 262496 237312
rect 168340 237272 262496 237300
rect 168340 237260 168346 237272
rect 262490 237260 262496 237272
rect 262548 237260 262554 237312
rect 61838 236716 61844 236768
rect 61896 236756 61902 236768
rect 73430 236756 73436 236768
rect 61896 236728 73436 236756
rect 61896 236716 61902 236728
rect 73430 236716 73436 236728
rect 73488 236716 73494 236768
rect 56318 236648 56324 236700
rect 56376 236688 56382 236700
rect 74626 236688 74632 236700
rect 56376 236660 74632 236688
rect 56376 236648 56382 236660
rect 74626 236648 74632 236660
rect 74684 236648 74690 236700
rect 74810 236648 74816 236700
rect 74868 236688 74874 236700
rect 84930 236688 84936 236700
rect 74868 236660 84936 236688
rect 74868 236648 74874 236660
rect 84930 236648 84936 236660
rect 84988 236648 84994 236700
rect 111058 236648 111064 236700
rect 111116 236688 111122 236700
rect 126422 236688 126428 236700
rect 111116 236660 126428 236688
rect 111116 236648 111122 236660
rect 126422 236648 126428 236660
rect 126480 236648 126486 236700
rect 206278 236648 206284 236700
rect 206336 236688 206342 236700
rect 209774 236688 209780 236700
rect 206336 236660 209780 236688
rect 206336 236648 206342 236660
rect 209774 236648 209780 236660
rect 209832 236648 209838 236700
rect 215938 236648 215944 236700
rect 215996 236688 216002 236700
rect 265158 236688 265164 236700
rect 215996 236660 265164 236688
rect 215996 236648 216002 236660
rect 265158 236648 265164 236660
rect 265216 236648 265222 236700
rect 95142 235968 95148 236020
rect 95200 236008 95206 236020
rect 98178 236008 98184 236020
rect 95200 235980 98184 236008
rect 95200 235968 95206 235980
rect 98178 235968 98184 235980
rect 98236 235968 98242 236020
rect 104618 235968 104624 236020
rect 104676 236008 104682 236020
rect 104986 236008 104992 236020
rect 104676 235980 104992 236008
rect 104676 235968 104682 235980
rect 104986 235968 104992 235980
rect 105044 235968 105050 236020
rect 200758 235968 200764 236020
rect 200816 236008 200822 236020
rect 201862 236008 201868 236020
rect 200816 235980 201868 236008
rect 200816 235968 200822 235980
rect 201862 235968 201868 235980
rect 201920 235968 201926 236020
rect 193674 235764 193680 235816
rect 193732 235804 193738 235816
rect 194778 235804 194784 235816
rect 193732 235776 194784 235804
rect 193732 235764 193738 235776
rect 194778 235764 194784 235776
rect 194836 235804 194842 235816
rect 197354 235804 197360 235816
rect 194836 235776 197360 235804
rect 194836 235764 194842 235776
rect 197354 235764 197360 235776
rect 197412 235764 197418 235816
rect 245562 235288 245568 235340
rect 245620 235328 245626 235340
rect 253198 235328 253204 235340
rect 245620 235300 253204 235328
rect 245620 235288 245626 235300
rect 253198 235288 253204 235300
rect 253256 235288 253262 235340
rect 3510 235220 3516 235272
rect 3568 235260 3574 235272
rect 39298 235260 39304 235272
rect 3568 235232 39304 235260
rect 3568 235220 3574 235232
rect 39298 235220 39304 235232
rect 39356 235220 39362 235272
rect 91186 235220 91192 235272
rect 91244 235260 91250 235272
rect 116578 235260 116584 235272
rect 91244 235232 116584 235260
rect 91244 235220 91250 235232
rect 116578 235220 116584 235232
rect 116636 235260 116642 235272
rect 124214 235260 124220 235272
rect 116636 235232 124220 235260
rect 116636 235220 116642 235232
rect 124214 235220 124220 235232
rect 124272 235220 124278 235272
rect 160002 235220 160008 235272
rect 160060 235260 160066 235272
rect 195146 235260 195152 235272
rect 160060 235232 195152 235260
rect 160060 235220 160066 235232
rect 195146 235220 195152 235232
rect 195204 235220 195210 235272
rect 205174 235220 205180 235272
rect 205232 235260 205238 235272
rect 219434 235260 219440 235272
rect 205232 235232 219440 235260
rect 205232 235220 205238 235232
rect 219434 235220 219440 235232
rect 219492 235220 219498 235272
rect 252462 235220 252468 235272
rect 252520 235260 252526 235272
rect 272058 235260 272064 235272
rect 252520 235232 272064 235260
rect 252520 235220 252526 235232
rect 272058 235220 272064 235232
rect 272116 235220 272122 235272
rect 96522 234608 96528 234660
rect 96580 234648 96586 234660
rect 100846 234648 100852 234660
rect 96580 234620 100852 234648
rect 96580 234608 96586 234620
rect 100846 234608 100852 234620
rect 100904 234608 100910 234660
rect 67450 234540 67456 234592
rect 67508 234580 67514 234592
rect 111150 234580 111156 234592
rect 67508 234552 111156 234580
rect 67508 234540 67514 234552
rect 111150 234540 111156 234552
rect 111208 234540 111214 234592
rect 159542 234540 159548 234592
rect 159600 234580 159606 234592
rect 268010 234580 268016 234592
rect 159600 234552 268016 234580
rect 159600 234540 159606 234552
rect 268010 234540 268016 234552
rect 268068 234540 268074 234592
rect 195146 234472 195152 234524
rect 195204 234512 195210 234524
rect 209038 234512 209044 234524
rect 195204 234484 209044 234512
rect 195204 234472 195210 234484
rect 209038 234472 209044 234484
rect 209096 234472 209102 234524
rect 228358 233860 228364 233912
rect 228416 233900 228422 233912
rect 255314 233900 255320 233912
rect 228416 233872 255320 233900
rect 228416 233860 228422 233872
rect 255314 233860 255320 233872
rect 255372 233860 255378 233912
rect 94774 233656 94780 233708
rect 94832 233696 94838 233708
rect 101398 233696 101404 233708
rect 94832 233668 101404 233696
rect 94832 233656 94838 233668
rect 101398 233656 101404 233668
rect 101456 233656 101462 233708
rect 71774 233180 71780 233232
rect 71832 233220 71838 233232
rect 73062 233220 73068 233232
rect 71832 233192 73068 233220
rect 71832 233180 71838 233192
rect 73062 233180 73068 233192
rect 73120 233220 73126 233232
rect 151354 233220 151360 233232
rect 73120 233192 151360 233220
rect 73120 233180 73126 233192
rect 151354 233180 151360 233192
rect 151412 233180 151418 233232
rect 176470 233180 176476 233232
rect 176528 233220 176534 233232
rect 269390 233220 269396 233232
rect 176528 233192 269396 233220
rect 176528 233180 176534 233192
rect 269390 233180 269396 233192
rect 269448 233180 269454 233232
rect 76006 233112 76012 233164
rect 76064 233152 76070 233164
rect 76558 233152 76564 233164
rect 76064 233124 76564 233152
rect 76064 233112 76070 233124
rect 76558 233112 76564 233124
rect 76616 233152 76622 233164
rect 116670 233152 116676 233164
rect 76616 233124 116676 233152
rect 76616 233112 76622 233124
rect 116670 233112 116676 233124
rect 116728 233112 116734 233164
rect 156690 233112 156696 233164
rect 156748 233152 156754 233164
rect 230474 233152 230480 233164
rect 156748 233124 230480 233152
rect 156748 233112 156754 233124
rect 230474 233112 230480 233124
rect 230532 233152 230538 233164
rect 231762 233152 231768 233164
rect 230532 233124 231768 233152
rect 230532 233112 230538 233124
rect 231762 233112 231768 233124
rect 231820 233112 231826 233164
rect 176010 232976 176016 233028
rect 176068 233016 176074 233028
rect 176470 233016 176476 233028
rect 176068 232988 176476 233016
rect 176068 232976 176074 232988
rect 176470 232976 176476 232988
rect 176528 232976 176534 233028
rect 254578 232500 254584 232552
rect 254636 232540 254642 232552
rect 580166 232540 580172 232552
rect 254636 232512 580172 232540
rect 254636 232500 254642 232512
rect 580166 232500 580172 232512
rect 580224 232500 580230 232552
rect 97258 231752 97264 231804
rect 97316 231792 97322 231804
rect 97902 231792 97908 231804
rect 97316 231764 97908 231792
rect 97316 231752 97322 231764
rect 97902 231752 97908 231764
rect 97960 231752 97966 231804
rect 184382 231752 184388 231804
rect 184440 231792 184446 231804
rect 261018 231792 261024 231804
rect 184440 231764 261024 231792
rect 184440 231752 184446 231764
rect 261018 231752 261024 231764
rect 261076 231752 261082 231804
rect 68278 231072 68284 231124
rect 68336 231112 68342 231124
rect 77478 231112 77484 231124
rect 68336 231084 77484 231112
rect 68336 231072 68342 231084
rect 77478 231072 77484 231084
rect 77536 231072 77542 231124
rect 240226 231072 240232 231124
rect 240284 231112 240290 231124
rect 278958 231112 278964 231124
rect 240284 231084 278964 231112
rect 240284 231072 240290 231084
rect 278958 231072 278964 231084
rect 279016 231072 279022 231124
rect 18598 230528 18604 230580
rect 18656 230568 18662 230580
rect 97258 230568 97264 230580
rect 18656 230540 97264 230568
rect 18656 230528 18662 230540
rect 97258 230528 97264 230540
rect 97316 230528 97322 230580
rect 77478 230460 77484 230512
rect 77536 230500 77542 230512
rect 182174 230500 182180 230512
rect 77536 230472 182180 230500
rect 77536 230460 77542 230472
rect 182174 230460 182180 230472
rect 182232 230500 182238 230512
rect 182910 230500 182916 230512
rect 182232 230472 182916 230500
rect 182232 230460 182238 230472
rect 182910 230460 182916 230472
rect 182968 230460 182974 230512
rect 67266 230392 67272 230444
rect 67324 230432 67330 230444
rect 108390 230432 108396 230444
rect 67324 230404 108396 230432
rect 67324 230392 67330 230404
rect 108390 230392 108396 230404
rect 108448 230392 108454 230444
rect 133230 230392 133236 230444
rect 133288 230432 133294 230444
rect 277394 230432 277400 230444
rect 133288 230404 277400 230432
rect 133288 230392 133294 230404
rect 277394 230392 277400 230404
rect 277452 230392 277458 230444
rect 89714 229712 89720 229764
rect 89772 229752 89778 229764
rect 111058 229752 111064 229764
rect 89772 229724 111064 229752
rect 89772 229712 89778 229724
rect 111058 229712 111064 229724
rect 111116 229752 111122 229764
rect 118694 229752 118700 229764
rect 111116 229724 118700 229752
rect 111116 229712 111122 229724
rect 118694 229712 118700 229724
rect 118752 229712 118758 229764
rect 218698 229712 218704 229764
rect 218756 229752 218762 229764
rect 222194 229752 222200 229764
rect 218756 229724 222200 229752
rect 218756 229712 218762 229724
rect 222194 229712 222200 229724
rect 222252 229712 222258 229764
rect 253198 229712 253204 229764
rect 253256 229752 253262 229764
rect 260834 229752 260840 229764
rect 253256 229724 260840 229752
rect 253256 229712 253262 229724
rect 260834 229712 260840 229724
rect 260892 229712 260898 229764
rect 112438 229032 112444 229084
rect 112496 229072 112502 229084
rect 215294 229072 215300 229084
rect 112496 229044 215300 229072
rect 112496 229032 112502 229044
rect 215294 229032 215300 229044
rect 215352 229032 215358 229084
rect 215294 228692 215300 228744
rect 215352 228732 215358 228744
rect 215938 228732 215944 228744
rect 215352 228704 215944 228732
rect 215352 228692 215358 228704
rect 215938 228692 215944 228704
rect 215996 228692 216002 228744
rect 80054 228352 80060 228404
rect 80112 228392 80118 228404
rect 111794 228392 111800 228404
rect 80112 228364 111800 228392
rect 80112 228352 80118 228364
rect 111794 228352 111800 228364
rect 111852 228392 111858 228404
rect 119430 228392 119436 228404
rect 111852 228364 119436 228392
rect 111852 228352 111858 228364
rect 119430 228352 119436 228364
rect 119488 228352 119494 228404
rect 149882 228352 149888 228404
rect 149940 228392 149946 228404
rect 238846 228392 238852 228404
rect 149940 228364 238852 228392
rect 149940 228352 149946 228364
rect 238846 228352 238852 228364
rect 238904 228392 238910 228404
rect 240042 228392 240048 228404
rect 238904 228364 240048 228392
rect 238904 228352 238910 228364
rect 240042 228352 240048 228364
rect 240100 228352 240106 228404
rect 262858 228352 262864 228404
rect 262916 228392 262922 228404
rect 270770 228392 270776 228404
rect 262916 228364 270776 228392
rect 262916 228352 262922 228364
rect 270770 228352 270776 228364
rect 270828 228352 270834 228404
rect 3418 227672 3424 227724
rect 3476 227712 3482 227724
rect 92474 227712 92480 227724
rect 3476 227684 92480 227712
rect 3476 227672 3482 227684
rect 92474 227672 92480 227684
rect 92532 227672 92538 227724
rect 148502 227060 148508 227112
rect 148560 227100 148566 227112
rect 237374 227100 237380 227112
rect 148560 227072 237380 227100
rect 148560 227060 148566 227072
rect 237374 227060 237380 227072
rect 237432 227060 237438 227112
rect 258810 227060 258816 227112
rect 258868 227100 258874 227112
rect 274818 227100 274824 227112
rect 258868 227072 274824 227100
rect 258868 227060 258874 227072
rect 274818 227060 274824 227072
rect 274876 227060 274882 227112
rect 65794 226992 65800 227044
rect 65852 227032 65858 227044
rect 260926 227032 260932 227044
rect 65852 227004 260932 227032
rect 65852 226992 65858 227004
rect 260926 226992 260932 227004
rect 260984 226992 260990 227044
rect 92474 226312 92480 226364
rect 92532 226352 92538 226364
rect 93118 226352 93124 226364
rect 92532 226324 93124 226352
rect 92532 226312 92538 226324
rect 93118 226312 93124 226324
rect 93176 226312 93182 226364
rect 236086 225632 236092 225684
rect 236144 225672 236150 225684
rect 283006 225672 283012 225684
rect 236144 225644 283012 225672
rect 236144 225632 236150 225644
rect 283006 225632 283012 225644
rect 283064 225672 283070 225684
rect 283064 225644 287054 225672
rect 283064 225632 283070 225644
rect 65978 225564 65984 225616
rect 66036 225604 66042 225616
rect 169110 225604 169116 225616
rect 66036 225576 169116 225604
rect 66036 225564 66042 225576
rect 169110 225564 169116 225576
rect 169168 225564 169174 225616
rect 213178 225564 213184 225616
rect 213236 225604 213242 225616
rect 263870 225604 263876 225616
rect 213236 225576 263876 225604
rect 213236 225564 213242 225576
rect 263870 225564 263876 225576
rect 263928 225564 263934 225616
rect 287026 225604 287054 225644
rect 580258 225604 580264 225616
rect 287026 225576 580264 225604
rect 580258 225564 580264 225576
rect 580316 225564 580322 225616
rect 170766 224272 170772 224324
rect 170824 224312 170830 224324
rect 170824 224284 200114 224312
rect 170824 224272 170830 224284
rect 53558 224204 53564 224256
rect 53616 224244 53622 224256
rect 177390 224244 177396 224256
rect 53616 224216 177396 224244
rect 53616 224204 53622 224216
rect 177390 224204 177396 224216
rect 177448 224204 177454 224256
rect 200086 224244 200114 224284
rect 240778 224272 240784 224324
rect 240836 224312 240842 224324
rect 258166 224312 258172 224324
rect 240836 224284 258172 224312
rect 240836 224272 240842 224284
rect 258166 224272 258172 224284
rect 258224 224272 258230 224324
rect 213914 224244 213920 224256
rect 200086 224216 213920 224244
rect 213914 224204 213920 224216
rect 213972 224244 213978 224256
rect 265618 224244 265624 224256
rect 213972 224216 265624 224244
rect 213972 224204 213978 224216
rect 265618 224204 265624 224216
rect 265676 224204 265682 224256
rect 88334 223524 88340 223576
rect 88392 223564 88398 223576
rect 121454 223564 121460 223576
rect 88392 223536 121460 223564
rect 88392 223524 88398 223536
rect 121454 223524 121460 223536
rect 121512 223524 121518 223576
rect 152550 222912 152556 222964
rect 152608 222952 152614 222964
rect 220814 222952 220820 222964
rect 152608 222924 220820 222952
rect 152608 222912 152614 222924
rect 220814 222912 220820 222924
rect 220872 222952 220878 222964
rect 222102 222952 222108 222964
rect 220872 222924 222108 222952
rect 220872 222912 220878 222924
rect 222102 222912 222108 222924
rect 222160 222912 222166 222964
rect 63218 222844 63224 222896
rect 63276 222884 63282 222896
rect 159450 222884 159456 222896
rect 63276 222856 159456 222884
rect 63276 222844 63282 222856
rect 159450 222844 159456 222856
rect 159508 222844 159514 222896
rect 163682 222844 163688 222896
rect 163740 222884 163746 222896
rect 237374 222884 237380 222896
rect 163740 222856 237380 222884
rect 163740 222844 163746 222856
rect 237374 222844 237380 222856
rect 237432 222844 237438 222896
rect 67358 222096 67364 222148
rect 67416 222136 67422 222148
rect 269298 222136 269304 222148
rect 67416 222108 269304 222136
rect 67416 222096 67422 222108
rect 269298 222096 269304 222108
rect 269356 222096 269362 222148
rect 222838 221416 222844 221468
rect 222896 221456 222902 221468
rect 254118 221456 254124 221468
rect 222896 221428 254124 221456
rect 222896 221416 222902 221428
rect 254118 221416 254124 221428
rect 254176 221416 254182 221468
rect 171042 220804 171048 220856
rect 171100 220844 171106 220856
rect 173342 220844 173348 220856
rect 171100 220816 173348 220844
rect 171100 220804 171106 220816
rect 173342 220804 173348 220816
rect 173400 220804 173406 220856
rect 113818 220736 113824 220788
rect 113876 220776 113882 220788
rect 236086 220776 236092 220788
rect 113876 220748 236092 220776
rect 113876 220736 113882 220748
rect 236086 220736 236092 220748
rect 236144 220736 236150 220788
rect 100110 220056 100116 220108
rect 100168 220096 100174 220108
rect 277486 220096 277492 220108
rect 100168 220068 277492 220096
rect 100168 220056 100174 220068
rect 277486 220056 277492 220068
rect 277544 220096 277550 220108
rect 277670 220096 277676 220108
rect 277544 220068 277676 220096
rect 277544 220056 277550 220068
rect 277670 220056 277676 220068
rect 277728 220056 277734 220108
rect 288434 219376 288440 219428
rect 288492 219416 288498 219428
rect 579890 219416 579896 219428
rect 288492 219388 579896 219416
rect 288492 219376 288498 219388
rect 579890 219376 579896 219388
rect 579948 219376 579954 219428
rect 77938 218764 77944 218816
rect 77996 218804 78002 218816
rect 87598 218804 87604 218816
rect 77996 218776 87604 218804
rect 77996 218764 78002 218776
rect 87598 218764 87604 218776
rect 87656 218764 87662 218816
rect 103422 218764 103428 218816
rect 103480 218804 103486 218816
rect 184198 218804 184204 218816
rect 103480 218776 184204 218804
rect 103480 218764 103486 218776
rect 184198 218764 184204 218776
rect 184256 218764 184262 218816
rect 60642 218696 60648 218748
rect 60700 218736 60706 218748
rect 156690 218736 156696 218748
rect 60700 218708 156696 218736
rect 60700 218696 60706 218708
rect 156690 218696 156696 218708
rect 156748 218736 156754 218748
rect 254578 218736 254584 218748
rect 156748 218708 254584 218736
rect 156748 218696 156754 218708
rect 254578 218696 254584 218708
rect 254636 218696 254642 218748
rect 104250 217948 104256 218000
rect 104308 217988 104314 218000
rect 240778 217988 240784 218000
rect 104308 217960 240784 217988
rect 104308 217948 104314 217960
rect 240778 217948 240784 217960
rect 240836 217948 240842 218000
rect 158622 217880 158628 217932
rect 158680 217920 158686 217932
rect 272150 217920 272156 217932
rect 158680 217892 272156 217920
rect 158680 217880 158686 217892
rect 272150 217880 272156 217892
rect 272208 217880 272214 217932
rect 48130 217268 48136 217320
rect 48188 217308 48194 217320
rect 77294 217308 77300 217320
rect 48188 217280 77300 217308
rect 48188 217268 48194 217280
rect 77294 217268 77300 217280
rect 77352 217268 77358 217320
rect 88242 217268 88248 217320
rect 88300 217308 88306 217320
rect 154482 217308 154488 217320
rect 88300 217280 154488 217308
rect 88300 217268 88306 217280
rect 154482 217268 154488 217280
rect 154540 217268 154546 217320
rect 118602 215976 118608 216028
rect 118660 216016 118666 216028
rect 185762 216016 185768 216028
rect 118660 215988 185768 216016
rect 118660 215976 118666 215988
rect 185762 215976 185768 215988
rect 185820 215976 185826 216028
rect 187050 215976 187056 216028
rect 187108 216016 187114 216028
rect 251818 216016 251824 216028
rect 187108 215988 251824 216016
rect 187108 215976 187114 215988
rect 251818 215976 251824 215988
rect 251876 215976 251882 216028
rect 177390 215908 177396 215960
rect 177448 215948 177454 215960
rect 250438 215948 250444 215960
rect 177448 215920 250444 215948
rect 177448 215908 177454 215920
rect 250438 215908 250444 215920
rect 250496 215948 250502 215960
rect 259638 215948 259644 215960
rect 250496 215920 259644 215948
rect 250496 215908 250502 215920
rect 259638 215908 259644 215920
rect 259696 215908 259702 215960
rect 91094 215228 91100 215280
rect 91152 215268 91158 215280
rect 170490 215268 170496 215280
rect 91152 215240 170496 215268
rect 91152 215228 91158 215240
rect 170490 215228 170496 215240
rect 170548 215268 170554 215280
rect 227714 215268 227720 215280
rect 170548 215240 227720 215268
rect 170548 215228 170554 215240
rect 227714 215228 227720 215240
rect 227772 215228 227778 215280
rect 227714 214752 227720 214804
rect 227772 214792 227778 214804
rect 228450 214792 228456 214804
rect 227772 214764 228456 214792
rect 227772 214752 227778 214764
rect 228450 214752 228456 214764
rect 228508 214752 228514 214804
rect 100202 214548 100208 214600
rect 100260 214588 100266 214600
rect 267826 214588 267832 214600
rect 100260 214560 267832 214588
rect 100260 214548 100266 214560
rect 267826 214548 267832 214560
rect 267884 214548 267890 214600
rect 98086 213868 98092 213920
rect 98144 213908 98150 213920
rect 98730 213908 98736 213920
rect 98144 213880 98736 213908
rect 98144 213868 98150 213880
rect 98730 213868 98736 213880
rect 98788 213868 98794 213920
rect 93854 213256 93860 213308
rect 93912 213296 93918 213308
rect 121546 213296 121552 213308
rect 93912 213268 121552 213296
rect 93912 213256 93918 213268
rect 121546 213256 121552 213268
rect 121604 213256 121610 213308
rect 98730 213188 98736 213240
rect 98788 213228 98794 213240
rect 206370 213228 206376 213240
rect 98788 213200 206376 213228
rect 98788 213188 98794 213200
rect 206370 213188 206376 213200
rect 206428 213188 206434 213240
rect 121546 212508 121552 212560
rect 121604 212548 121610 212560
rect 259546 212548 259552 212560
rect 121604 212520 259552 212548
rect 121604 212508 121610 212520
rect 259546 212508 259552 212520
rect 259604 212508 259610 212560
rect 254578 211760 254584 211812
rect 254636 211800 254642 211812
rect 267918 211800 267924 211812
rect 254636 211772 267924 211800
rect 254636 211760 254642 211772
rect 267918 211760 267924 211772
rect 267976 211760 267982 211812
rect 96614 211080 96620 211132
rect 96672 211120 96678 211132
rect 102318 211120 102324 211132
rect 96672 211092 102324 211120
rect 96672 211080 96678 211092
rect 102318 211080 102324 211092
rect 102376 211080 102382 211132
rect 154482 211080 154488 211132
rect 154540 211120 154546 211132
rect 224954 211120 224960 211132
rect 154540 211092 224960 211120
rect 154540 211080 154546 211092
rect 224954 211080 224960 211092
rect 225012 211080 225018 211132
rect 53558 210400 53564 210452
rect 53616 210440 53622 210452
rect 73246 210440 73252 210452
rect 53616 210412 73252 210440
rect 53616 210400 53622 210412
rect 73246 210400 73252 210412
rect 73304 210400 73310 210452
rect 88242 210400 88248 210452
rect 88300 210440 88306 210452
rect 102134 210440 102140 210452
rect 88300 210412 102140 210440
rect 88300 210400 88306 210412
rect 102134 210400 102140 210412
rect 102192 210400 102198 210452
rect 102318 209788 102324 209840
rect 102376 209828 102382 209840
rect 270586 209828 270592 209840
rect 102376 209800 270592 209828
rect 102376 209788 102382 209800
rect 270586 209788 270592 209800
rect 270644 209788 270650 209840
rect 102226 209720 102232 209772
rect 102284 209760 102290 209772
rect 263686 209760 263692 209772
rect 102284 209732 263692 209760
rect 102284 209720 102290 209732
rect 263686 209720 263692 209732
rect 263744 209720 263750 209772
rect 88150 209040 88156 209092
rect 88208 209080 88214 209092
rect 120074 209080 120080 209092
rect 88208 209052 120080 209080
rect 88208 209040 88214 209052
rect 120074 209040 120080 209052
rect 120132 209040 120138 209092
rect 224218 209040 224224 209092
rect 224276 209080 224282 209092
rect 253934 209080 253940 209092
rect 224276 209052 253940 209080
rect 224276 209040 224282 209052
rect 253934 209040 253940 209052
rect 253992 209040 253998 209092
rect 98638 208360 98644 208412
rect 98696 208400 98702 208412
rect 102226 208400 102232 208412
rect 98696 208372 102232 208400
rect 98696 208360 98702 208372
rect 102226 208360 102232 208372
rect 102284 208360 102290 208412
rect 175182 208360 175188 208412
rect 175240 208400 175246 208412
rect 180058 208400 180064 208412
rect 175240 208372 180064 208400
rect 175240 208360 175246 208372
rect 180058 208360 180064 208372
rect 180116 208360 180122 208412
rect 86954 207680 86960 207732
rect 87012 207720 87018 207732
rect 110506 207720 110512 207732
rect 87012 207692 110512 207720
rect 87012 207680 87018 207692
rect 110506 207680 110512 207692
rect 110564 207680 110570 207732
rect 97258 207612 97264 207664
rect 97316 207652 97322 207664
rect 266446 207652 266452 207664
rect 97316 207624 266452 207652
rect 97316 207612 97322 207624
rect 266446 207612 266452 207624
rect 266504 207612 266510 207664
rect 110506 207000 110512 207052
rect 110564 207040 110570 207052
rect 256694 207040 256700 207052
rect 110564 207012 256700 207040
rect 110564 207000 110570 207012
rect 256694 207000 256700 207012
rect 256752 207000 256758 207052
rect 79962 206252 79968 206304
rect 80020 206292 80026 206304
rect 91094 206292 91100 206304
rect 80020 206264 91100 206292
rect 80020 206252 80026 206264
rect 91094 206252 91100 206264
rect 91152 206252 91158 206304
rect 93118 206252 93124 206304
rect 93176 206292 93182 206304
rect 274634 206292 274640 206304
rect 93176 206264 274640 206292
rect 93176 206252 93182 206264
rect 274634 206252 274640 206264
rect 274692 206252 274698 206304
rect 91094 205640 91100 205692
rect 91152 205680 91158 205692
rect 92382 205680 92388 205692
rect 91152 205652 92388 205680
rect 91152 205640 91158 205652
rect 92382 205640 92388 205652
rect 92440 205680 92446 205692
rect 176010 205680 176016 205692
rect 92440 205652 176016 205680
rect 92440 205640 92446 205652
rect 176010 205640 176016 205652
rect 176068 205640 176074 205692
rect 95234 204892 95240 204944
rect 95292 204932 95298 204944
rect 95878 204932 95884 204944
rect 95292 204904 95884 204932
rect 95292 204892 95298 204904
rect 95878 204892 95884 204904
rect 95936 204932 95942 204944
rect 262214 204932 262220 204944
rect 95936 204904 262220 204932
rect 95936 204892 95942 204904
rect 262214 204892 262220 204904
rect 262272 204932 262278 204944
rect 262582 204932 262588 204944
rect 262272 204904 262588 204932
rect 262272 204892 262278 204904
rect 262582 204892 262588 204904
rect 262640 204892 262646 204944
rect 3418 204212 3424 204264
rect 3476 204252 3482 204264
rect 7558 204252 7564 204264
rect 3476 204224 7564 204252
rect 3476 204212 3482 204224
rect 7558 204212 7564 204224
rect 7616 204212 7622 204264
rect 158070 204212 158076 204264
rect 158128 204252 158134 204264
rect 271966 204252 271972 204264
rect 158128 204224 271972 204252
rect 158128 204212 158134 204224
rect 271966 204212 271972 204224
rect 272024 204212 272030 204264
rect 169110 203532 169116 203584
rect 169168 203572 169174 203584
rect 178862 203572 178868 203584
rect 169168 203544 178868 203572
rect 169168 203532 169174 203544
rect 178862 203532 178868 203544
rect 178920 203532 178926 203584
rect 99374 202784 99380 202836
rect 99432 202824 99438 202836
rect 100202 202824 100208 202836
rect 99432 202796 100208 202824
rect 99432 202784 99438 202796
rect 100202 202784 100208 202796
rect 100260 202784 100266 202836
rect 147122 202784 147128 202836
rect 147180 202824 147186 202836
rect 241514 202824 241520 202836
rect 147180 202796 241520 202824
rect 147180 202784 147186 202796
rect 241514 202784 241520 202796
rect 241572 202784 241578 202836
rect 3234 202104 3240 202156
rect 3292 202144 3298 202156
rect 99374 202144 99380 202156
rect 3292 202116 99380 202144
rect 3292 202104 3298 202116
rect 99374 202104 99380 202116
rect 99432 202104 99438 202156
rect 188338 201424 188344 201476
rect 188396 201464 188402 201476
rect 188890 201464 188896 201476
rect 188396 201436 188896 201464
rect 188396 201424 188402 201436
rect 188890 201424 188896 201436
rect 188948 201464 188954 201476
rect 257338 201464 257344 201476
rect 188948 201436 257344 201464
rect 188948 201424 188954 201436
rect 257338 201424 257344 201436
rect 257396 201424 257402 201476
rect 192938 199384 192944 199436
rect 192996 199424 193002 199436
rect 249058 199424 249064 199436
rect 192996 199396 249064 199424
rect 192996 199384 193002 199396
rect 249058 199384 249064 199396
rect 249116 199384 249122 199436
rect 117958 197276 117964 197328
rect 118016 197316 118022 197328
rect 223574 197316 223580 197328
rect 118016 197288 223580 197316
rect 118016 197276 118022 197288
rect 223574 197276 223580 197288
rect 223632 197276 223638 197328
rect 223574 196664 223580 196716
rect 223632 196704 223638 196716
rect 224218 196704 224224 196716
rect 223632 196676 224224 196704
rect 223632 196664 223638 196676
rect 224218 196664 224224 196676
rect 224276 196664 224282 196716
rect 20622 196596 20628 196648
rect 20680 196636 20686 196648
rect 120718 196636 120724 196648
rect 20680 196608 120724 196636
rect 20680 196596 20686 196608
rect 120718 196596 120724 196608
rect 120776 196596 120782 196648
rect 233878 196596 233884 196648
rect 233936 196636 233942 196648
rect 244366 196636 244372 196648
rect 233936 196608 244372 196636
rect 233936 196596 233942 196608
rect 244366 196596 244372 196608
rect 244424 196596 244430 196648
rect 108298 195916 108304 195968
rect 108356 195956 108362 195968
rect 220906 195956 220912 195968
rect 108356 195928 220912 195956
rect 108356 195916 108362 195928
rect 220906 195916 220912 195928
rect 220964 195956 220970 195968
rect 221826 195956 221832 195968
rect 220964 195928 221832 195956
rect 220964 195916 220970 195928
rect 221826 195916 221832 195928
rect 221884 195916 221890 195968
rect 84930 195236 84936 195288
rect 84988 195276 84994 195288
rect 106274 195276 106280 195288
rect 84988 195248 106280 195276
rect 84988 195236 84994 195248
rect 106274 195236 106280 195248
rect 106332 195236 106338 195288
rect 240778 194556 240784 194608
rect 240836 194596 240842 194608
rect 580166 194596 580172 194608
rect 240836 194568 580172 194596
rect 240836 194556 240842 194568
rect 580166 194556 580172 194568
rect 580224 194556 580230 194608
rect 44082 193808 44088 193860
rect 44140 193848 44146 193860
rect 149790 193848 149796 193860
rect 44140 193820 149796 193848
rect 44140 193808 44146 193820
rect 149790 193808 149796 193820
rect 149848 193808 149854 193860
rect 188982 193808 188988 193860
rect 189040 193848 189046 193860
rect 574738 193848 574744 193860
rect 189040 193820 574744 193848
rect 189040 193808 189046 193820
rect 574738 193808 574744 193820
rect 574796 193808 574802 193860
rect 84838 192516 84844 192568
rect 84896 192556 84902 192568
rect 115382 192556 115388 192568
rect 84896 192528 115388 192556
rect 84896 192516 84902 192528
rect 115382 192516 115388 192528
rect 115440 192516 115446 192568
rect 3878 192448 3884 192500
rect 3936 192488 3942 192500
rect 133138 192488 133144 192500
rect 3936 192460 133144 192488
rect 3936 192448 3942 192460
rect 133138 192448 133144 192460
rect 133196 192448 133202 192500
rect 229830 192448 229836 192500
rect 229888 192488 229894 192500
rect 266538 192488 266544 192500
rect 229888 192460 266544 192488
rect 229888 192448 229894 192460
rect 266538 192448 266544 192460
rect 266596 192448 266602 192500
rect 221826 191768 221832 191820
rect 221884 191808 221890 191820
rect 225138 191808 225144 191820
rect 221884 191780 225144 191808
rect 221884 191768 221890 191780
rect 225138 191768 225144 191780
rect 225196 191768 225202 191820
rect 59262 191088 59268 191140
rect 59320 191128 59326 191140
rect 173250 191128 173256 191140
rect 59320 191100 173256 191128
rect 59320 191088 59326 191100
rect 173250 191088 173256 191100
rect 173308 191088 173314 191140
rect 190362 191088 190368 191140
rect 190420 191128 190426 191140
rect 263778 191128 263784 191140
rect 190420 191100 263784 191128
rect 190420 191088 190426 191100
rect 263778 191088 263784 191100
rect 263836 191088 263842 191140
rect 3418 188980 3424 189032
rect 3476 189020 3482 189032
rect 18598 189020 18604 189032
rect 3476 188992 18604 189020
rect 3476 188980 3482 188992
rect 18598 188980 18604 188992
rect 18656 188980 18662 189032
rect 27522 188300 27528 188352
rect 27580 188340 27586 188352
rect 148410 188340 148416 188352
rect 27580 188312 148416 188340
rect 27580 188300 27586 188312
rect 148410 188300 148416 188312
rect 148468 188300 148474 188352
rect 193766 188300 193772 188352
rect 193824 188340 193830 188352
rect 235994 188340 236000 188352
rect 193824 188312 236000 188340
rect 193824 188300 193830 188312
rect 235994 188300 236000 188312
rect 236052 188300 236058 188352
rect 87598 187008 87604 187060
rect 87656 187048 87662 187060
rect 104158 187048 104164 187060
rect 87656 187020 104164 187048
rect 87656 187008 87662 187020
rect 104158 187008 104164 187020
rect 104216 187008 104222 187060
rect 5442 186940 5448 186992
rect 5500 186980 5506 186992
rect 155310 186980 155316 186992
rect 5500 186952 155316 186980
rect 5500 186940 5506 186952
rect 155310 186940 155316 186952
rect 155368 186940 155374 186992
rect 184290 186940 184296 186992
rect 184348 186980 184354 186992
rect 200758 186980 200764 186992
rect 184348 186952 200764 186980
rect 184348 186940 184354 186952
rect 200758 186940 200764 186952
rect 200816 186940 200822 186992
rect 240778 186940 240784 186992
rect 240836 186980 240842 186992
rect 276290 186980 276296 186992
rect 240836 186952 276296 186980
rect 240836 186940 240842 186952
rect 276290 186940 276296 186952
rect 276348 186940 276354 186992
rect 17218 185580 17224 185632
rect 17276 185620 17282 185632
rect 144178 185620 144184 185632
rect 17276 185592 144184 185620
rect 17276 185580 17282 185592
rect 144178 185580 144184 185592
rect 144236 185580 144242 185632
rect 213178 185580 213184 185632
rect 213236 185620 213242 185632
rect 235258 185620 235264 185632
rect 213236 185592 235264 185620
rect 213236 185580 213242 185592
rect 235258 185580 235264 185592
rect 235316 185580 235322 185632
rect 86862 184220 86868 184272
rect 86920 184260 86926 184272
rect 97350 184260 97356 184272
rect 86920 184232 97356 184260
rect 86920 184220 86926 184232
rect 97350 184220 97356 184232
rect 97408 184220 97414 184272
rect 28902 184152 28908 184204
rect 28960 184192 28966 184204
rect 189718 184192 189724 184204
rect 28960 184164 189724 184192
rect 28960 184152 28966 184164
rect 189718 184152 189724 184164
rect 189776 184152 189782 184204
rect 88978 182792 88984 182844
rect 89036 182832 89042 182844
rect 120166 182832 120172 182844
rect 89036 182804 120172 182832
rect 89036 182792 89042 182804
rect 120166 182792 120172 182804
rect 120224 182792 120230 182844
rect 133138 181432 133144 181484
rect 133196 181472 133202 181484
rect 206278 181472 206284 181484
rect 133196 181444 206284 181472
rect 133196 181432 133202 181444
rect 206278 181432 206284 181444
rect 206336 181432 206342 181484
rect 91002 180072 91008 180124
rect 91060 180112 91066 180124
rect 117314 180112 117320 180124
rect 91060 180084 117320 180112
rect 91060 180072 91066 180084
rect 117314 180072 117320 180084
rect 117372 180072 117378 180124
rect 99190 179392 99196 179444
rect 99248 179432 99254 179444
rect 226426 179432 226432 179444
rect 99248 179404 226432 179432
rect 99248 179392 99254 179404
rect 226426 179392 226432 179404
rect 226484 179392 226490 179444
rect 92290 178644 92296 178696
rect 92348 178684 92354 178696
rect 118694 178684 118700 178696
rect 92348 178656 118700 178684
rect 92348 178644 92354 178656
rect 118694 178644 118700 178656
rect 118752 178644 118758 178696
rect 238018 178644 238024 178696
rect 238076 178684 238082 178696
rect 238662 178684 238668 178696
rect 238076 178656 238668 178684
rect 238076 178644 238082 178656
rect 238662 178644 238668 178656
rect 238720 178684 238726 178696
rect 580166 178684 580172 178696
rect 238720 178656 580172 178684
rect 238720 178644 238726 178656
rect 580166 178644 580172 178656
rect 580224 178644 580230 178696
rect 71038 178032 71044 178084
rect 71096 178072 71102 178084
rect 159542 178072 159548 178084
rect 71096 178044 159548 178072
rect 71096 178032 71102 178044
rect 159542 178032 159548 178044
rect 159600 178032 159606 178084
rect 75362 177352 75368 177404
rect 75420 177392 75426 177404
rect 128998 177392 129004 177404
rect 75420 177364 129004 177392
rect 75420 177352 75426 177364
rect 128998 177352 129004 177364
rect 129056 177352 129062 177404
rect 197998 177352 198004 177404
rect 198056 177392 198062 177404
rect 226702 177392 226708 177404
rect 198056 177364 226708 177392
rect 198056 177352 198062 177364
rect 226702 177352 226708 177364
rect 226760 177352 226766 177404
rect 80790 177284 80796 177336
rect 80848 177324 80854 177336
rect 106458 177324 106464 177336
rect 80848 177296 106464 177324
rect 80848 177284 80854 177296
rect 106458 177284 106464 177296
rect 106516 177324 106522 177336
rect 219526 177324 219532 177336
rect 106516 177296 219532 177324
rect 106516 177284 106522 177296
rect 219526 177284 219532 177296
rect 219584 177324 219590 177336
rect 219710 177324 219716 177336
rect 219584 177296 219716 177324
rect 219584 177284 219590 177296
rect 219710 177284 219716 177296
rect 219768 177284 219774 177336
rect 154022 175312 154028 175364
rect 154080 175352 154086 175364
rect 204254 175352 204260 175364
rect 154080 175324 204260 175352
rect 154080 175312 154086 175324
rect 204254 175312 204260 175324
rect 204312 175352 204318 175364
rect 204898 175352 204904 175364
rect 204312 175324 204904 175352
rect 204312 175312 204318 175324
rect 204898 175312 204904 175324
rect 204956 175312 204962 175364
rect 89714 175244 89720 175296
rect 89772 175284 89778 175296
rect 219434 175284 219440 175296
rect 89772 175256 219440 175284
rect 89772 175244 89778 175256
rect 219434 175244 219440 175256
rect 219492 175284 219498 175296
rect 220078 175284 220084 175296
rect 219492 175256 220084 175284
rect 219492 175244 219498 175256
rect 220078 175244 220084 175256
rect 220136 175244 220142 175296
rect 85574 174496 85580 174548
rect 85632 174536 85638 174548
rect 195974 174536 195980 174548
rect 85632 174508 195980 174536
rect 85632 174496 85638 174508
rect 195974 174496 195980 174508
rect 196032 174536 196038 174548
rect 215938 174536 215944 174548
rect 196032 174508 215944 174536
rect 196032 174496 196038 174508
rect 215938 174496 215944 174508
rect 215996 174496 216002 174548
rect 153930 173884 153936 173936
rect 153988 173924 153994 173936
rect 222194 173924 222200 173936
rect 153988 173896 222200 173924
rect 153988 173884 153994 173896
rect 222194 173884 222200 173896
rect 222252 173924 222258 173936
rect 222930 173924 222936 173936
rect 222252 173896 222936 173924
rect 222252 173884 222258 173896
rect 222930 173884 222936 173896
rect 222988 173884 222994 173936
rect 80698 173136 80704 173188
rect 80756 173176 80762 173188
rect 160922 173176 160928 173188
rect 80756 173148 160928 173176
rect 80756 173136 80762 173148
rect 160922 173136 160928 173148
rect 160980 173176 160986 173188
rect 195238 173176 195244 173188
rect 160980 173148 195244 173176
rect 160980 173136 160986 173148
rect 195238 173136 195244 173148
rect 195296 173136 195302 173188
rect 206370 173136 206376 173188
rect 206428 173176 206434 173188
rect 227806 173176 227812 173188
rect 206428 173148 227812 173176
rect 206428 173136 206434 173148
rect 227806 173136 227812 173148
rect 227864 173136 227870 173188
rect 75914 171776 75920 171828
rect 75972 171816 75978 171828
rect 156598 171816 156604 171828
rect 75972 171788 156604 171816
rect 75972 171776 75978 171788
rect 156598 171776 156604 171788
rect 156656 171816 156662 171828
rect 202874 171816 202880 171828
rect 156656 171788 202880 171816
rect 156656 171776 156662 171788
rect 202874 171776 202880 171788
rect 202932 171776 202938 171828
rect 104618 171096 104624 171148
rect 104676 171136 104682 171148
rect 210418 171136 210424 171148
rect 104676 171108 210424 171136
rect 104676 171096 104682 171108
rect 210418 171096 210424 171108
rect 210476 171096 210482 171148
rect 211154 171096 211160 171148
rect 211212 171136 211218 171148
rect 317414 171136 317420 171148
rect 211212 171108 317420 171136
rect 211212 171096 211218 171108
rect 317414 171096 317420 171108
rect 317472 171096 317478 171148
rect 189718 170348 189724 170400
rect 189776 170388 189782 170400
rect 250438 170388 250444 170400
rect 189776 170360 250444 170388
rect 189776 170348 189782 170360
rect 250438 170348 250444 170360
rect 250496 170388 250502 170400
rect 582742 170388 582748 170400
rect 250496 170360 582748 170388
rect 250496 170348 250502 170360
rect 582742 170348 582748 170360
rect 582800 170348 582806 170400
rect 67818 169736 67824 169788
rect 67876 169776 67882 169788
rect 68554 169776 68560 169788
rect 67876 169748 68560 169776
rect 67876 169736 67882 169748
rect 68554 169736 68560 169748
rect 68612 169776 68618 169788
rect 194502 169776 194508 169788
rect 68612 169748 194508 169776
rect 68612 169736 68618 169748
rect 194502 169736 194508 169748
rect 194560 169736 194566 169788
rect 81526 168988 81532 169040
rect 81584 169028 81590 169040
rect 154022 169028 154028 169040
rect 81584 169000 154028 169028
rect 81584 168988 81590 169000
rect 154022 168988 154028 169000
rect 154080 168988 154086 169040
rect 154482 168988 154488 169040
rect 154540 169028 154546 169040
rect 162302 169028 162308 169040
rect 154540 169000 162308 169028
rect 154540 168988 154546 169000
rect 162302 168988 162308 169000
rect 162360 169028 162366 169040
rect 204990 169028 204996 169040
rect 162360 169000 204996 169028
rect 162360 168988 162366 169000
rect 204990 168988 204996 169000
rect 205048 168988 205054 169040
rect 193858 168376 193864 168428
rect 193916 168416 193922 168428
rect 194502 168416 194508 168428
rect 193916 168388 194508 168416
rect 193916 168376 193922 168388
rect 194502 168376 194508 168388
rect 194560 168416 194566 168428
rect 194560 168388 234108 168416
rect 194560 168376 194566 168388
rect 166442 168308 166448 168360
rect 166500 168348 166506 168360
rect 211154 168348 211160 168360
rect 166500 168320 211160 168348
rect 166500 168308 166506 168320
rect 211154 168308 211160 168320
rect 211212 168308 211218 168360
rect 234080 168348 234108 168388
rect 234522 168348 234528 168360
rect 234080 168320 234528 168348
rect 234522 168308 234528 168320
rect 234580 168348 234586 168360
rect 243538 168348 243544 168360
rect 234580 168320 243544 168348
rect 234580 168308 234586 168320
rect 243538 168308 243544 168320
rect 243596 168308 243602 168360
rect 82906 167628 82912 167680
rect 82964 167668 82970 167680
rect 166442 167668 166448 167680
rect 82964 167640 166448 167668
rect 82964 167628 82970 167640
rect 166442 167628 166448 167640
rect 166500 167628 166506 167680
rect 141602 167016 141608 167068
rect 141660 167056 141666 167068
rect 223574 167056 223580 167068
rect 141660 167028 223580 167056
rect 141660 167016 141666 167028
rect 223574 167016 223580 167028
rect 223632 167016 223638 167068
rect 200114 166336 200120 166388
rect 200172 166376 200178 166388
rect 229830 166376 229836 166388
rect 200172 166348 229836 166376
rect 200172 166336 200178 166348
rect 229830 166336 229836 166348
rect 229888 166336 229894 166388
rect 84194 166268 84200 166320
rect 84252 166308 84258 166320
rect 157978 166308 157984 166320
rect 84252 166280 157984 166308
rect 84252 166268 84258 166280
rect 157978 166268 157984 166280
rect 158036 166308 158042 166320
rect 213178 166308 213184 166320
rect 158036 166280 213184 166308
rect 158036 166268 158042 166280
rect 213178 166268 213184 166280
rect 213236 166268 213242 166320
rect 218054 166268 218060 166320
rect 218112 166308 218118 166320
rect 267734 166308 267740 166320
rect 218112 166280 267740 166308
rect 218112 166268 218118 166280
rect 267734 166268 267740 166280
rect 267792 166268 267798 166320
rect 54938 165588 54944 165640
rect 54996 165628 55002 165640
rect 190454 165628 190460 165640
rect 54996 165600 190460 165628
rect 54996 165588 55002 165600
rect 190454 165588 190460 165600
rect 190512 165628 190518 165640
rect 191190 165628 191196 165640
rect 190512 165600 191196 165628
rect 190512 165588 190518 165600
rect 191190 165588 191196 165600
rect 191248 165588 191254 165640
rect 92658 164840 92664 164892
rect 92716 164880 92722 164892
rect 153930 164880 153936 164892
rect 92716 164852 153936 164880
rect 92716 164840 92722 164852
rect 153930 164840 153936 164852
rect 153988 164840 153994 164892
rect 202874 164296 202880 164348
rect 202932 164336 202938 164348
rect 300118 164336 300124 164348
rect 202932 164308 300124 164336
rect 202932 164296 202938 164308
rect 300118 164296 300124 164308
rect 300176 164296 300182 164348
rect 100202 164228 100208 164280
rect 100260 164268 100266 164280
rect 100662 164268 100668 164280
rect 100260 164240 100668 164268
rect 100260 164228 100266 164240
rect 100662 164228 100668 164240
rect 100720 164268 100726 164280
rect 237466 164268 237472 164280
rect 100720 164240 237472 164268
rect 100720 164228 100726 164240
rect 237466 164228 237472 164240
rect 237524 164228 237530 164280
rect 77386 163548 77392 163600
rect 77444 163588 77450 163600
rect 154482 163588 154488 163600
rect 77444 163560 154488 163588
rect 77444 163548 77450 163560
rect 154482 163548 154488 163560
rect 154540 163548 154546 163600
rect 91738 163480 91744 163532
rect 91796 163520 91802 163532
rect 129090 163520 129096 163532
rect 91796 163492 129096 163520
rect 91796 163480 91802 163492
rect 129090 163480 129096 163492
rect 129148 163520 129154 163532
rect 220998 163520 221004 163532
rect 129148 163492 221004 163520
rect 129148 163480 129154 163492
rect 220998 163480 221004 163492
rect 221056 163480 221062 163532
rect 3418 162868 3424 162920
rect 3476 162908 3482 162920
rect 51810 162908 51816 162920
rect 3476 162880 51816 162908
rect 3476 162868 3482 162880
rect 51810 162868 51816 162880
rect 51868 162868 51874 162920
rect 153930 162868 153936 162920
rect 153988 162908 153994 162920
rect 218054 162908 218060 162920
rect 153988 162880 218060 162908
rect 153988 162868 153994 162880
rect 218054 162868 218060 162880
rect 218112 162868 218118 162920
rect 84102 162120 84108 162172
rect 84160 162160 84166 162172
rect 109034 162160 109040 162172
rect 84160 162132 109040 162160
rect 84160 162120 84166 162132
rect 109034 162120 109040 162132
rect 109092 162120 109098 162172
rect 243538 162120 243544 162172
rect 243596 162160 243602 162172
rect 274634 162160 274640 162172
rect 243596 162132 274640 162160
rect 243596 162120 243602 162132
rect 274634 162120 274640 162132
rect 274692 162120 274698 162172
rect 148410 161508 148416 161560
rect 148468 161548 148474 161560
rect 199378 161548 199384 161560
rect 148468 161520 199384 161548
rect 148468 161508 148474 161520
rect 199378 161508 199384 161520
rect 199436 161548 199442 161560
rect 233234 161548 233240 161560
rect 199436 161520 233240 161548
rect 199436 161508 199442 161520
rect 233234 161508 233240 161520
rect 233292 161508 233298 161560
rect 129182 161440 129188 161492
rect 129240 161480 129246 161492
rect 241698 161480 241704 161492
rect 129240 161452 241704 161480
rect 129240 161440 129246 161452
rect 241698 161440 241704 161452
rect 241756 161440 241762 161492
rect 193030 160760 193036 160812
rect 193088 160800 193094 160812
rect 245194 160800 245200 160812
rect 193088 160772 245200 160800
rect 193088 160760 193094 160772
rect 245194 160760 245200 160772
rect 245252 160760 245258 160812
rect 213270 160692 213276 160744
rect 213328 160732 213334 160744
rect 277578 160732 277584 160744
rect 213328 160704 277584 160732
rect 213328 160692 213334 160704
rect 277578 160692 277584 160704
rect 277636 160692 277642 160744
rect 176562 160148 176568 160200
rect 176620 160188 176626 160200
rect 196710 160188 196716 160200
rect 176620 160160 196716 160188
rect 176620 160148 176626 160160
rect 196710 160148 196716 160160
rect 196768 160148 196774 160200
rect 87598 160080 87604 160132
rect 87656 160120 87662 160132
rect 88242 160120 88248 160132
rect 87656 160092 88248 160120
rect 87656 160080 87662 160092
rect 88242 160080 88248 160092
rect 88300 160120 88306 160132
rect 182082 160120 182088 160132
rect 88300 160092 182088 160120
rect 88300 160080 88306 160092
rect 182082 160080 182088 160092
rect 182140 160080 182146 160132
rect 72970 159332 72976 159384
rect 73028 159372 73034 159384
rect 176562 159372 176568 159384
rect 73028 159344 176568 159372
rect 73028 159332 73034 159344
rect 176562 159332 176568 159344
rect 176620 159332 176626 159384
rect 229830 159332 229836 159384
rect 229888 159372 229894 159384
rect 287698 159372 287704 159384
rect 229888 159344 287704 159372
rect 229888 159332 229894 159344
rect 287698 159332 287704 159344
rect 287756 159332 287762 159384
rect 194594 158788 194600 158840
rect 194652 158828 194658 158840
rect 195238 158828 195244 158840
rect 194652 158800 195244 158828
rect 194652 158788 194658 158800
rect 195238 158788 195244 158800
rect 195296 158828 195302 158840
rect 250438 158828 250444 158840
rect 195296 158800 250444 158828
rect 195296 158788 195302 158800
rect 250438 158788 250444 158800
rect 250496 158788 250502 158840
rect 93854 158720 93860 158772
rect 93912 158760 93918 158772
rect 95142 158760 95148 158772
rect 93912 158732 95148 158760
rect 93912 158720 93918 158732
rect 95142 158720 95148 158732
rect 95200 158760 95206 158772
rect 223666 158760 223672 158772
rect 95200 158732 223672 158760
rect 95200 158720 95206 158732
rect 223666 158720 223672 158732
rect 223724 158720 223730 158772
rect 210418 158652 210424 158704
rect 210476 158692 210482 158704
rect 291286 158692 291292 158704
rect 210476 158664 291292 158692
rect 210476 158652 210482 158664
rect 291286 158652 291292 158664
rect 291344 158652 291350 158704
rect 45370 157972 45376 158024
rect 45428 158012 45434 158024
rect 63494 158012 63500 158024
rect 45428 157984 63500 158012
rect 45428 157972 45434 157984
rect 63494 157972 63500 157984
rect 63552 157972 63558 158024
rect 186222 157972 186228 158024
rect 186280 158012 186286 158024
rect 208394 158012 208400 158024
rect 186280 157984 208400 158012
rect 186280 157972 186286 157984
rect 208394 157972 208400 157984
rect 208452 157972 208458 158024
rect 291286 157972 291292 158024
rect 291344 158012 291350 158024
rect 582926 158012 582932 158024
rect 291344 157984 582932 158012
rect 291344 157972 291350 157984
rect 582926 157972 582932 157984
rect 582984 157972 582990 158024
rect 209774 157428 209780 157480
rect 209832 157468 209838 157480
rect 210418 157468 210424 157480
rect 209832 157440 210424 157468
rect 209832 157428 209838 157440
rect 210418 157428 210424 157440
rect 210476 157428 210482 157480
rect 63494 157360 63500 157412
rect 63552 157400 63558 157412
rect 64598 157400 64604 157412
rect 63552 157372 64604 157400
rect 63552 157360 63558 157372
rect 64598 157360 64604 157372
rect 64656 157400 64662 157412
rect 189902 157400 189908 157412
rect 64656 157372 189908 157400
rect 64656 157360 64662 157372
rect 189902 157360 189908 157372
rect 189960 157360 189966 157412
rect 202138 157360 202144 157412
rect 202196 157400 202202 157412
rect 202782 157400 202788 157412
rect 202196 157372 202788 157400
rect 202196 157360 202202 157372
rect 202782 157360 202788 157372
rect 202840 157400 202846 157412
rect 230566 157400 230572 157412
rect 202840 157372 230572 157400
rect 202840 157360 202846 157372
rect 230566 157360 230572 157372
rect 230624 157360 230630 157412
rect 206278 156680 206284 156732
rect 206336 156720 206342 156732
rect 252462 156720 252468 156732
rect 206336 156692 252468 156720
rect 206336 156680 206342 156692
rect 252462 156680 252468 156692
rect 252520 156720 252526 156732
rect 255958 156720 255964 156732
rect 252520 156692 255964 156720
rect 252520 156680 252526 156692
rect 255958 156680 255964 156692
rect 256016 156680 256022 156732
rect 220814 156612 220820 156664
rect 220872 156652 220878 156664
rect 582650 156652 582656 156664
rect 220872 156624 582656 156652
rect 220872 156612 220878 156624
rect 582650 156612 582656 156624
rect 582708 156612 582714 156664
rect 57698 156000 57704 156052
rect 57756 156040 57762 156052
rect 162210 156040 162216 156052
rect 57756 156012 162216 156040
rect 57756 156000 57762 156012
rect 162210 156000 162216 156012
rect 162268 156000 162274 156052
rect 71774 155932 71780 155984
rect 71832 155972 71838 155984
rect 72878 155972 72884 155984
rect 71832 155944 72884 155972
rect 71832 155932 71838 155944
rect 72878 155932 72884 155944
rect 72936 155972 72942 155984
rect 197446 155972 197452 155984
rect 72936 155944 197452 155972
rect 72936 155932 72942 155944
rect 197446 155932 197452 155944
rect 197504 155932 197510 155984
rect 70578 155252 70584 155304
rect 70636 155292 70642 155304
rect 74626 155292 74632 155304
rect 70636 155264 74632 155292
rect 70636 155252 70642 155264
rect 74626 155252 74632 155264
rect 74684 155292 74690 155304
rect 183002 155292 183008 155304
rect 74684 155264 183008 155292
rect 74684 155252 74690 155264
rect 183002 155252 183008 155264
rect 183060 155252 183066 155304
rect 43990 155184 43996 155236
rect 44048 155224 44054 155236
rect 178770 155224 178776 155236
rect 44048 155196 178776 155224
rect 44048 155184 44054 155196
rect 178770 155184 178776 155196
rect 178828 155184 178834 155236
rect 212718 154504 212724 154556
rect 212776 154544 212782 154556
rect 213178 154544 213184 154556
rect 212776 154516 213184 154544
rect 212776 154504 212782 154516
rect 213178 154504 213184 154516
rect 213236 154504 213242 154556
rect 88334 153892 88340 153944
rect 88392 153932 88398 153944
rect 153930 153932 153936 153944
rect 88392 153904 153936 153932
rect 88392 153892 88398 153904
rect 153930 153892 153936 153904
rect 153988 153892 153994 153944
rect 57882 153824 57888 153876
rect 57940 153864 57946 153876
rect 187050 153864 187056 153876
rect 57940 153836 187056 153864
rect 57940 153824 57946 153836
rect 187050 153824 187056 153836
rect 187108 153824 187114 153876
rect 187142 153280 187148 153332
rect 187200 153320 187206 153332
rect 224402 153320 224408 153332
rect 187200 153292 224408 153320
rect 187200 153280 187206 153292
rect 224402 153280 224408 153292
rect 224460 153280 224466 153332
rect 212718 153212 212724 153264
rect 212776 153252 212782 153264
rect 295334 153252 295340 153264
rect 212776 153224 295340 153252
rect 212776 153212 212782 153224
rect 295334 153212 295340 153224
rect 295392 153212 295398 153264
rect 215386 153144 215392 153196
rect 215444 153184 215450 153196
rect 259454 153184 259460 153196
rect 215444 153156 259460 153184
rect 215444 153144 215450 153156
rect 259454 153144 259460 153156
rect 259512 153144 259518 153196
rect 182082 152532 182088 152584
rect 182140 152572 182146 152584
rect 216674 152572 216680 152584
rect 182140 152544 216680 152572
rect 182140 152532 182146 152544
rect 216674 152532 216680 152544
rect 216732 152532 216738 152584
rect 54846 152464 54852 152516
rect 54904 152504 54910 152516
rect 184290 152504 184296 152516
rect 54904 152476 184296 152504
rect 54904 152464 54910 152476
rect 184290 152464 184296 152476
rect 184348 152464 184354 152516
rect 184198 151784 184204 151836
rect 184256 151824 184262 151836
rect 202046 151824 202052 151836
rect 184256 151796 202052 151824
rect 184256 151784 184262 151796
rect 202046 151784 202052 151796
rect 202104 151784 202110 151836
rect 180242 150492 180248 150544
rect 180300 150532 180306 150544
rect 214006 150532 214012 150544
rect 180300 150504 214012 150532
rect 180300 150492 180306 150504
rect 214006 150492 214012 150504
rect 214064 150492 214070 150544
rect 215478 150492 215484 150544
rect 215536 150532 215542 150544
rect 215938 150532 215944 150544
rect 215536 150504 215944 150532
rect 215536 150492 215542 150504
rect 215938 150492 215944 150504
rect 215996 150532 216002 150544
rect 251174 150532 251180 150544
rect 215996 150504 251180 150532
rect 215996 150492 216002 150504
rect 251174 150492 251180 150504
rect 251232 150492 251238 150544
rect 127618 150424 127624 150476
rect 127676 150464 127682 150476
rect 220906 150464 220912 150476
rect 127676 150436 220912 150464
rect 127676 150424 127682 150436
rect 220906 150424 220912 150436
rect 220964 150424 220970 150476
rect 208486 150356 208492 150408
rect 208544 150396 208550 150408
rect 209130 150396 209136 150408
rect 208544 150368 209136 150396
rect 208544 150356 208550 150368
rect 209130 150356 209136 150368
rect 209188 150396 209194 150408
rect 281718 150396 281724 150408
rect 209188 150368 281724 150396
rect 209188 150356 209194 150368
rect 281718 150356 281724 150368
rect 281776 150356 281782 150408
rect 89622 149744 89628 149796
rect 89680 149784 89686 149796
rect 127618 149784 127624 149796
rect 89680 149756 127624 149784
rect 89680 149744 89686 149756
rect 127618 149744 127624 149756
rect 127676 149744 127682 149796
rect 67726 149676 67732 149728
rect 67784 149716 67790 149728
rect 77478 149716 77484 149728
rect 67784 149688 77484 149716
rect 67784 149676 67790 149688
rect 77478 149676 77484 149688
rect 77536 149676 77542 149728
rect 124858 149676 124864 149728
rect 124916 149716 124922 149728
rect 240134 149716 240140 149728
rect 124916 149688 240140 149716
rect 124916 149676 124922 149688
rect 240134 149676 240140 149688
rect 240192 149716 240198 149728
rect 240778 149716 240784 149728
rect 240192 149688 240784 149716
rect 240192 149676 240198 149688
rect 240778 149676 240784 149688
rect 240836 149676 240842 149728
rect 77570 149132 77576 149184
rect 77628 149172 77634 149184
rect 80790 149172 80796 149184
rect 77628 149144 80796 149172
rect 77628 149132 77634 149144
rect 80790 149132 80796 149144
rect 80848 149132 80854 149184
rect 86310 149132 86316 149184
rect 86368 149172 86374 149184
rect 88978 149172 88984 149184
rect 86368 149144 88984 149172
rect 86368 149132 86374 149144
rect 88978 149132 88984 149144
rect 89036 149132 89042 149184
rect 67542 149064 67548 149116
rect 67600 149104 67606 149116
rect 105630 149104 105636 149116
rect 67600 149076 105636 149104
rect 67600 149064 67606 149076
rect 105630 149064 105636 149076
rect 105688 149064 105694 149116
rect 212442 148996 212448 149048
rect 212500 149036 212506 149048
rect 271874 149036 271880 149048
rect 212500 149008 271880 149036
rect 212500 148996 212506 149008
rect 271874 148996 271880 149008
rect 271932 148996 271938 149048
rect 183002 148384 183008 148436
rect 183060 148424 183066 148436
rect 196066 148424 196072 148436
rect 183060 148396 196072 148424
rect 183060 148384 183066 148396
rect 196066 148384 196072 148396
rect 196124 148384 196130 148436
rect 162210 148316 162216 148368
rect 162268 148356 162274 148368
rect 211798 148356 211804 148368
rect 162268 148328 211804 148356
rect 162268 148316 162274 148328
rect 211798 148316 211804 148328
rect 211856 148316 211862 148368
rect 61930 147704 61936 147756
rect 61988 147744 61994 147756
rect 127618 147744 127624 147756
rect 61988 147716 127624 147744
rect 61988 147704 61994 147716
rect 127618 147704 127624 147716
rect 127676 147704 127682 147756
rect 76190 147636 76196 147688
rect 76248 147676 76254 147688
rect 159450 147676 159456 147688
rect 76248 147648 159456 147676
rect 76248 147636 76254 147648
rect 159450 147636 159456 147648
rect 159508 147636 159514 147688
rect 205174 147636 205180 147688
rect 205232 147676 205238 147688
rect 260098 147676 260104 147688
rect 205232 147648 260104 147676
rect 205232 147636 205238 147648
rect 260098 147636 260104 147648
rect 260156 147636 260162 147688
rect 194594 146956 194600 147008
rect 194652 146996 194658 147008
rect 195054 146996 195060 147008
rect 194652 146968 195060 146996
rect 194652 146956 194658 146968
rect 195054 146956 195060 146968
rect 195112 146956 195118 147008
rect 200206 146956 200212 147008
rect 200264 146996 200270 147008
rect 200942 146996 200948 147008
rect 200264 146968 200948 146996
rect 200264 146956 200270 146968
rect 200942 146956 200948 146968
rect 201000 146956 201006 147008
rect 223666 146956 223672 147008
rect 223724 146996 223730 147008
rect 224586 146996 224592 147008
rect 223724 146968 224592 146996
rect 223724 146956 223730 146968
rect 224586 146956 224592 146968
rect 224644 146956 224650 147008
rect 60458 146888 60464 146940
rect 60516 146928 60522 146940
rect 161014 146928 161020 146940
rect 60516 146900 161020 146928
rect 60516 146888 60522 146900
rect 161014 146888 161020 146900
rect 161072 146888 161078 146940
rect 214006 146888 214012 146940
rect 214064 146928 214070 146940
rect 225046 146928 225052 146940
rect 214064 146900 225052 146928
rect 214064 146888 214070 146900
rect 225046 146888 225052 146900
rect 225104 146888 225110 146940
rect 226518 146888 226524 146940
rect 226576 146928 226582 146940
rect 264974 146928 264980 146940
rect 226576 146900 264980 146928
rect 226576 146888 226582 146900
rect 264974 146888 264980 146900
rect 265032 146888 265038 146940
rect 165522 146344 165528 146396
rect 165580 146384 165586 146396
rect 193766 146384 193772 146396
rect 165580 146356 193772 146384
rect 165580 146344 165586 146356
rect 193766 146344 193772 146356
rect 193824 146344 193830 146396
rect 98822 146276 98828 146328
rect 98880 146316 98886 146328
rect 99282 146316 99288 146328
rect 98880 146288 99288 146316
rect 98880 146276 98886 146288
rect 99282 146276 99288 146288
rect 99340 146316 99346 146328
rect 230658 146316 230664 146328
rect 99340 146288 230664 146316
rect 99340 146276 99346 146288
rect 230658 146276 230664 146288
rect 230716 146276 230722 146328
rect 196710 146208 196716 146260
rect 196768 146248 196774 146260
rect 199194 146248 199200 146260
rect 196768 146220 199200 146248
rect 196768 146208 196774 146220
rect 199194 146208 199200 146220
rect 199252 146208 199258 146260
rect 191650 145868 191656 145920
rect 191708 145908 191714 145920
rect 193858 145908 193864 145920
rect 191708 145880 193864 145908
rect 191708 145868 191714 145880
rect 193858 145868 193864 145880
rect 193916 145868 193922 145920
rect 3326 145528 3332 145580
rect 3384 145568 3390 145580
rect 95694 145568 95700 145580
rect 3384 145540 95700 145568
rect 3384 145528 3390 145540
rect 95694 145528 95700 145540
rect 95752 145528 95758 145580
rect 180150 145528 180156 145580
rect 180208 145568 180214 145580
rect 188338 145568 188344 145580
rect 180208 145540 188344 145568
rect 180208 145528 180214 145540
rect 188338 145528 188344 145540
rect 188396 145528 188402 145580
rect 234522 145528 234528 145580
rect 234580 145568 234586 145580
rect 340138 145568 340144 145580
rect 234580 145540 340144 145568
rect 234580 145528 234586 145540
rect 340138 145528 340144 145540
rect 340196 145528 340202 145580
rect 63126 144984 63132 145036
rect 63184 145024 63190 145036
rect 63310 145024 63316 145036
rect 63184 144996 63316 145024
rect 63184 144984 63190 144996
rect 63310 144984 63316 144996
rect 63368 145024 63374 145036
rect 138750 145024 138756 145036
rect 63368 144996 138756 145024
rect 63368 144984 63374 144996
rect 138750 144984 138756 144996
rect 138808 144984 138814 145036
rect 206462 144984 206468 145036
rect 206520 145024 206526 145036
rect 235258 145024 235264 145036
rect 206520 144996 235264 145024
rect 206520 144984 206526 144996
rect 235258 144984 235264 144996
rect 235316 144984 235322 145036
rect 95418 144916 95424 144968
rect 95476 144956 95482 144968
rect 95694 144956 95700 144968
rect 95476 144928 95700 144956
rect 95476 144916 95482 144928
rect 95694 144916 95700 144928
rect 95752 144956 95758 144968
rect 226518 144956 226524 144968
rect 95752 144928 226524 144956
rect 95752 144916 95758 144928
rect 226518 144916 226524 144928
rect 226576 144916 226582 144968
rect 51810 144848 51816 144900
rect 51868 144888 51874 144900
rect 87598 144888 87604 144900
rect 51868 144860 87604 144888
rect 51868 144848 51874 144860
rect 87598 144848 87604 144860
rect 87656 144848 87662 144900
rect 97442 144848 97448 144900
rect 97500 144888 97506 144900
rect 100202 144888 100208 144900
rect 97500 144860 100208 144888
rect 97500 144848 97506 144860
rect 100202 144848 100208 144860
rect 100260 144848 100266 144900
rect 73798 144168 73804 144220
rect 73856 144208 73862 144220
rect 165522 144208 165528 144220
rect 73856 144180 165528 144208
rect 73856 144168 73862 144180
rect 165522 144168 165528 144180
rect 165580 144168 165586 144220
rect 186866 143624 186872 143676
rect 186924 143664 186930 143676
rect 225598 143664 225604 143676
rect 186924 143636 225604 143664
rect 186924 143624 186930 143636
rect 225598 143624 225604 143636
rect 225656 143624 225662 143676
rect 156598 143556 156604 143608
rect 156656 143596 156662 143608
rect 211246 143596 211252 143608
rect 156656 143568 211252 143596
rect 156656 143556 156662 143568
rect 211246 143556 211252 143568
rect 211304 143556 211310 143608
rect 220078 143556 220084 143608
rect 220136 143596 220142 143608
rect 246298 143596 246304 143608
rect 220136 143568 246304 143596
rect 220136 143556 220142 143568
rect 246298 143556 246304 143568
rect 246356 143556 246362 143608
rect 219526 143080 219532 143132
rect 219584 143120 219590 143132
rect 220722 143120 220728 143132
rect 219584 143092 220728 143120
rect 219584 143080 219590 143092
rect 220722 143080 220728 143092
rect 220780 143080 220786 143132
rect 218238 142944 218244 142996
rect 218296 142984 218302 142996
rect 218698 142984 218704 142996
rect 218296 142956 218704 142984
rect 218296 142944 218302 142956
rect 218698 142944 218704 142956
rect 218756 142944 218762 142996
rect 92566 142808 92572 142860
rect 92624 142848 92630 142860
rect 149698 142848 149704 142860
rect 92624 142820 149704 142848
rect 92624 142808 92630 142820
rect 149698 142808 149704 142820
rect 149756 142848 149762 142860
rect 221918 142848 221924 142860
rect 149756 142820 221924 142848
rect 149756 142808 149762 142820
rect 221918 142808 221924 142820
rect 221976 142808 221982 142860
rect 60550 142196 60556 142248
rect 60608 142236 60614 142248
rect 93210 142236 93216 142248
rect 60608 142208 93216 142236
rect 60608 142196 60614 142208
rect 93210 142196 93216 142208
rect 93268 142196 93274 142248
rect 223206 142196 223212 142248
rect 223264 142236 223270 142248
rect 238018 142236 238024 142248
rect 223264 142208 238024 142236
rect 223264 142196 223270 142208
rect 238018 142196 238024 142208
rect 238076 142196 238082 142248
rect 46198 142128 46204 142180
rect 46256 142168 46262 142180
rect 88702 142168 88708 142180
rect 46256 142140 88708 142168
rect 46256 142128 46262 142140
rect 88702 142128 88708 142140
rect 88760 142128 88766 142180
rect 204898 142128 204904 142180
rect 204956 142168 204962 142180
rect 209774 142168 209780 142180
rect 204956 142140 209780 142168
rect 204956 142128 204962 142140
rect 209774 142128 209780 142140
rect 209832 142128 209838 142180
rect 218238 142128 218244 142180
rect 218296 142168 218302 142180
rect 280890 142168 280896 142180
rect 218296 142140 280896 142168
rect 218296 142128 218302 142140
rect 280890 142128 280896 142140
rect 280948 142128 280954 142180
rect 63310 141516 63316 141568
rect 63368 141556 63374 141568
rect 76558 141556 76564 141568
rect 63368 141528 76564 141556
rect 63368 141516 63374 141528
rect 76558 141516 76564 141528
rect 76616 141516 76622 141568
rect 76190 141448 76196 141500
rect 76248 141488 76254 141500
rect 159358 141488 159364 141500
rect 76248 141460 159364 141488
rect 76248 141448 76254 141460
rect 159358 141448 159364 141460
rect 159416 141488 159422 141500
rect 203150 141488 203156 141500
rect 159416 141460 203156 141488
rect 159416 141448 159422 141460
rect 203150 141448 203156 141460
rect 203208 141448 203214 141500
rect 39850 141380 39856 141432
rect 39908 141420 39914 141432
rect 72326 141420 72332 141432
rect 39908 141392 72332 141420
rect 39908 141380 39914 141392
rect 72326 141380 72332 141392
rect 72384 141380 72390 141432
rect 75822 141380 75828 141432
rect 75880 141420 75886 141432
rect 170582 141420 170588 141432
rect 75880 141392 170588 141420
rect 75880 141380 75886 141392
rect 170582 141380 170588 141392
rect 170640 141420 170646 141432
rect 202598 141420 202604 141432
rect 170640 141392 202604 141420
rect 170640 141380 170646 141392
rect 202598 141380 202604 141392
rect 202656 141380 202662 141432
rect 219434 141380 219440 141432
rect 219492 141420 219498 141432
rect 258718 141420 258724 141432
rect 219492 141392 258724 141420
rect 219492 141380 219498 141392
rect 258718 141380 258724 141392
rect 258776 141380 258782 141432
rect 203426 140768 203432 140820
rect 203484 140808 203490 140820
rect 289078 140808 289084 140820
rect 203484 140780 289084 140808
rect 203484 140768 203490 140780
rect 289078 140768 289084 140780
rect 289136 140768 289142 140820
rect 214650 140604 214656 140616
rect 200086 140576 214656 140604
rect 188982 140428 188988 140480
rect 189040 140468 189046 140480
rect 194778 140468 194784 140480
rect 189040 140440 194784 140468
rect 189040 140428 189046 140440
rect 194778 140428 194784 140440
rect 194836 140428 194842 140480
rect 64782 140020 64788 140072
rect 64840 140060 64846 140072
rect 76650 140060 76656 140072
rect 64840 140032 76656 140060
rect 64840 140020 64846 140032
rect 76650 140020 76656 140032
rect 76708 140020 76714 140072
rect 85942 140020 85948 140072
rect 86000 140060 86006 140072
rect 174630 140060 174636 140072
rect 86000 140032 174636 140060
rect 86000 140020 86006 140032
rect 174630 140020 174636 140032
rect 174688 140020 174694 140072
rect 59078 139408 59084 139460
rect 59136 139448 59142 139460
rect 104250 139448 104256 139460
rect 59136 139420 104256 139448
rect 59136 139408 59142 139420
rect 104250 139408 104256 139420
rect 104308 139408 104314 139460
rect 174630 139408 174636 139460
rect 174688 139448 174694 139460
rect 200086 139448 200114 140576
rect 214650 140564 214656 140576
rect 214708 140564 214714 140616
rect 213730 140496 213736 140548
rect 213788 140496 213794 140548
rect 174688 139420 200114 139448
rect 174688 139408 174694 139420
rect 213748 139380 213776 140496
rect 214834 140428 214840 140480
rect 214892 140468 214898 140480
rect 214892 140440 219434 140468
rect 214892 140428 214898 140440
rect 219406 139448 219434 140440
rect 224494 140428 224500 140480
rect 224552 140468 224558 140480
rect 227898 140468 227904 140480
rect 224552 140440 227904 140468
rect 224552 140428 224558 140440
rect 227898 140428 227904 140440
rect 227956 140428 227962 140480
rect 249058 139448 249064 139460
rect 219406 139420 249064 139448
rect 249058 139408 249064 139420
rect 249116 139408 249122 139460
rect 213748 139352 219434 139380
rect 219406 138768 219434 139352
rect 316034 138768 316040 138780
rect 219406 138740 316040 138768
rect 316034 138728 316040 138740
rect 316092 138728 316098 138780
rect 51718 138660 51724 138712
rect 51776 138700 51782 138712
rect 71222 138700 71228 138712
rect 51776 138672 71228 138700
rect 51776 138660 51782 138672
rect 71222 138660 71228 138672
rect 71280 138660 71286 138712
rect 88518 138660 88524 138712
rect 88576 138700 88582 138712
rect 185578 138700 185584 138712
rect 88576 138672 185584 138700
rect 88576 138660 88582 138672
rect 185578 138660 185584 138672
rect 185636 138660 185642 138712
rect 226610 138660 226616 138712
rect 226668 138700 226674 138712
rect 230474 138700 230480 138712
rect 226668 138672 230480 138700
rect 226668 138660 226674 138672
rect 230474 138660 230480 138672
rect 230532 138700 230538 138712
rect 582558 138700 582564 138712
rect 230532 138672 582564 138700
rect 230532 138660 230538 138672
rect 582558 138660 582564 138672
rect 582616 138660 582622 138712
rect 77386 138048 77392 138100
rect 77444 138088 77450 138100
rect 77938 138088 77944 138100
rect 77444 138060 77944 138088
rect 77444 138048 77450 138060
rect 77938 138048 77944 138060
rect 77996 138048 78002 138100
rect 82906 138048 82912 138100
rect 82964 138088 82970 138100
rect 83550 138088 83556 138100
rect 82964 138060 83556 138088
rect 82964 138048 82970 138060
rect 83550 138048 83556 138060
rect 83608 138048 83614 138100
rect 89714 138048 89720 138100
rect 89772 138088 89778 138100
rect 90174 138088 90180 138100
rect 89772 138060 90180 138088
rect 89772 138048 89778 138060
rect 90174 138048 90180 138060
rect 90232 138048 90238 138100
rect 92382 138048 92388 138100
rect 92440 138088 92446 138100
rect 92566 138088 92572 138100
rect 92440 138060 92572 138088
rect 92440 138048 92446 138060
rect 92566 138048 92572 138060
rect 92624 138048 92630 138100
rect 64506 137980 64512 138032
rect 64564 138020 64570 138032
rect 81434 138020 81440 138032
rect 64564 137992 81440 138020
rect 64564 137980 64570 137992
rect 81434 137980 81440 137992
rect 81492 137980 81498 138032
rect 3234 137912 3240 137964
rect 3292 137952 3298 137964
rect 72970 137952 72976 137964
rect 3292 137924 72976 137952
rect 3292 137912 3298 137924
rect 72970 137912 72976 137924
rect 73028 137912 73034 137964
rect 190086 137776 190092 137828
rect 190144 137816 190150 137828
rect 192570 137816 192576 137828
rect 190144 137788 192576 137816
rect 190144 137776 190150 137788
rect 192570 137776 192576 137788
rect 192628 137776 192634 137828
rect 97350 137300 97356 137352
rect 97408 137340 97414 137352
rect 100846 137340 100852 137352
rect 97408 137312 100852 137340
rect 97408 137300 97414 137312
rect 100846 137300 100852 137312
rect 100904 137300 100910 137352
rect 88702 137232 88708 137284
rect 88760 137272 88766 137284
rect 96798 137272 96804 137284
rect 88760 137244 96804 137272
rect 88760 137232 88766 137244
rect 96798 137232 96804 137244
rect 96856 137232 96862 137284
rect 169202 137232 169208 137284
rect 169260 137272 169266 137284
rect 187142 137272 187148 137284
rect 169260 137244 187148 137272
rect 169260 137232 169266 137244
rect 187142 137232 187148 137244
rect 187200 137232 187206 137284
rect 226610 137232 226616 137284
rect 226668 137272 226674 137284
rect 233234 137272 233240 137284
rect 226668 137244 233240 137272
rect 226668 137232 226674 137244
rect 233234 137232 233240 137244
rect 233292 137272 233298 137284
rect 233878 137272 233884 137284
rect 233292 137244 233884 137272
rect 233292 137232 233298 137244
rect 233878 137232 233884 137244
rect 233936 137232 233942 137284
rect 72970 136688 72976 136740
rect 73028 136728 73034 136740
rect 73154 136728 73160 136740
rect 73028 136700 73160 136728
rect 73028 136688 73034 136700
rect 73154 136688 73160 136700
rect 73212 136688 73218 136740
rect 74442 136688 74448 136740
rect 74500 136728 74506 136740
rect 75178 136728 75184 136740
rect 74500 136700 75184 136728
rect 74500 136688 74506 136700
rect 75178 136688 75184 136700
rect 75236 136688 75242 136740
rect 81066 136688 81072 136740
rect 81124 136728 81130 136740
rect 83458 136728 83464 136740
rect 81124 136700 83464 136728
rect 81124 136688 81130 136700
rect 83458 136688 83464 136700
rect 83516 136688 83522 136740
rect 85206 136688 85212 136740
rect 85264 136728 85270 136740
rect 86310 136728 86316 136740
rect 85264 136700 86316 136728
rect 85264 136688 85270 136700
rect 86310 136688 86316 136700
rect 86368 136688 86374 136740
rect 66070 136620 66076 136672
rect 66128 136660 66134 136672
rect 141694 136660 141700 136672
rect 66128 136632 141700 136660
rect 66128 136620 66134 136632
rect 141694 136620 141700 136632
rect 141752 136620 141758 136672
rect 88334 136552 88340 136604
rect 88392 136592 88398 136604
rect 89622 136592 89628 136604
rect 88392 136564 89628 136592
rect 88392 136552 88398 136564
rect 89622 136552 89628 136564
rect 89680 136592 89686 136604
rect 91186 136592 91192 136604
rect 89680 136564 91192 136592
rect 89680 136552 89686 136564
rect 91186 136552 91192 136564
rect 91244 136552 91250 136604
rect 171870 136552 171876 136604
rect 171928 136592 171934 136604
rect 191650 136592 191656 136604
rect 171928 136564 191656 136592
rect 171928 136552 171934 136564
rect 191650 136552 191656 136564
rect 191708 136552 191714 136604
rect 88610 136008 88616 136060
rect 88668 136048 88674 136060
rect 89254 136048 89260 136060
rect 88668 136020 89260 136048
rect 88668 136008 88674 136020
rect 89254 136008 89260 136020
rect 89312 136008 89318 136060
rect 93762 135940 93768 135992
rect 93820 135980 93826 135992
rect 141602 135980 141608 135992
rect 93820 135952 141608 135980
rect 93820 135940 93826 135952
rect 141602 135940 141608 135952
rect 141660 135940 141666 135992
rect 3418 135872 3424 135924
rect 3476 135912 3482 135924
rect 88334 135912 88340 135924
rect 3476 135884 88340 135912
rect 3476 135872 3482 135884
rect 88334 135872 88340 135884
rect 88392 135872 88398 135924
rect 94222 135872 94228 135924
rect 94280 135912 94286 135924
rect 151262 135912 151268 135924
rect 94280 135884 151268 135912
rect 94280 135872 94286 135884
rect 151262 135872 151268 135884
rect 151320 135872 151326 135924
rect 159358 135872 159364 135924
rect 159416 135912 159422 135924
rect 169110 135912 169116 135924
rect 159416 135884 169116 135912
rect 159416 135872 159422 135884
rect 169110 135872 169116 135884
rect 169168 135872 169174 135924
rect 67266 135260 67272 135312
rect 67324 135300 67330 135312
rect 94866 135300 94872 135312
rect 67324 135272 94872 135300
rect 67324 135260 67330 135272
rect 94866 135260 94872 135272
rect 94924 135260 94930 135312
rect 180150 135260 180156 135312
rect 180208 135300 180214 135312
rect 191650 135300 191656 135312
rect 180208 135272 191656 135300
rect 180208 135260 180214 135272
rect 191650 135260 191656 135272
rect 191708 135260 191714 135312
rect 226794 135192 226800 135244
rect 226852 135232 226858 135244
rect 278774 135232 278780 135244
rect 226852 135204 278780 135232
rect 226852 135192 226858 135204
rect 278774 135192 278780 135204
rect 278832 135232 278838 135244
rect 280062 135232 280068 135244
rect 278832 135204 280068 135232
rect 278832 135192 278838 135204
rect 280062 135192 280068 135204
rect 280120 135192 280126 135244
rect 69566 134988 69572 135040
rect 69624 135028 69630 135040
rect 73798 135028 73804 135040
rect 69624 135000 73804 135028
rect 69624 134988 69630 135000
rect 73798 134988 73804 135000
rect 73856 134988 73862 135040
rect 68646 134784 68652 134836
rect 68704 134824 68710 134836
rect 69658 134824 69664 134836
rect 68704 134796 69664 134824
rect 68704 134784 68710 134796
rect 69658 134784 69664 134796
rect 69716 134784 69722 134836
rect 93210 134580 93216 134632
rect 93268 134620 93274 134632
rect 147122 134620 147128 134632
rect 93268 134592 147128 134620
rect 93268 134580 93274 134592
rect 147122 134580 147128 134592
rect 147180 134580 147186 134632
rect 94866 134512 94872 134564
rect 94924 134552 94930 134564
rect 174630 134552 174636 134564
rect 94924 134524 174636 134552
rect 94924 134512 94930 134524
rect 174630 134512 174636 134524
rect 174688 134512 174694 134564
rect 280062 134512 280068 134564
rect 280120 134552 280126 134564
rect 307018 134552 307024 134564
rect 280120 134524 307024 134552
rect 280120 134512 280126 134524
rect 307018 134512 307024 134524
rect 307076 134512 307082 134564
rect 173802 133832 173808 133884
rect 173860 133872 173866 133884
rect 192478 133872 192484 133884
rect 173860 133844 192484 133872
rect 173860 133832 173866 133844
rect 192478 133832 192484 133844
rect 192536 133832 192542 133884
rect 226610 133696 226616 133748
rect 226668 133736 226674 133748
rect 229186 133736 229192 133748
rect 226668 133708 229192 133736
rect 226668 133696 226674 133708
rect 229186 133696 229192 133708
rect 229244 133696 229250 133748
rect 96614 133152 96620 133204
rect 96672 133192 96678 133204
rect 184382 133192 184388 133204
rect 96672 133164 184388 133192
rect 96672 133152 96678 133164
rect 184382 133152 184388 133164
rect 184440 133152 184446 133204
rect 225598 133152 225604 133204
rect 225656 133192 225662 133204
rect 273438 133192 273444 133204
rect 225656 133164 273444 133192
rect 225656 133152 225662 133164
rect 273438 133152 273444 133164
rect 273496 133152 273502 133204
rect 50982 132404 50988 132456
rect 51040 132444 51046 132456
rect 66254 132444 66260 132456
rect 51040 132416 66260 132444
rect 51040 132404 51046 132416
rect 66254 132404 66260 132416
rect 66312 132404 66318 132456
rect 138750 132404 138756 132456
rect 138808 132444 138814 132456
rect 190454 132444 190460 132456
rect 138808 132416 190460 132444
rect 138808 132404 138814 132416
rect 190454 132404 190460 132416
rect 190512 132444 190518 132456
rect 191098 132444 191104 132456
rect 190512 132416 191104 132444
rect 190512 132404 190518 132416
rect 191098 132404 191104 132416
rect 191156 132404 191162 132456
rect 235258 132404 235264 132456
rect 235316 132444 235322 132456
rect 280798 132444 280804 132456
rect 235316 132416 280804 132444
rect 235316 132404 235322 132416
rect 280798 132404 280804 132416
rect 280856 132404 280862 132456
rect 64690 132336 64696 132388
rect 64748 132376 64754 132388
rect 66346 132376 66352 132388
rect 64748 132348 66352 132376
rect 64748 132336 64754 132348
rect 66346 132336 66352 132348
rect 66404 132336 66410 132388
rect 96706 132336 96712 132388
rect 96764 132376 96770 132388
rect 148410 132376 148416 132388
rect 96764 132348 148416 132376
rect 96764 132336 96770 132348
rect 148410 132336 148416 132348
rect 148468 132336 148474 132388
rect 226334 132336 226340 132388
rect 226392 132376 226398 132388
rect 238846 132376 238852 132388
rect 226392 132348 238852 132376
rect 226392 132336 226398 132348
rect 238846 132336 238852 132348
rect 238904 132336 238910 132388
rect 280798 131724 280804 131776
rect 280856 131764 280862 131776
rect 305638 131764 305644 131776
rect 280856 131736 305644 131764
rect 280856 131724 280862 131736
rect 305638 131724 305644 131736
rect 305696 131724 305702 131776
rect 57790 131044 57796 131096
rect 57848 131084 57854 131096
rect 66254 131084 66260 131096
rect 57848 131056 66260 131084
rect 57848 131044 57854 131056
rect 66254 131044 66260 131056
rect 66312 131044 66318 131096
rect 156690 131044 156696 131096
rect 156748 131084 156754 131096
rect 190822 131084 190828 131096
rect 156748 131056 190828 131084
rect 156748 131044 156754 131056
rect 190822 131044 190828 131056
rect 190880 131044 190886 131096
rect 226334 131044 226340 131096
rect 226392 131084 226398 131096
rect 266354 131084 266360 131096
rect 226392 131056 266360 131084
rect 226392 131044 226398 131056
rect 266354 131044 266360 131056
rect 266412 131044 266418 131096
rect 96614 130568 96620 130620
rect 96672 130608 96678 130620
rect 102778 130608 102784 130620
rect 96672 130580 102784 130608
rect 96672 130568 96678 130580
rect 102778 130568 102784 130580
rect 102836 130568 102842 130620
rect 107010 130432 107016 130484
rect 107068 130472 107074 130484
rect 152550 130472 152556 130484
rect 107068 130444 152556 130472
rect 107068 130432 107074 130444
rect 152550 130432 152556 130444
rect 152608 130432 152614 130484
rect 96706 130364 96712 130416
rect 96764 130404 96770 130416
rect 188430 130404 188436 130416
rect 96764 130376 188436 130404
rect 96764 130364 96770 130376
rect 188430 130364 188436 130376
rect 188488 130364 188494 130416
rect 96706 129684 96712 129736
rect 96764 129724 96770 129736
rect 181530 129724 181536 129736
rect 96764 129696 181536 129724
rect 96764 129684 96770 129696
rect 181530 129684 181536 129696
rect 181588 129684 181594 129736
rect 227070 129684 227076 129736
rect 227128 129724 227134 129736
rect 227898 129724 227904 129736
rect 227128 129696 227904 129724
rect 227128 129684 227134 129696
rect 227898 129684 227904 129696
rect 227956 129724 227962 129736
rect 276382 129724 276388 129736
rect 227956 129696 276388 129724
rect 227956 129684 227962 129696
rect 276382 129684 276388 129696
rect 276440 129724 276446 129736
rect 278038 129724 278044 129736
rect 276440 129696 278044 129724
rect 276440 129684 276446 129696
rect 278038 129684 278044 129696
rect 278096 129684 278102 129736
rect 102778 129004 102784 129056
rect 102836 129044 102842 129056
rect 156598 129044 156604 129056
rect 102836 129016 156604 129044
rect 102836 129004 102842 129016
rect 156598 129004 156604 129016
rect 156656 129004 156662 129056
rect 225322 128868 225328 128920
rect 225380 128908 225386 128920
rect 228450 128908 228456 128920
rect 225380 128880 228456 128908
rect 225380 128868 225386 128880
rect 228450 128868 228456 128880
rect 228508 128868 228514 128920
rect 61654 128664 61660 128716
rect 61712 128704 61718 128716
rect 66254 128704 66260 128716
rect 61712 128676 66260 128704
rect 61712 128664 61718 128676
rect 66254 128664 66260 128676
rect 66312 128664 66318 128716
rect 189074 128664 189080 128716
rect 189132 128704 189138 128716
rect 191650 128704 191656 128716
rect 189132 128676 191656 128704
rect 189132 128664 189138 128676
rect 191650 128664 191656 128676
rect 191708 128664 191714 128716
rect 64598 128256 64604 128308
rect 64656 128296 64662 128308
rect 66898 128296 66904 128308
rect 64656 128268 66904 128296
rect 64656 128256 64662 128268
rect 66898 128256 66904 128268
rect 66956 128256 66962 128308
rect 97626 128256 97632 128308
rect 97684 128296 97690 128308
rect 147030 128296 147036 128308
rect 97684 128268 147036 128296
rect 97684 128256 97690 128268
rect 147030 128256 147036 128268
rect 147088 128256 147094 128308
rect 226794 128256 226800 128308
rect 226852 128296 226858 128308
rect 237374 128296 237380 128308
rect 226852 128268 237380 128296
rect 226852 128256 226858 128268
rect 237374 128256 237380 128268
rect 237432 128256 237438 128308
rect 237374 127576 237380 127628
rect 237432 127616 237438 127628
rect 331858 127616 331864 127628
rect 237432 127588 331864 127616
rect 237432 127576 237438 127588
rect 331858 127576 331864 127588
rect 331916 127576 331922 127628
rect 181530 126964 181536 127016
rect 181588 127004 181594 127016
rect 191650 127004 191656 127016
rect 181588 126976 191656 127004
rect 181588 126964 181594 126976
rect 191650 126964 191656 126976
rect 191708 126964 191714 127016
rect 54938 126896 54944 126948
rect 54996 126936 55002 126948
rect 66898 126936 66904 126948
rect 54996 126908 66904 126936
rect 54996 126896 55002 126908
rect 66898 126896 66904 126908
rect 66956 126896 66962 126948
rect 97902 126896 97908 126948
rect 97960 126936 97966 126948
rect 152642 126936 152648 126948
rect 97960 126908 152648 126936
rect 97960 126896 97966 126908
rect 152642 126896 152648 126908
rect 152700 126896 152706 126948
rect 226610 126896 226616 126948
rect 226668 126936 226674 126948
rect 229094 126936 229100 126948
rect 226668 126908 229100 126936
rect 226668 126896 226674 126908
rect 229094 126896 229100 126908
rect 229152 126936 229158 126948
rect 281626 126936 281632 126948
rect 229152 126908 281632 126936
rect 229152 126896 229158 126908
rect 281626 126896 281632 126908
rect 281684 126896 281690 126948
rect 61838 126828 61844 126880
rect 61896 126868 61902 126880
rect 66806 126868 66812 126880
rect 61896 126840 66812 126868
rect 61896 126828 61902 126840
rect 66806 126828 66812 126840
rect 66864 126828 66870 126880
rect 226518 126828 226524 126880
rect 226576 126868 226582 126880
rect 241698 126868 241704 126880
rect 226576 126840 241704 126868
rect 226576 126828 226582 126840
rect 241698 126828 241704 126840
rect 241756 126868 241762 126880
rect 287330 126868 287336 126880
rect 241756 126840 287336 126868
rect 241756 126828 241762 126840
rect 287330 126828 287336 126840
rect 287388 126868 287394 126880
rect 288342 126868 288348 126880
rect 287388 126840 288348 126868
rect 287388 126828 287394 126840
rect 288342 126828 288348 126840
rect 288400 126828 288406 126880
rect 176010 126216 176016 126268
rect 176068 126256 176074 126268
rect 185578 126256 185584 126268
rect 176068 126228 185584 126256
rect 176068 126216 176074 126228
rect 185578 126216 185584 126228
rect 185636 126216 185642 126268
rect 288342 126216 288348 126268
rect 288400 126256 288406 126268
rect 353294 126256 353300 126268
rect 288400 126228 353300 126256
rect 288400 126216 288406 126228
rect 353294 126216 353300 126228
rect 353352 126216 353358 126268
rect 190086 125780 190092 125792
rect 189092 125752 190092 125780
rect 97810 125536 97816 125588
rect 97868 125576 97874 125588
rect 180242 125576 180248 125588
rect 97868 125548 180248 125576
rect 97868 125536 97874 125548
rect 180242 125536 180248 125548
rect 180300 125536 180306 125588
rect 189092 125576 189120 125752
rect 190086 125740 190092 125752
rect 190144 125780 190150 125792
rect 191006 125780 191012 125792
rect 190144 125752 191012 125780
rect 190144 125740 190150 125752
rect 191006 125740 191012 125752
rect 191064 125740 191070 125792
rect 190086 125604 190092 125656
rect 190144 125644 190150 125656
rect 193122 125644 193128 125656
rect 190144 125616 193128 125644
rect 190144 125604 190150 125616
rect 193122 125604 193128 125616
rect 193180 125604 193186 125656
rect 180766 125548 189120 125576
rect 97902 125468 97908 125520
rect 97960 125508 97966 125520
rect 144178 125508 144184 125520
rect 97960 125480 144184 125508
rect 97960 125468 97966 125480
rect 144178 125468 144184 125480
rect 144236 125468 144242 125520
rect 147122 125468 147128 125520
rect 147180 125508 147186 125520
rect 180766 125508 180794 125548
rect 226794 125536 226800 125588
rect 226852 125576 226858 125588
rect 231946 125576 231952 125588
rect 226852 125548 231952 125576
rect 226852 125536 226858 125548
rect 231946 125536 231952 125548
rect 232004 125576 232010 125588
rect 276198 125576 276204 125588
rect 232004 125548 276204 125576
rect 232004 125536 232010 125548
rect 276198 125536 276204 125548
rect 276256 125536 276262 125588
rect 147180 125480 180794 125508
rect 147180 125468 147186 125480
rect 63218 125332 63224 125384
rect 63276 125372 63282 125384
rect 66806 125372 66812 125384
rect 63276 125344 66812 125372
rect 63276 125332 63282 125344
rect 66806 125332 66812 125344
rect 66864 125332 66870 125384
rect 53466 124856 53472 124908
rect 53524 124896 53530 124908
rect 66806 124896 66812 124908
rect 53524 124868 66812 124896
rect 53524 124856 53530 124868
rect 66806 124856 66812 124868
rect 66864 124856 66870 124908
rect 246482 124856 246488 124908
rect 246540 124896 246546 124908
rect 298094 124896 298100 124908
rect 246540 124868 298100 124896
rect 246540 124856 246546 124868
rect 298094 124856 298100 124868
rect 298152 124856 298158 124908
rect 97902 124108 97908 124160
rect 97960 124148 97966 124160
rect 169202 124148 169208 124160
rect 97960 124120 169208 124148
rect 97960 124108 97966 124120
rect 169202 124108 169208 124120
rect 169260 124108 169266 124160
rect 226610 124108 226616 124160
rect 226668 124148 226674 124160
rect 231854 124148 231860 124160
rect 226668 124120 231860 124148
rect 226668 124108 226674 124120
rect 231854 124108 231860 124120
rect 231912 124148 231918 124160
rect 280154 124148 280160 124160
rect 231912 124120 280160 124148
rect 231912 124108 231918 124120
rect 280154 124108 280160 124120
rect 280212 124148 280218 124160
rect 582834 124148 582840 124160
rect 280212 124120 582840 124148
rect 280212 124108 280218 124120
rect 582834 124108 582840 124120
rect 582892 124108 582898 124160
rect 110966 123428 110972 123480
rect 111024 123468 111030 123480
rect 126330 123468 126336 123480
rect 111024 123440 126336 123468
rect 111024 123428 111030 123440
rect 126330 123428 126336 123440
rect 126388 123428 126394 123480
rect 141694 123428 141700 123480
rect 141752 123468 141758 123480
rect 180610 123468 180616 123480
rect 141752 123440 180616 123468
rect 141752 123428 141758 123440
rect 180610 123428 180616 123440
rect 180668 123468 180674 123480
rect 189074 123468 189080 123480
rect 180668 123440 189080 123468
rect 180668 123428 180674 123440
rect 189074 123428 189080 123440
rect 189132 123428 189138 123480
rect 182358 122816 182364 122868
rect 182416 122856 182422 122868
rect 193030 122856 193036 122868
rect 182416 122828 193036 122856
rect 182416 122816 182422 122828
rect 193030 122816 193036 122828
rect 193088 122816 193094 122868
rect 57698 122748 57704 122800
rect 57756 122788 57762 122800
rect 66346 122788 66352 122800
rect 57756 122760 66352 122788
rect 57756 122748 57762 122760
rect 66346 122748 66352 122760
rect 66404 122748 66410 122800
rect 97902 122748 97908 122800
rect 97960 122788 97966 122800
rect 129090 122788 129096 122800
rect 97960 122760 129096 122788
rect 97960 122748 97966 122760
rect 129090 122748 129096 122760
rect 129148 122748 129154 122800
rect 162302 122748 162308 122800
rect 162360 122788 162366 122800
rect 181530 122788 181536 122800
rect 162360 122760 181536 122788
rect 162360 122748 162366 122760
rect 181530 122748 181536 122760
rect 181588 122748 181594 122800
rect 226610 122748 226616 122800
rect 226668 122788 226674 122800
rect 237650 122788 237656 122800
rect 226668 122760 237656 122788
rect 226668 122748 226674 122760
rect 237650 122748 237656 122760
rect 237708 122748 237714 122800
rect 97442 122680 97448 122732
rect 97500 122720 97506 122732
rect 124950 122720 124956 122732
rect 97500 122692 124956 122720
rect 97500 122680 97506 122692
rect 124950 122680 124956 122692
rect 125008 122680 125014 122732
rect 238110 122136 238116 122188
rect 238168 122176 238174 122188
rect 246390 122176 246396 122188
rect 238168 122148 246396 122176
rect 238168 122136 238174 122148
rect 246390 122136 246396 122148
rect 246448 122136 246454 122188
rect 228450 122068 228456 122120
rect 228508 122108 228514 122120
rect 267918 122108 267924 122120
rect 228508 122080 267924 122108
rect 228508 122068 228514 122080
rect 267918 122068 267924 122080
rect 267976 122068 267982 122120
rect 181622 121932 181628 121984
rect 181680 121972 181686 121984
rect 187142 121972 187148 121984
rect 181680 121944 187148 121972
rect 181680 121932 181686 121944
rect 187142 121932 187148 121944
rect 187200 121932 187206 121984
rect 184290 121592 184296 121644
rect 184348 121632 184354 121644
rect 184842 121632 184848 121644
rect 184348 121604 184848 121632
rect 184348 121592 184354 121604
rect 184842 121592 184848 121604
rect 184900 121632 184906 121644
rect 191558 121632 191564 121644
rect 184900 121604 191564 121632
rect 184900 121592 184906 121604
rect 191558 121592 191564 121604
rect 191616 121592 191622 121644
rect 43990 121388 43996 121440
rect 44048 121428 44054 121440
rect 66806 121428 66812 121440
rect 44048 121400 66812 121428
rect 44048 121388 44054 121400
rect 66806 121388 66812 121400
rect 66864 121388 66870 121440
rect 97534 121388 97540 121440
rect 97592 121428 97598 121440
rect 110966 121428 110972 121440
rect 97592 121400 110972 121428
rect 97592 121388 97598 121400
rect 110966 121388 110972 121400
rect 111024 121388 111030 121440
rect 178770 121388 178776 121440
rect 178828 121428 178834 121440
rect 190086 121428 190092 121440
rect 178828 121400 190092 121428
rect 178828 121388 178834 121400
rect 190086 121388 190092 121400
rect 190144 121388 190150 121440
rect 226610 121388 226616 121440
rect 226668 121428 226674 121440
rect 237558 121428 237564 121440
rect 226668 121400 237564 121428
rect 226668 121388 226674 121400
rect 237558 121388 237564 121400
rect 237616 121388 237622 121440
rect 60550 121320 60556 121372
rect 60608 121360 60614 121372
rect 66898 121360 66904 121372
rect 60608 121332 66904 121360
rect 60608 121320 60614 121332
rect 66898 121320 66904 121332
rect 66956 121320 66962 121372
rect 97626 121048 97632 121100
rect 97684 121088 97690 121100
rect 102778 121088 102784 121100
rect 97684 121060 102784 121088
rect 97684 121048 97690 121060
rect 102778 121048 102784 121060
rect 102836 121048 102842 121100
rect 104250 120708 104256 120760
rect 104308 120748 104314 120760
rect 178034 120748 178040 120760
rect 104308 120720 178040 120748
rect 104308 120708 104314 120720
rect 178034 120708 178040 120720
rect 178092 120708 178098 120760
rect 233878 120708 233884 120760
rect 233936 120748 233942 120760
rect 282178 120748 282184 120760
rect 233936 120720 282184 120748
rect 233936 120708 233942 120720
rect 282178 120708 282184 120720
rect 282236 120708 282242 120760
rect 187694 120096 187700 120148
rect 187752 120136 187758 120148
rect 190822 120136 190828 120148
rect 187752 120108 190828 120136
rect 187752 120096 187758 120108
rect 190822 120096 190828 120108
rect 190880 120096 190886 120148
rect 60458 120028 60464 120080
rect 60516 120068 60522 120080
rect 66806 120068 66812 120080
rect 60516 120040 66812 120068
rect 60516 120028 60522 120040
rect 66806 120028 66812 120040
rect 66864 120028 66870 120080
rect 97166 120028 97172 120080
rect 97224 120068 97230 120080
rect 109678 120068 109684 120080
rect 97224 120040 109684 120068
rect 97224 120028 97230 120040
rect 109678 120028 109684 120040
rect 109736 120028 109742 120080
rect 160922 120028 160928 120080
rect 160980 120068 160986 120080
rect 160980 120040 180794 120068
rect 160980 120028 160986 120040
rect 59170 119960 59176 120012
rect 59228 120000 59234 120012
rect 66898 120000 66904 120012
rect 59228 119972 66904 120000
rect 59228 119960 59234 119972
rect 66898 119960 66904 119972
rect 66956 119960 66962 120012
rect 180766 120000 180794 120040
rect 187050 120028 187056 120080
rect 187108 120068 187114 120080
rect 191558 120068 191564 120080
rect 187108 120040 191564 120068
rect 187108 120028 187114 120040
rect 191558 120028 191564 120040
rect 191616 120028 191622 120080
rect 189718 120000 189724 120012
rect 180766 119972 189724 120000
rect 189718 119960 189724 119972
rect 189776 119960 189782 120012
rect 226610 119620 226616 119672
rect 226668 119660 226674 119672
rect 230566 119660 230572 119672
rect 226668 119632 230572 119660
rect 226668 119620 226674 119632
rect 230566 119620 230572 119632
rect 230624 119620 230630 119672
rect 229830 119348 229836 119400
rect 229888 119388 229894 119400
rect 313274 119388 313280 119400
rect 229888 119360 313280 119388
rect 229888 119348 229894 119360
rect 313274 119348 313280 119360
rect 313332 119348 313338 119400
rect 54846 118600 54852 118652
rect 54904 118640 54910 118652
rect 66806 118640 66812 118652
rect 54904 118612 66812 118640
rect 54904 118600 54910 118612
rect 66806 118600 66812 118612
rect 66864 118600 66870 118652
rect 97810 118600 97816 118652
rect 97868 118640 97874 118652
rect 155310 118640 155316 118652
rect 97868 118612 155316 118640
rect 97868 118600 97874 118612
rect 155310 118600 155316 118612
rect 155368 118600 155374 118652
rect 184842 118600 184848 118652
rect 184900 118640 184906 118652
rect 186958 118640 186964 118652
rect 184900 118612 186964 118640
rect 184900 118600 184906 118612
rect 186958 118600 186964 118612
rect 187016 118600 187022 118652
rect 56410 118532 56416 118584
rect 56468 118572 56474 118584
rect 66898 118572 66904 118584
rect 56468 118544 66904 118572
rect 56468 118532 56474 118544
rect 66898 118532 66904 118544
rect 66956 118532 66962 118584
rect 97902 118532 97908 118584
rect 97960 118572 97966 118584
rect 107010 118572 107016 118584
rect 97960 118544 107016 118572
rect 97960 118532 97966 118544
rect 107010 118532 107016 118544
rect 107068 118532 107074 118584
rect 226794 117988 226800 118040
rect 226852 118028 226858 118040
rect 235994 118028 236000 118040
rect 226852 118000 236000 118028
rect 226852 117988 226858 118000
rect 235994 117988 236000 118000
rect 236052 117988 236058 118040
rect 178034 117920 178040 117972
rect 178092 117960 178098 117972
rect 179322 117960 179328 117972
rect 178092 117932 179328 117960
rect 178092 117920 178098 117932
rect 179322 117920 179328 117932
rect 179380 117960 179386 117972
rect 190822 117960 190828 117972
rect 179380 117932 190828 117960
rect 179380 117920 179386 117932
rect 190822 117920 190828 117932
rect 190880 117920 190886 117972
rect 226610 117920 226616 117972
rect 226668 117960 226674 117972
rect 240134 117960 240140 117972
rect 226668 117932 240140 117960
rect 226668 117920 226674 117932
rect 240134 117920 240140 117932
rect 240192 117960 240198 117972
rect 240778 117960 240784 117972
rect 240192 117932 240784 117960
rect 240192 117920 240198 117932
rect 240778 117920 240784 117932
rect 240836 117920 240842 117972
rect 186314 117308 186320 117360
rect 186372 117348 186378 117360
rect 191558 117348 191564 117360
rect 186372 117320 191564 117348
rect 186372 117308 186378 117320
rect 191558 117308 191564 117320
rect 191616 117308 191622 117360
rect 63126 117240 63132 117292
rect 63184 117280 63190 117292
rect 66622 117280 66628 117292
rect 63184 117252 66628 117280
rect 63184 117240 63190 117252
rect 66622 117240 66628 117252
rect 66680 117240 66686 117292
rect 97902 117240 97908 117292
rect 97960 117280 97966 117292
rect 149790 117280 149796 117292
rect 97960 117252 149796 117280
rect 97960 117240 97966 117252
rect 149790 117240 149796 117252
rect 149848 117240 149854 117292
rect 159450 117240 159456 117292
rect 159508 117280 159514 117292
rect 187694 117280 187700 117292
rect 159508 117252 187700 117280
rect 159508 117240 159514 117252
rect 187694 117240 187700 117252
rect 187752 117240 187758 117292
rect 182910 117172 182916 117224
rect 182968 117212 182974 117224
rect 191374 117212 191380 117224
rect 182968 117184 191380 117212
rect 182968 117172 182974 117184
rect 191374 117172 191380 117184
rect 191432 117172 191438 117224
rect 226978 116628 226984 116680
rect 227036 116668 227042 116680
rect 238754 116668 238760 116680
rect 227036 116640 238760 116668
rect 227036 116628 227042 116640
rect 238754 116628 238760 116640
rect 238812 116628 238818 116680
rect 231762 116560 231768 116612
rect 231820 116600 231826 116612
rect 261018 116600 261024 116612
rect 231820 116572 261024 116600
rect 231820 116560 231826 116572
rect 261018 116560 261024 116572
rect 261076 116560 261082 116612
rect 188430 116016 188436 116068
rect 188488 116056 188494 116068
rect 191558 116056 191564 116068
rect 188488 116028 191564 116056
rect 188488 116016 188494 116028
rect 191558 116016 191564 116028
rect 191616 116016 191622 116068
rect 226610 115948 226616 116000
rect 226668 115988 226674 116000
rect 230474 115988 230480 116000
rect 226668 115960 230480 115988
rect 226668 115948 226674 115960
rect 230474 115948 230480 115960
rect 230532 115988 230538 116000
rect 231762 115988 231768 116000
rect 230532 115960 231768 115988
rect 230532 115948 230538 115960
rect 231762 115948 231768 115960
rect 231820 115948 231826 116000
rect 57882 115880 57888 115932
rect 57940 115920 57946 115932
rect 66806 115920 66812 115932
rect 57940 115892 66812 115920
rect 57940 115880 57946 115892
rect 66806 115880 66812 115892
rect 66864 115880 66870 115932
rect 97534 115880 97540 115932
rect 97592 115920 97598 115932
rect 124858 115920 124864 115932
rect 97592 115892 124864 115920
rect 97592 115880 97598 115892
rect 124858 115880 124864 115892
rect 124916 115880 124922 115932
rect 127618 115880 127624 115932
rect 127676 115920 127682 115932
rect 170122 115920 170128 115932
rect 127676 115892 170128 115920
rect 127676 115880 127682 115892
rect 170122 115880 170128 115892
rect 170180 115880 170186 115932
rect 97166 115676 97172 115728
rect 97224 115716 97230 115728
rect 100754 115716 100760 115728
rect 97224 115688 100760 115716
rect 97224 115676 97230 115688
rect 100754 115676 100760 115688
rect 100812 115676 100818 115728
rect 61930 115404 61936 115456
rect 61988 115444 61994 115456
rect 66898 115444 66904 115456
rect 61988 115416 66904 115444
rect 61988 115404 61994 115416
rect 66898 115404 66904 115416
rect 66956 115404 66962 115456
rect 187602 115404 187608 115456
rect 187660 115444 187666 115456
rect 191006 115444 191012 115456
rect 187660 115416 191012 115444
rect 187660 115404 187666 115416
rect 191006 115404 191012 115416
rect 191064 115404 191070 115456
rect 227990 115268 227996 115320
rect 228048 115308 228054 115320
rect 277394 115308 277400 115320
rect 228048 115280 277400 115308
rect 228048 115268 228054 115280
rect 277394 115268 277400 115280
rect 277452 115268 277458 115320
rect 170122 115200 170128 115252
rect 170180 115240 170186 115252
rect 171042 115240 171048 115252
rect 170180 115212 171048 115240
rect 170180 115200 170186 115212
rect 171042 115200 171048 115212
rect 171100 115240 171106 115252
rect 184842 115240 184848 115252
rect 171100 115212 184848 115240
rect 171100 115200 171106 115212
rect 184842 115200 184848 115212
rect 184900 115240 184906 115252
rect 186314 115240 186320 115252
rect 184900 115212 186320 115240
rect 184900 115200 184906 115212
rect 186314 115200 186320 115212
rect 186372 115200 186378 115252
rect 235994 115200 236000 115252
rect 236052 115240 236058 115252
rect 304258 115240 304264 115252
rect 236052 115212 304264 115240
rect 236052 115200 236058 115212
rect 304258 115200 304264 115212
rect 304316 115200 304322 115252
rect 59078 114452 59084 114504
rect 59136 114492 59142 114504
rect 66806 114492 66812 114504
rect 59136 114464 66812 114492
rect 59136 114452 59142 114464
rect 66806 114452 66812 114464
rect 66864 114452 66870 114504
rect 178862 114452 178868 114504
rect 178920 114492 178926 114504
rect 191558 114492 191564 114504
rect 178920 114464 191564 114492
rect 178920 114452 178926 114464
rect 191558 114452 191564 114464
rect 191616 114452 191622 114504
rect 184474 114112 184480 114164
rect 184532 114152 184538 114164
rect 186222 114152 186228 114164
rect 184532 114124 186228 114152
rect 184532 114112 184538 114124
rect 186222 114112 186228 114124
rect 186280 114112 186286 114164
rect 226518 113840 226524 113892
rect 226576 113880 226582 113892
rect 230658 113880 230664 113892
rect 226576 113852 230664 113880
rect 226576 113840 226582 113852
rect 230658 113840 230664 113852
rect 230716 113840 230722 113892
rect 7558 113772 7564 113824
rect 7616 113812 7622 113824
rect 63218 113812 63224 113824
rect 7616 113784 63224 113812
rect 7616 113772 7622 113784
rect 63218 113772 63224 113784
rect 63276 113812 63282 113824
rect 66898 113812 66904 113824
rect 63276 113784 66904 113812
rect 63276 113772 63282 113784
rect 66898 113772 66904 113784
rect 66956 113772 66962 113824
rect 244918 113772 244924 113824
rect 244976 113812 244982 113824
rect 254578 113812 254584 113824
rect 244976 113784 254584 113812
rect 244976 113772 244982 113784
rect 254578 113772 254584 113784
rect 254636 113772 254642 113824
rect 97534 113160 97540 113212
rect 97592 113200 97598 113212
rect 178770 113200 178776 113212
rect 97592 113172 178776 113200
rect 97592 113160 97598 113172
rect 178770 113160 178776 113172
rect 178828 113160 178834 113212
rect 186222 113160 186228 113212
rect 186280 113200 186286 113212
rect 190822 113200 190828 113212
rect 186280 113172 190828 113200
rect 186280 113160 186286 113172
rect 190822 113160 190828 113172
rect 190880 113160 190886 113212
rect 227806 113160 227812 113212
rect 227864 113200 227870 113212
rect 229830 113200 229836 113212
rect 227864 113172 229836 113200
rect 227864 113160 227870 113172
rect 229830 113160 229836 113172
rect 229888 113160 229894 113212
rect 157978 113092 157984 113144
rect 158036 113132 158042 113144
rect 191558 113132 191564 113144
rect 158036 113104 191564 113132
rect 158036 113092 158042 113104
rect 191558 113092 191564 113104
rect 191616 113092 191622 113144
rect 226610 113092 226616 113144
rect 226668 113132 226674 113144
rect 277486 113132 277492 113144
rect 226668 113104 277492 113132
rect 226668 113092 226674 113104
rect 277486 113092 277492 113104
rect 277544 113132 277550 113144
rect 278682 113132 278688 113144
rect 277544 113104 278688 113132
rect 277544 113092 277550 113104
rect 278682 113092 278688 113104
rect 278740 113092 278746 113144
rect 50798 112412 50804 112464
rect 50856 112452 50862 112464
rect 67174 112452 67180 112464
rect 50856 112424 67180 112452
rect 50856 112412 50862 112424
rect 67174 112412 67180 112424
rect 67232 112412 67238 112464
rect 278682 112412 278688 112464
rect 278740 112452 278746 112464
rect 324314 112452 324320 112464
rect 278740 112424 324320 112452
rect 278740 112412 278746 112424
rect 324314 112412 324320 112424
rect 324372 112412 324378 112464
rect 96706 111868 96712 111920
rect 96764 111908 96770 111920
rect 98730 111908 98736 111920
rect 96764 111880 98736 111908
rect 96764 111868 96770 111880
rect 98730 111868 98736 111880
rect 98788 111868 98794 111920
rect 97902 111800 97908 111852
rect 97960 111840 97966 111852
rect 184290 111840 184296 111852
rect 97960 111812 184296 111840
rect 97960 111800 97966 111812
rect 184290 111800 184296 111812
rect 184348 111800 184354 111852
rect 56502 111732 56508 111784
rect 56560 111772 56566 111784
rect 66898 111772 66904 111784
rect 56560 111744 66904 111772
rect 56560 111732 56566 111744
rect 66898 111732 66904 111744
rect 66956 111732 66962 111784
rect 96706 111732 96712 111784
rect 96764 111772 96770 111784
rect 98822 111772 98828 111784
rect 96764 111744 98828 111772
rect 96764 111732 96770 111744
rect 98822 111732 98828 111744
rect 98880 111732 98886 111784
rect 118694 111732 118700 111784
rect 118752 111772 118758 111784
rect 167730 111772 167736 111784
rect 118752 111744 167736 111772
rect 118752 111732 118758 111744
rect 167730 111732 167736 111744
rect 167788 111732 167794 111784
rect 177390 111732 177396 111784
rect 177448 111772 177454 111784
rect 191190 111772 191196 111784
rect 177448 111744 191196 111772
rect 177448 111732 177454 111744
rect 191190 111732 191196 111744
rect 191248 111732 191254 111784
rect 226702 111732 226708 111784
rect 226760 111772 226766 111784
rect 244366 111772 244372 111784
rect 226760 111744 244372 111772
rect 226760 111732 226766 111744
rect 244366 111732 244372 111744
rect 244424 111732 244430 111784
rect 98730 111120 98736 111172
rect 98788 111160 98794 111172
rect 118694 111160 118700 111172
rect 98788 111132 118700 111160
rect 98788 111120 98794 111132
rect 118694 111120 118700 111132
rect 118752 111120 118758 111172
rect 101398 111052 101404 111104
rect 101456 111092 101462 111104
rect 188430 111092 188436 111104
rect 101456 111064 188436 111092
rect 101456 111052 101462 111064
rect 188430 111052 188436 111064
rect 188488 111052 188494 111104
rect 244366 111052 244372 111104
rect 244424 111092 244430 111104
rect 291838 111092 291844 111104
rect 244424 111064 291844 111092
rect 244424 111052 244430 111064
rect 291838 111052 291844 111064
rect 291896 111052 291902 111104
rect 64506 110372 64512 110424
rect 64564 110412 64570 110424
rect 66806 110412 66812 110424
rect 64564 110384 66812 110412
rect 64564 110372 64570 110384
rect 66806 110372 66812 110384
rect 66864 110372 66870 110424
rect 97902 110372 97908 110424
rect 97960 110412 97966 110424
rect 184198 110412 184204 110424
rect 97960 110384 184204 110412
rect 97960 110372 97966 110384
rect 184198 110372 184204 110384
rect 184256 110372 184262 110424
rect 105630 110304 105636 110356
rect 105688 110344 105694 110356
rect 191006 110344 191012 110356
rect 105688 110316 191012 110344
rect 105688 110304 105694 110316
rect 191006 110304 191012 110316
rect 191064 110304 191070 110356
rect 97074 110236 97080 110288
rect 97132 110276 97138 110288
rect 100110 110276 100116 110288
rect 97132 110248 100116 110276
rect 97132 110236 97138 110248
rect 100110 110236 100116 110248
rect 100168 110236 100174 110288
rect 226978 109692 226984 109744
rect 227036 109732 227042 109744
rect 263686 109732 263692 109744
rect 227036 109704 263692 109732
rect 227036 109692 227042 109704
rect 263686 109692 263692 109704
rect 263744 109692 263750 109744
rect 65518 109012 65524 109064
rect 65576 109052 65582 109064
rect 65978 109052 65984 109064
rect 65576 109024 65984 109052
rect 65576 109012 65582 109024
rect 65978 109012 65984 109024
rect 66036 109012 66042 109064
rect 115382 108944 115388 108996
rect 115440 108984 115446 108996
rect 164142 108984 164148 108996
rect 115440 108956 164148 108984
rect 115440 108944 115446 108956
rect 164142 108944 164148 108956
rect 164200 108944 164206 108996
rect 226610 108944 226616 108996
rect 226668 108984 226674 108996
rect 229738 108984 229744 108996
rect 226668 108956 229744 108984
rect 226668 108944 226674 108956
rect 229738 108944 229744 108956
rect 229796 108944 229802 108996
rect 155310 108876 155316 108928
rect 155368 108916 155374 108928
rect 158622 108916 158628 108928
rect 155368 108888 158628 108916
rect 155368 108876 155374 108888
rect 158622 108876 158628 108888
rect 158680 108916 158686 108928
rect 190270 108916 190276 108928
rect 158680 108888 190276 108916
rect 158680 108876 158686 108888
rect 190270 108876 190276 108888
rect 190328 108876 190334 108928
rect 164142 108264 164148 108316
rect 164200 108304 164206 108316
rect 177390 108304 177396 108316
rect 164200 108276 177396 108304
rect 164200 108264 164206 108276
rect 177390 108264 177396 108276
rect 177448 108264 177454 108316
rect 236730 108264 236736 108316
rect 236788 108304 236794 108316
rect 259546 108304 259552 108316
rect 236788 108276 259552 108304
rect 236788 108264 236794 108276
rect 259546 108264 259552 108276
rect 259604 108264 259610 108316
rect 240042 108128 240048 108180
rect 240100 108168 240106 108180
rect 241514 108168 241520 108180
rect 240100 108140 241520 108168
rect 240100 108128 240106 108140
rect 241514 108128 241520 108140
rect 241572 108128 241578 108180
rect 97994 108060 98000 108112
rect 98052 108100 98058 108112
rect 98914 108100 98920 108112
rect 98052 108072 98920 108100
rect 98052 108060 98058 108072
rect 98914 108060 98920 108072
rect 98972 108060 98978 108112
rect 98914 107652 98920 107704
rect 98972 107692 98978 107704
rect 152550 107692 152556 107704
rect 98972 107664 152556 107692
rect 98972 107652 98978 107664
rect 152550 107652 152556 107664
rect 152608 107652 152614 107704
rect 166902 107584 166908 107636
rect 166960 107624 166966 107636
rect 190638 107624 190644 107636
rect 166960 107596 190644 107624
rect 166960 107584 166966 107596
rect 190638 107584 190644 107596
rect 190696 107584 190702 107636
rect 226702 107584 226708 107636
rect 226760 107624 226766 107636
rect 288526 107624 288532 107636
rect 226760 107596 288532 107624
rect 226760 107584 226766 107596
rect 288526 107584 288532 107596
rect 288584 107624 288590 107636
rect 289722 107624 289728 107636
rect 288584 107596 289728 107624
rect 288584 107584 288590 107596
rect 289722 107584 289728 107596
rect 289780 107584 289786 107636
rect 100110 106904 100116 106956
rect 100168 106944 100174 106956
rect 110506 106944 110512 106956
rect 100168 106916 110512 106944
rect 100168 106904 100174 106916
rect 110506 106904 110512 106916
rect 110564 106904 110570 106956
rect 289722 106904 289728 106956
rect 289780 106944 289786 106956
rect 342898 106944 342904 106956
rect 289780 106916 342904 106944
rect 289780 106904 289786 106916
rect 342898 106904 342904 106916
rect 342956 106904 342962 106956
rect 97902 106360 97908 106412
rect 97960 106400 97966 106412
rect 157978 106400 157984 106412
rect 97960 106372 157984 106400
rect 97960 106360 97966 106372
rect 157978 106360 157984 106372
rect 158036 106360 158042 106412
rect 7558 106292 7564 106344
rect 7616 106332 7622 106344
rect 66806 106332 66812 106344
rect 7616 106304 66812 106332
rect 7616 106292 7622 106304
rect 66806 106292 66812 106304
rect 66864 106292 66870 106344
rect 123570 106292 123576 106344
rect 123628 106332 123634 106344
rect 185762 106332 185768 106344
rect 123628 106304 185768 106332
rect 123628 106292 123634 106304
rect 185762 106292 185768 106304
rect 185820 106292 185826 106344
rect 96798 106224 96804 106276
rect 96856 106264 96862 106276
rect 100018 106264 100024 106276
rect 96856 106236 100024 106264
rect 96856 106224 96862 106236
rect 100018 106224 100024 106236
rect 100076 106224 100082 106276
rect 174630 106224 174636 106276
rect 174688 106264 174694 106276
rect 191006 106264 191012 106276
rect 174688 106236 191012 106264
rect 174688 106224 174694 106236
rect 191006 106224 191012 106236
rect 191064 106224 191070 106276
rect 46842 105544 46848 105596
rect 46900 105584 46906 105596
rect 66070 105584 66076 105596
rect 46900 105556 66076 105584
rect 46900 105544 46906 105556
rect 66070 105544 66076 105556
rect 66128 105584 66134 105596
rect 66622 105584 66628 105596
rect 66128 105556 66628 105584
rect 66128 105544 66134 105556
rect 66622 105544 66628 105556
rect 66680 105544 66686 105596
rect 97994 105544 98000 105596
rect 98052 105584 98058 105596
rect 123570 105584 123576 105596
rect 98052 105556 123576 105584
rect 98052 105544 98058 105556
rect 123570 105544 123576 105556
rect 123628 105544 123634 105596
rect 271782 105544 271788 105596
rect 271840 105584 271846 105596
rect 291470 105584 291476 105596
rect 271840 105556 291476 105584
rect 271840 105544 271846 105556
rect 291470 105544 291476 105556
rect 291528 105544 291534 105596
rect 188890 104864 188896 104916
rect 188948 104904 188954 104916
rect 191558 104904 191564 104916
rect 188948 104876 191564 104904
rect 188948 104864 188954 104876
rect 191558 104864 191564 104876
rect 191616 104864 191622 104916
rect 226702 104864 226708 104916
rect 226760 104904 226766 104916
rect 271782 104904 271788 104916
rect 226760 104876 271788 104904
rect 226760 104864 226766 104876
rect 271782 104864 271788 104876
rect 271840 104864 271846 104916
rect 53650 104796 53656 104848
rect 53708 104836 53714 104848
rect 66806 104836 66812 104848
rect 53708 104808 66812 104836
rect 53708 104796 53714 104808
rect 66806 104796 66812 104808
rect 66864 104796 66870 104848
rect 227438 104116 227444 104168
rect 227496 104156 227502 104168
rect 267826 104156 267832 104168
rect 227496 104128 267832 104156
rect 227496 104116 227502 104128
rect 267826 104116 267832 104128
rect 267884 104116 267890 104168
rect 102042 103504 102048 103556
rect 102100 103544 102106 103556
rect 174630 103544 174636 103556
rect 102100 103516 174636 103544
rect 102100 103504 102106 103516
rect 174630 103504 174636 103516
rect 174688 103504 174694 103556
rect 187050 103504 187056 103556
rect 187108 103544 187114 103556
rect 193214 103544 193220 103556
rect 187108 103516 193220 103544
rect 187108 103504 187114 103516
rect 193214 103504 193220 103516
rect 193272 103504 193278 103556
rect 226518 103504 226524 103556
rect 226576 103544 226582 103556
rect 231854 103544 231860 103556
rect 226576 103516 231860 103544
rect 226576 103504 226582 103516
rect 231854 103504 231860 103516
rect 231912 103544 231918 103556
rect 323578 103544 323584 103556
rect 231912 103516 323584 103544
rect 231912 103504 231918 103516
rect 323578 103504 323584 103516
rect 323636 103504 323642 103556
rect 63402 103436 63408 103488
rect 63460 103476 63466 103488
rect 67818 103476 67824 103488
rect 63460 103448 67824 103476
rect 63460 103436 63466 103448
rect 67818 103436 67824 103448
rect 67876 103436 67882 103488
rect 97902 103436 97908 103488
rect 97960 103476 97966 103488
rect 129734 103476 129740 103488
rect 97960 103448 129740 103476
rect 97960 103436 97966 103448
rect 129734 103436 129740 103448
rect 129792 103436 129798 103488
rect 97810 103368 97816 103420
rect 97868 103408 97874 103420
rect 102042 103408 102048 103420
rect 97868 103380 102048 103408
rect 97868 103368 97874 103380
rect 102042 103368 102048 103380
rect 102100 103368 102106 103420
rect 55030 102756 55036 102808
rect 55088 102796 55094 102808
rect 61746 102796 61752 102808
rect 55088 102768 61752 102796
rect 55088 102756 55094 102768
rect 61746 102756 61752 102768
rect 61804 102796 61810 102808
rect 66806 102796 66812 102808
rect 61804 102768 66812 102796
rect 61804 102756 61810 102768
rect 66806 102756 66812 102768
rect 66864 102756 66870 102808
rect 129734 102756 129740 102808
rect 129792 102796 129798 102808
rect 187234 102796 187240 102808
rect 129792 102768 187240 102796
rect 129792 102756 129798 102768
rect 187234 102756 187240 102768
rect 187292 102756 187298 102808
rect 227898 102756 227904 102808
rect 227956 102796 227962 102808
rect 258810 102796 258816 102808
rect 227956 102768 258816 102796
rect 227956 102756 227962 102768
rect 258810 102756 258816 102768
rect 258868 102756 258874 102808
rect 278038 102756 278044 102808
rect 278096 102796 278102 102808
rect 299474 102796 299480 102808
rect 278096 102768 299480 102796
rect 278096 102756 278102 102768
rect 299474 102756 299480 102768
rect 299532 102756 299538 102808
rect 188982 102212 188988 102264
rect 189040 102252 189046 102264
rect 191466 102252 191472 102264
rect 189040 102224 191472 102252
rect 189040 102212 189046 102224
rect 191466 102212 191472 102224
rect 191524 102212 191530 102264
rect 188522 102144 188528 102196
rect 188580 102184 188586 102196
rect 191558 102184 191564 102196
rect 188580 102156 191564 102184
rect 188580 102144 188586 102156
rect 191558 102144 191564 102156
rect 191616 102144 191622 102196
rect 226610 102144 226616 102196
rect 226668 102184 226674 102196
rect 226668 102156 229094 102184
rect 226668 102144 226674 102156
rect 96706 102076 96712 102128
rect 96764 102116 96770 102128
rect 98914 102116 98920 102128
rect 96764 102088 98920 102116
rect 96764 102076 96770 102088
rect 98914 102076 98920 102088
rect 98972 102076 98978 102128
rect 106274 102076 106280 102128
rect 106332 102116 106338 102128
rect 169662 102116 169668 102128
rect 106332 102088 169668 102116
rect 106332 102076 106338 102088
rect 169662 102076 169668 102088
rect 169720 102076 169726 102128
rect 229066 102116 229094 102156
rect 229738 102116 229744 102128
rect 229066 102088 229744 102116
rect 229738 102076 229744 102088
rect 229796 102116 229802 102128
rect 287054 102116 287060 102128
rect 229796 102088 287060 102116
rect 229796 102076 229802 102088
rect 287054 102076 287060 102088
rect 287112 102116 287118 102128
rect 288342 102116 288348 102128
rect 287112 102088 288348 102116
rect 287112 102076 287118 102088
rect 288342 102076 288348 102088
rect 288400 102076 288406 102128
rect 96706 101804 96712 101856
rect 96764 101844 96770 101856
rect 99374 101844 99380 101856
rect 96764 101816 99380 101844
rect 96764 101804 96770 101816
rect 99374 101804 99380 101816
rect 99432 101804 99438 101856
rect 41230 101396 41236 101448
rect 41288 101436 41294 101448
rect 65978 101436 65984 101448
rect 41288 101408 65984 101436
rect 41288 101396 41294 101408
rect 65978 101396 65984 101408
rect 66036 101436 66042 101448
rect 66530 101436 66536 101448
rect 66036 101408 66536 101436
rect 66036 101396 66042 101408
rect 66530 101396 66536 101408
rect 66588 101396 66594 101448
rect 101490 101396 101496 101448
rect 101548 101436 101554 101448
rect 106274 101436 106280 101448
rect 101548 101408 106280 101436
rect 101548 101396 101554 101408
rect 106274 101396 106280 101408
rect 106332 101396 106338 101448
rect 169662 101396 169668 101448
rect 169720 101436 169726 101448
rect 182910 101436 182916 101448
rect 169720 101408 182916 101436
rect 169720 101396 169726 101408
rect 182910 101396 182916 101408
rect 182968 101396 182974 101448
rect 288342 101396 288348 101448
rect 288400 101436 288406 101448
rect 321646 101436 321652 101448
rect 288400 101408 321652 101436
rect 288400 101396 288406 101408
rect 321646 101396 321652 101408
rect 321704 101396 321710 101448
rect 61838 100716 61844 100768
rect 61896 100756 61902 100768
rect 66806 100756 66812 100768
rect 61896 100728 66812 100756
rect 61896 100716 61902 100728
rect 66806 100716 66812 100728
rect 66864 100716 66870 100768
rect 98822 100716 98828 100768
rect 98880 100756 98886 100768
rect 190638 100756 190644 100768
rect 98880 100728 190644 100756
rect 98880 100716 98886 100728
rect 190638 100716 190644 100728
rect 190696 100716 190702 100768
rect 188338 100648 188344 100700
rect 188396 100688 188402 100700
rect 191742 100688 191748 100700
rect 188396 100660 191748 100688
rect 188396 100648 188402 100660
rect 191742 100648 191748 100660
rect 191800 100648 191806 100700
rect 230382 99968 230388 100020
rect 230440 100008 230446 100020
rect 240042 100008 240048 100020
rect 230440 99980 240048 100008
rect 230440 99968 230446 99980
rect 240042 99968 240048 99980
rect 240100 100008 240106 100020
rect 320818 100008 320824 100020
rect 240100 99980 320824 100008
rect 240100 99968 240106 99980
rect 320818 99968 320824 99980
rect 320876 99968 320882 100020
rect 185670 99560 185676 99612
rect 185728 99600 185734 99612
rect 191558 99600 191564 99612
rect 185728 99572 191564 99600
rect 185728 99560 185734 99572
rect 191558 99560 191564 99572
rect 191616 99560 191622 99612
rect 55858 99424 55864 99476
rect 55916 99464 55922 99476
rect 64598 99464 64604 99476
rect 55916 99436 64604 99464
rect 55916 99424 55922 99436
rect 64598 99424 64604 99436
rect 64656 99464 64662 99476
rect 66714 99464 66720 99476
rect 64656 99436 66720 99464
rect 64656 99424 64662 99436
rect 66714 99424 66720 99436
rect 66772 99424 66778 99476
rect 225138 99424 225144 99476
rect 225196 99464 225202 99476
rect 242802 99464 242808 99476
rect 225196 99436 242808 99464
rect 225196 99424 225202 99436
rect 242802 99424 242808 99436
rect 242860 99424 242866 99476
rect 97902 99356 97908 99408
rect 97960 99396 97966 99408
rect 185854 99396 185860 99408
rect 97960 99368 185860 99396
rect 97960 99356 97966 99368
rect 185854 99356 185860 99368
rect 185912 99356 185918 99408
rect 226426 99356 226432 99408
rect 226484 99396 226490 99408
rect 229094 99396 229100 99408
rect 226484 99368 229100 99396
rect 226484 99356 226490 99368
rect 229094 99356 229100 99368
rect 229152 99396 229158 99408
rect 230382 99396 230388 99408
rect 229152 99368 230388 99396
rect 229152 99356 229158 99368
rect 230382 99356 230388 99368
rect 230440 99356 230446 99408
rect 97902 99016 97908 99068
rect 97960 99056 97966 99068
rect 100754 99056 100760 99068
rect 97960 99028 100760 99056
rect 97960 99016 97966 99028
rect 100754 99016 100760 99028
rect 100812 99016 100818 99068
rect 97902 98132 97908 98184
rect 97960 98172 97966 98184
rect 188430 98172 188436 98184
rect 97960 98144 188436 98172
rect 97960 98132 97966 98144
rect 188430 98132 188436 98144
rect 188488 98132 188494 98184
rect 101582 98064 101588 98116
rect 101640 98104 101646 98116
rect 171042 98104 171048 98116
rect 101640 98076 171048 98104
rect 101640 98064 101646 98076
rect 171042 98064 171048 98076
rect 171100 98064 171106 98116
rect 187694 97996 187700 98048
rect 187752 98036 187758 98048
rect 191742 98036 191748 98048
rect 187752 98008 191748 98036
rect 187752 97996 187758 98008
rect 191742 97996 191748 98008
rect 191800 97996 191806 98048
rect 226702 97996 226708 98048
rect 226760 98036 226766 98048
rect 250530 98036 250536 98048
rect 226760 98008 250536 98036
rect 226760 97996 226766 98008
rect 250530 97996 250536 98008
rect 250588 98036 250594 98048
rect 250588 98008 250760 98036
rect 250588 97996 250594 98008
rect 3418 97928 3424 97980
rect 3476 97968 3482 97980
rect 46198 97968 46204 97980
rect 3476 97940 46204 97968
rect 3476 97928 3482 97940
rect 46198 97928 46204 97940
rect 46256 97928 46262 97980
rect 187142 97928 187148 97980
rect 187200 97968 187206 97980
rect 190638 97968 190644 97980
rect 187200 97940 190644 97968
rect 187200 97928 187206 97940
rect 190638 97928 190644 97940
rect 190696 97928 190702 97980
rect 250732 97968 250760 98008
rect 253198 97968 253204 97980
rect 250732 97940 253204 97968
rect 253198 97928 253204 97940
rect 253256 97928 253262 97980
rect 100018 97248 100024 97300
rect 100076 97288 100082 97300
rect 187694 97288 187700 97300
rect 100076 97260 187700 97288
rect 100076 97248 100082 97260
rect 187694 97248 187700 97260
rect 187752 97248 187758 97300
rect 96706 96840 96712 96892
rect 96764 96880 96770 96892
rect 98638 96880 98644 96892
rect 96764 96852 98644 96880
rect 96764 96840 96770 96852
rect 98638 96840 98644 96852
rect 98696 96840 98702 96892
rect 226334 96568 226340 96620
rect 226392 96608 226398 96620
rect 240870 96608 240876 96620
rect 226392 96580 240876 96608
rect 226392 96568 226398 96580
rect 240870 96568 240876 96580
rect 240928 96568 240934 96620
rect 226886 95888 226892 95940
rect 226944 95928 226950 95940
rect 266446 95928 266452 95940
rect 226944 95900 266452 95928
rect 226944 95888 226950 95900
rect 266446 95888 266452 95900
rect 266504 95888 266510 95940
rect 97810 95276 97816 95328
rect 97868 95316 97874 95328
rect 187602 95316 187608 95328
rect 97868 95288 187608 95316
rect 97868 95276 97874 95288
rect 187602 95276 187608 95288
rect 187660 95276 187666 95328
rect 64690 95208 64696 95260
rect 64748 95248 64754 95260
rect 66898 95248 66904 95260
rect 64748 95220 66904 95248
rect 64748 95208 64754 95220
rect 66898 95208 66904 95220
rect 66956 95208 66962 95260
rect 97902 95208 97908 95260
rect 97960 95248 97966 95260
rect 190454 95248 190460 95260
rect 97960 95220 190460 95248
rect 97960 95208 97966 95220
rect 190454 95208 190460 95220
rect 190512 95208 190518 95260
rect 59262 95140 59268 95192
rect 59320 95180 59326 95192
rect 66806 95180 66812 95192
rect 59320 95152 66812 95180
rect 59320 95140 59326 95152
rect 66806 95140 66812 95152
rect 66864 95140 66870 95192
rect 94866 94460 94872 94512
rect 94924 94500 94930 94512
rect 117314 94500 117320 94512
rect 94924 94472 117320 94500
rect 94924 94460 94930 94472
rect 117314 94460 117320 94472
rect 117372 94500 117378 94512
rect 193398 94500 193404 94512
rect 117372 94472 193404 94500
rect 117372 94460 117378 94472
rect 193398 94460 193404 94472
rect 193456 94460 193462 94512
rect 242802 94460 242808 94512
rect 242860 94500 242866 94512
rect 277394 94500 277400 94512
rect 242860 94472 277400 94500
rect 242860 94460 242866 94472
rect 277394 94460 277400 94472
rect 277452 94460 277458 94512
rect 97902 93644 97908 93696
rect 97960 93684 97966 93696
rect 102318 93684 102324 93696
rect 97960 93656 102324 93684
rect 97960 93644 97966 93656
rect 102318 93644 102324 93656
rect 102376 93644 102382 93696
rect 94682 93508 94688 93560
rect 94740 93548 94746 93560
rect 95878 93548 95884 93560
rect 94740 93520 95884 93548
rect 94740 93508 94746 93520
rect 95878 93508 95884 93520
rect 95936 93508 95942 93560
rect 171042 93168 171048 93220
rect 171100 93208 171106 93220
rect 191742 93208 191748 93220
rect 171100 93180 191748 93208
rect 171100 93168 171106 93180
rect 191742 93168 191748 93180
rect 191800 93208 191806 93220
rect 193766 93208 193772 93220
rect 191800 93180 193772 93208
rect 191800 93168 191806 93180
rect 193766 93168 193772 93180
rect 193824 93168 193830 93220
rect 95142 93100 95148 93152
rect 95200 93140 95206 93152
rect 120166 93140 120172 93152
rect 95200 93112 120172 93140
rect 95200 93100 95206 93112
rect 120166 93100 120172 93112
rect 120224 93140 120230 93152
rect 184382 93140 184388 93152
rect 120224 93112 184388 93140
rect 120224 93100 120230 93112
rect 184382 93100 184388 93112
rect 184440 93100 184446 93152
rect 185854 93100 185860 93152
rect 185912 93140 185918 93152
rect 205082 93140 205088 93152
rect 185912 93112 205088 93140
rect 185912 93100 185918 93112
rect 205082 93100 205088 93112
rect 205140 93100 205146 93152
rect 67542 92828 67548 92880
rect 67600 92868 67606 92880
rect 68370 92868 68376 92880
rect 67600 92840 68376 92868
rect 67600 92828 67606 92840
rect 68370 92828 68376 92840
rect 68428 92828 68434 92880
rect 95234 92800 95240 92812
rect 93826 92772 95240 92800
rect 68922 92692 68928 92744
rect 68980 92732 68986 92744
rect 70256 92732 70262 92744
rect 68980 92704 70262 92732
rect 68980 92692 68986 92704
rect 70256 92692 70262 92704
rect 70314 92692 70320 92744
rect 88656 92692 88662 92744
rect 88714 92732 88720 92744
rect 93826 92732 93854 92772
rect 95234 92760 95240 92772
rect 95292 92760 95298 92812
rect 88714 92704 93854 92732
rect 88714 92692 88720 92704
rect 81618 92556 81624 92608
rect 81676 92596 81682 92608
rect 82584 92596 82590 92608
rect 81676 92568 82590 92596
rect 81676 92556 81682 92568
rect 82584 92556 82590 92568
rect 82642 92556 82648 92608
rect 89898 92556 89904 92608
rect 89956 92596 89962 92608
rect 90680 92596 90686 92608
rect 89956 92568 90686 92596
rect 89956 92556 89962 92568
rect 90680 92556 90686 92568
rect 90738 92556 90744 92608
rect 62022 92488 62028 92540
rect 62080 92528 62086 92540
rect 67542 92528 67548 92540
rect 62080 92500 67548 92528
rect 62080 92488 62086 92500
rect 67542 92488 67548 92500
rect 67600 92488 67606 92540
rect 222838 92488 222844 92540
rect 222896 92528 222902 92540
rect 225230 92528 225236 92540
rect 222896 92500 225236 92528
rect 222896 92488 222902 92500
rect 225230 92488 225236 92500
rect 225288 92488 225294 92540
rect 52362 92420 52368 92472
rect 52420 92460 52426 92472
rect 74718 92460 74724 92472
rect 52420 92432 74724 92460
rect 52420 92420 52426 92432
rect 74718 92420 74724 92432
rect 74776 92420 74782 92472
rect 95142 92460 95148 92472
rect 85592 92432 95148 92460
rect 85592 92404 85620 92432
rect 95142 92420 95148 92432
rect 95200 92420 95206 92472
rect 190454 92420 190460 92472
rect 190512 92460 190518 92472
rect 226794 92460 226800 92472
rect 190512 92432 226800 92460
rect 190512 92420 190518 92432
rect 226794 92420 226800 92432
rect 226852 92420 226858 92472
rect 64782 92352 64788 92404
rect 64840 92392 64846 92404
rect 76282 92392 76288 92404
rect 64840 92364 76288 92392
rect 64840 92352 64846 92364
rect 76282 92352 76288 92364
rect 76340 92352 76346 92404
rect 85574 92352 85580 92404
rect 85632 92352 85638 92404
rect 88150 92352 88156 92404
rect 88208 92392 88214 92404
rect 94866 92392 94872 92404
rect 88208 92364 94872 92392
rect 88208 92352 88214 92364
rect 94866 92352 94872 92364
rect 94924 92352 94930 92404
rect 179414 92352 179420 92404
rect 179472 92392 179478 92404
rect 180702 92392 180708 92404
rect 179472 92364 180708 92392
rect 179472 92352 179478 92364
rect 180702 92352 180708 92364
rect 180760 92392 180766 92404
rect 210418 92392 210424 92404
rect 180760 92364 210424 92392
rect 180760 92352 180766 92364
rect 210418 92352 210424 92364
rect 210476 92392 210482 92404
rect 211062 92392 211068 92404
rect 210476 92364 211068 92392
rect 210476 92352 210482 92364
rect 211062 92352 211068 92364
rect 211120 92352 211126 92404
rect 95142 91060 95148 91112
rect 95200 91100 95206 91112
rect 120074 91100 120080 91112
rect 95200 91072 120080 91100
rect 95200 91060 95206 91072
rect 120074 91060 120080 91072
rect 120132 91060 120138 91112
rect 220722 91060 220728 91112
rect 220780 91100 220786 91112
rect 224954 91100 224960 91112
rect 220780 91072 224960 91100
rect 220780 91060 220786 91072
rect 224954 91060 224960 91072
rect 225012 91060 225018 91112
rect 84654 90992 84660 91044
rect 84712 91032 84718 91044
rect 100846 91032 100852 91044
rect 84712 91004 100852 91032
rect 84712 90992 84718 91004
rect 100846 90992 100852 91004
rect 100904 91032 100910 91044
rect 212166 91032 212172 91044
rect 100904 91004 212172 91032
rect 100904 90992 100910 91004
rect 212166 90992 212172 91004
rect 212224 90992 212230 91044
rect 213270 90992 213276 91044
rect 213328 91032 213334 91044
rect 228358 91032 228364 91044
rect 213328 91004 228364 91032
rect 213328 90992 213334 91004
rect 228358 90992 228364 91004
rect 228416 90992 228422 91044
rect 63310 90924 63316 90976
rect 63368 90964 63374 90976
rect 63368 90936 64874 90964
rect 63368 90924 63374 90936
rect 64846 90896 64874 90936
rect 78950 90924 78956 90976
rect 79008 90964 79014 90976
rect 110414 90964 110420 90976
rect 79008 90936 110420 90964
rect 79008 90924 79014 90936
rect 110414 90924 110420 90936
rect 110472 90924 110478 90976
rect 75730 90896 75736 90908
rect 64846 90868 75736 90896
rect 75730 90856 75736 90868
rect 75788 90856 75794 90908
rect 223758 90788 223764 90840
rect 223816 90828 223822 90840
rect 224862 90828 224868 90840
rect 223816 90800 224868 90828
rect 223816 90788 223822 90800
rect 224862 90788 224868 90800
rect 224920 90788 224926 90840
rect 222470 90244 222476 90296
rect 222528 90284 222534 90296
rect 226334 90284 226340 90296
rect 222528 90256 226340 90284
rect 222528 90244 222534 90256
rect 226334 90244 226340 90256
rect 226392 90244 226398 90296
rect 69198 89700 69204 89752
rect 69256 89740 69262 89752
rect 71038 89740 71044 89752
rect 69256 89712 71044 89740
rect 69256 89700 69262 89712
rect 71038 89700 71044 89712
rect 71096 89700 71102 89752
rect 73062 89700 73068 89752
rect 73120 89740 73126 89752
rect 74258 89740 74264 89752
rect 73120 89712 74264 89740
rect 73120 89700 73126 89712
rect 74258 89700 74264 89712
rect 74316 89700 74322 89752
rect 110414 89700 110420 89752
rect 110472 89740 110478 89752
rect 111150 89740 111156 89752
rect 110472 89712 111156 89740
rect 110472 89700 110478 89712
rect 111150 89700 111156 89712
rect 111208 89700 111214 89752
rect 111242 89700 111248 89752
rect 111300 89740 111306 89752
rect 111794 89740 111800 89752
rect 111300 89712 111800 89740
rect 111300 89700 111306 89712
rect 111794 89700 111800 89712
rect 111852 89700 111858 89752
rect 214650 89700 214656 89752
rect 214708 89740 214714 89752
rect 218790 89740 218796 89752
rect 214708 89712 218796 89740
rect 214708 89700 214714 89712
rect 218790 89700 218796 89712
rect 218848 89700 218854 89752
rect 53558 89632 53564 89684
rect 53616 89672 53622 89684
rect 73154 89672 73160 89684
rect 53616 89644 73160 89672
rect 53616 89632 53622 89644
rect 73154 89632 73160 89644
rect 73212 89672 73218 89684
rect 73706 89672 73712 89684
rect 73212 89644 73712 89672
rect 73212 89632 73218 89644
rect 73706 89632 73712 89644
rect 73764 89632 73770 89684
rect 89254 89632 89260 89684
rect 89312 89672 89318 89684
rect 111058 89672 111064 89684
rect 89312 89644 111064 89672
rect 89312 89632 89318 89644
rect 111058 89632 111064 89644
rect 111116 89672 111122 89684
rect 217686 89672 217692 89684
rect 111116 89644 217692 89672
rect 111116 89632 111122 89644
rect 217686 89632 217692 89644
rect 217744 89632 217750 89684
rect 221366 89632 221372 89684
rect 221424 89672 221430 89684
rect 236730 89672 236736 89684
rect 221424 89644 236736 89672
rect 221424 89632 221430 89644
rect 236730 89632 236736 89644
rect 236788 89632 236794 89684
rect 88702 89564 88708 89616
rect 88760 89604 88766 89616
rect 89530 89604 89536 89616
rect 88760 89576 89536 89604
rect 88760 89564 88766 89576
rect 89530 89564 89536 89576
rect 89588 89564 89594 89616
rect 114370 89564 114376 89616
rect 114428 89604 114434 89616
rect 204990 89604 204996 89616
rect 114428 89576 204996 89604
rect 114428 89564 114434 89576
rect 204990 89564 204996 89576
rect 205048 89564 205054 89616
rect 205082 89564 205088 89616
rect 205140 89604 205146 89616
rect 229094 89604 229100 89616
rect 205140 89576 229100 89604
rect 205140 89564 205146 89576
rect 229094 89564 229100 89576
rect 229152 89564 229158 89616
rect 73154 89020 73160 89072
rect 73212 89060 73218 89072
rect 77938 89060 77944 89072
rect 73212 89032 77944 89060
rect 73212 89020 73218 89032
rect 77938 89020 77944 89032
rect 77996 89020 78002 89072
rect 67450 88952 67456 89004
rect 67508 88992 67514 89004
rect 87598 88992 87604 89004
rect 67508 88964 87604 88992
rect 67508 88952 67514 88964
rect 87598 88952 87604 88964
rect 87656 88952 87662 89004
rect 194686 88544 194692 88596
rect 194744 88544 194750 88596
rect 194704 88392 194732 88544
rect 194686 88340 194692 88392
rect 194744 88340 194750 88392
rect 63218 88272 63224 88324
rect 63276 88312 63282 88324
rect 101398 88312 101404 88324
rect 63276 88284 101404 88312
rect 63276 88272 63282 88284
rect 101398 88272 101404 88284
rect 101456 88272 101462 88324
rect 120074 88272 120080 88324
rect 120132 88312 120138 88324
rect 214006 88312 214012 88324
rect 120132 88284 214012 88312
rect 120132 88272 120138 88284
rect 214006 88272 214012 88284
rect 214064 88272 214070 88324
rect 72326 88204 72332 88256
rect 72384 88244 72390 88256
rect 96982 88244 96988 88256
rect 72384 88216 96988 88244
rect 72384 88204 72390 88216
rect 96982 88204 96988 88216
rect 97040 88204 97046 88256
rect 203702 88204 203708 88256
rect 203760 88244 203766 88256
rect 204990 88244 204996 88256
rect 203760 88216 204996 88244
rect 203760 88204 203766 88216
rect 204990 88204 204996 88216
rect 205048 88204 205054 88256
rect 206278 88204 206284 88256
rect 206336 88244 206342 88256
rect 207382 88244 207388 88256
rect 206336 88216 207388 88244
rect 206336 88204 206342 88216
rect 207382 88204 207388 88216
rect 207440 88204 207446 88256
rect 226794 87592 226800 87644
rect 226852 87632 226858 87644
rect 241514 87632 241520 87644
rect 226852 87604 241520 87632
rect 226852 87592 226858 87604
rect 241514 87592 241520 87604
rect 241572 87592 241578 87644
rect 80974 86912 80980 86964
rect 81032 86952 81038 86964
rect 115382 86952 115388 86964
rect 81032 86924 115388 86952
rect 81032 86912 81038 86924
rect 115382 86912 115388 86924
rect 115440 86912 115446 86964
rect 218238 86952 218244 86964
rect 122806 86924 218244 86952
rect 89806 86844 89812 86896
rect 89864 86884 89870 86896
rect 116578 86884 116584 86896
rect 89864 86856 116584 86884
rect 89864 86844 89870 86856
rect 116578 86844 116584 86856
rect 116636 86884 116642 86896
rect 122806 86884 122834 86924
rect 218238 86912 218244 86924
rect 218296 86912 218302 86964
rect 116636 86856 122834 86884
rect 116636 86844 116642 86856
rect 185762 86844 185768 86896
rect 185820 86884 185826 86896
rect 225046 86884 225052 86896
rect 185820 86856 225052 86884
rect 185820 86844 185826 86856
rect 225046 86844 225052 86856
rect 225104 86844 225110 86896
rect 3142 85484 3148 85536
rect 3200 85524 3206 85536
rect 65518 85524 65524 85536
rect 3200 85496 65524 85524
rect 3200 85484 3206 85496
rect 65518 85484 65524 85496
rect 65576 85484 65582 85536
rect 87230 85484 87236 85536
rect 87288 85524 87294 85536
rect 121454 85524 121460 85536
rect 87288 85496 121460 85524
rect 87288 85484 87294 85496
rect 121454 85484 121460 85496
rect 121512 85524 121518 85536
rect 215294 85524 215300 85536
rect 121512 85496 215300 85524
rect 121512 85484 121518 85496
rect 215294 85484 215300 85496
rect 215352 85484 215358 85536
rect 217318 85484 217324 85536
rect 217376 85524 217382 85536
rect 244274 85524 244280 85536
rect 217376 85496 244280 85524
rect 217376 85484 217382 85496
rect 244274 85484 244280 85496
rect 244332 85484 244338 85536
rect 75454 85416 75460 85468
rect 75512 85456 75518 85468
rect 101490 85456 101496 85468
rect 75512 85428 101496 85456
rect 75512 85416 75518 85428
rect 101490 85416 101496 85428
rect 101548 85416 101554 85468
rect 193214 85416 193220 85468
rect 193272 85456 193278 85468
rect 216030 85456 216036 85468
rect 193272 85428 216036 85456
rect 193272 85416 193278 85428
rect 216030 85416 216036 85428
rect 216088 85416 216094 85468
rect 244274 84804 244280 84856
rect 244332 84844 244338 84856
rect 245562 84844 245568 84856
rect 244332 84816 245568 84844
rect 244332 84804 244338 84816
rect 245562 84804 245568 84816
rect 245620 84844 245626 84856
rect 256050 84844 256056 84856
rect 245620 84816 256056 84844
rect 245620 84804 245626 84816
rect 256050 84804 256056 84816
rect 256108 84804 256114 84856
rect 71038 84124 71044 84176
rect 71096 84164 71102 84176
rect 101582 84164 101588 84176
rect 71096 84136 101588 84164
rect 71096 84124 71102 84136
rect 101582 84124 101588 84136
rect 101640 84124 101646 84176
rect 107654 84164 107660 84176
rect 103486 84136 107660 84164
rect 80054 84056 80060 84108
rect 80112 84096 80118 84108
rect 103486 84096 103514 84136
rect 107654 84124 107660 84136
rect 107712 84164 107718 84176
rect 205634 84164 205640 84176
rect 107712 84136 205640 84164
rect 107712 84124 107718 84136
rect 205634 84124 205640 84136
rect 205692 84164 205698 84176
rect 206922 84164 206928 84176
rect 205692 84136 206928 84164
rect 205692 84124 205698 84136
rect 206922 84124 206928 84136
rect 206980 84124 206986 84176
rect 80112 84068 103514 84096
rect 80112 84056 80118 84068
rect 191650 83512 191656 83564
rect 191708 83552 191714 83564
rect 266998 83552 267004 83564
rect 191708 83524 267004 83552
rect 191708 83512 191714 83524
rect 266998 83512 267004 83524
rect 267056 83512 267062 83564
rect 210418 83444 210424 83496
rect 210476 83484 210482 83496
rect 582834 83484 582840 83496
rect 210476 83456 582840 83484
rect 210476 83444 210482 83456
rect 582834 83444 582840 83456
rect 582892 83444 582898 83496
rect 65978 82764 65984 82816
rect 66036 82804 66042 82816
rect 155494 82804 155500 82816
rect 66036 82776 155500 82804
rect 66036 82764 66042 82776
rect 155494 82764 155500 82776
rect 155552 82764 155558 82816
rect 187234 82764 187240 82816
rect 187292 82804 187298 82816
rect 229738 82804 229744 82816
rect 187292 82776 229744 82804
rect 187292 82764 187298 82776
rect 229738 82764 229744 82776
rect 229796 82764 229802 82816
rect 76006 82696 76012 82748
rect 76064 82736 76070 82748
rect 104158 82736 104164 82748
rect 76064 82708 104164 82736
rect 76064 82696 76070 82708
rect 104158 82696 104164 82708
rect 104216 82696 104222 82748
rect 200390 82084 200396 82136
rect 200448 82124 200454 82136
rect 245654 82124 245660 82136
rect 200448 82096 245660 82124
rect 200448 82084 200454 82096
rect 245654 82084 245660 82096
rect 245712 82084 245718 82136
rect 281534 82084 281540 82136
rect 281592 82124 281598 82136
rect 322934 82124 322940 82136
rect 281592 82096 322940 82124
rect 281592 82084 281598 82096
rect 322934 82084 322940 82096
rect 322992 82084 322998 82136
rect 65518 81404 65524 81456
rect 65576 81444 65582 81456
rect 65978 81444 65984 81456
rect 65576 81416 65984 81444
rect 65576 81404 65582 81416
rect 65978 81404 65984 81416
rect 66036 81404 66042 81456
rect 87598 81336 87604 81388
rect 87656 81376 87662 81388
rect 189902 81376 189908 81388
rect 87656 81348 189908 81376
rect 87656 81336 87662 81348
rect 189902 81336 189908 81348
rect 189960 81336 189966 81388
rect 80146 81268 80152 81320
rect 80204 81308 80210 81320
rect 111242 81308 111248 81320
rect 80204 81280 111248 81308
rect 80204 81268 80210 81280
rect 111242 81268 111248 81280
rect 111300 81268 111306 81320
rect 167730 81268 167736 81320
rect 167788 81308 167794 81320
rect 214558 81308 214564 81320
rect 167788 81280 214564 81308
rect 167788 81268 167794 81280
rect 214558 81268 214564 81280
rect 214616 81268 214622 81320
rect 198734 80044 198740 80096
rect 198792 80084 198798 80096
rect 244274 80084 244280 80096
rect 198792 80056 244280 80084
rect 198792 80044 198798 80056
rect 244274 80044 244280 80056
rect 244332 80044 244338 80096
rect 67726 79976 67732 80028
rect 67784 80016 67790 80028
rect 184198 80016 184204 80028
rect 67784 79988 184204 80016
rect 67784 79976 67790 79988
rect 184198 79976 184204 79988
rect 184256 80016 184262 80028
rect 184474 80016 184480 80028
rect 184256 79988 184480 80016
rect 184256 79976 184262 79988
rect 184474 79976 184480 79988
rect 184532 79976 184538 80028
rect 81710 79908 81716 79960
rect 81768 79948 81774 79960
rect 115290 79948 115296 79960
rect 81768 79920 115296 79948
rect 81768 79908 81774 79920
rect 115290 79908 115296 79920
rect 115348 79908 115354 79960
rect 177390 79908 177396 79960
rect 177448 79948 177454 79960
rect 207014 79948 207020 79960
rect 177448 79920 207020 79948
rect 177448 79908 177454 79920
rect 207014 79908 207020 79920
rect 207072 79908 207078 79960
rect 207014 79500 207020 79552
rect 207072 79540 207078 79552
rect 207658 79540 207664 79552
rect 207072 79512 207664 79540
rect 207072 79500 207078 79512
rect 207658 79500 207664 79512
rect 207716 79500 207722 79552
rect 190362 79296 190368 79348
rect 190420 79336 190426 79348
rect 284294 79336 284300 79348
rect 190420 79308 284300 79336
rect 190420 79296 190426 79308
rect 284294 79296 284300 79308
rect 284352 79296 284358 79348
rect 97442 78616 97448 78668
rect 97500 78656 97506 78668
rect 225138 78656 225144 78668
rect 97500 78628 225144 78656
rect 97500 78616 97506 78628
rect 225138 78616 225144 78628
rect 225196 78616 225202 78668
rect 97350 78548 97356 78600
rect 97408 78588 97414 78600
rect 222838 78588 222844 78600
rect 97408 78560 222844 78588
rect 97408 78548 97414 78560
rect 222838 78548 222844 78560
rect 222896 78548 222902 78600
rect 81618 77188 81624 77240
rect 81676 77228 81682 77240
rect 109034 77228 109040 77240
rect 81676 77200 109040 77228
rect 81676 77188 81682 77200
rect 109034 77188 109040 77200
rect 109092 77228 109098 77240
rect 209774 77228 209780 77240
rect 109092 77200 209780 77228
rect 109092 77188 109098 77200
rect 209774 77188 209780 77200
rect 209832 77188 209838 77240
rect 206922 77120 206928 77172
rect 206980 77160 206986 77172
rect 262858 77160 262864 77172
rect 206980 77132 262864 77160
rect 206980 77120 206986 77132
rect 262858 77120 262864 77132
rect 262916 77120 262922 77172
rect 71682 76508 71688 76560
rect 71740 76548 71746 76560
rect 171778 76548 171784 76560
rect 71740 76520 171784 76548
rect 71740 76508 71746 76520
rect 171778 76508 171784 76520
rect 171836 76508 171842 76560
rect 77938 75828 77944 75880
rect 77996 75868 78002 75880
rect 198734 75868 198740 75880
rect 77996 75840 198740 75868
rect 77996 75828 78002 75840
rect 198734 75828 198740 75840
rect 198792 75828 198798 75880
rect 227898 75868 227904 75880
rect 219406 75840 227904 75868
rect 152550 75760 152556 75812
rect 152608 75800 152614 75812
rect 219406 75800 219434 75840
rect 227898 75828 227904 75840
rect 227956 75868 227962 75880
rect 228358 75868 228364 75880
rect 227956 75840 228364 75868
rect 227956 75828 227962 75840
rect 228358 75828 228364 75840
rect 228416 75828 228422 75880
rect 152608 75772 219434 75800
rect 152608 75760 152614 75772
rect 84194 74468 84200 74520
rect 84252 74508 84258 74520
rect 115934 74508 115940 74520
rect 84252 74480 115940 74508
rect 84252 74468 84258 74480
rect 115934 74468 115940 74480
rect 115992 74508 115998 74520
rect 212534 74508 212540 74520
rect 115992 74480 212540 74508
rect 115992 74468 115998 74480
rect 212534 74468 212540 74480
rect 212592 74468 212598 74520
rect 215938 73788 215944 73840
rect 215996 73828 216002 73840
rect 248414 73828 248420 73840
rect 215996 73800 248420 73828
rect 215996 73788 216002 73800
rect 248414 73788 248420 73800
rect 248472 73788 248478 73840
rect 69842 73108 69848 73160
rect 69900 73148 69906 73160
rect 196158 73148 196164 73160
rect 69900 73120 196164 73148
rect 69900 73108 69906 73120
rect 196158 73108 196164 73120
rect 196216 73108 196222 73160
rect 212534 73108 212540 73160
rect 212592 73148 212598 73160
rect 282914 73148 282920 73160
rect 212592 73120 282920 73148
rect 212592 73108 212598 73120
rect 282914 73108 282920 73120
rect 282972 73108 282978 73160
rect 174630 73040 174636 73092
rect 174688 73080 174694 73092
rect 231854 73080 231860 73092
rect 174688 73052 231860 73080
rect 174688 73040 174694 73052
rect 231854 73040 231860 73052
rect 231912 73040 231918 73092
rect 282914 72428 282920 72480
rect 282972 72468 282978 72480
rect 333974 72468 333980 72480
rect 282972 72440 333980 72468
rect 282972 72428 282978 72440
rect 333974 72428 333980 72440
rect 334032 72428 334038 72480
rect 67818 71680 67824 71732
rect 67876 71720 67882 71732
rect 187694 71720 187700 71732
rect 67876 71692 187700 71720
rect 67876 71680 67882 71692
rect 187694 71680 187700 71692
rect 187752 71680 187758 71732
rect 196618 71680 196624 71732
rect 196676 71720 196682 71732
rect 244918 71720 244924 71732
rect 196676 71692 244924 71720
rect 196676 71680 196682 71692
rect 244918 71680 244924 71692
rect 244976 71680 244982 71732
rect 195974 71340 195980 71392
rect 196032 71380 196038 71392
rect 196618 71380 196624 71392
rect 196032 71352 196624 71380
rect 196032 71340 196038 71352
rect 196618 71340 196624 71352
rect 196676 71340 196682 71392
rect 89622 71000 89628 71052
rect 89680 71040 89686 71052
rect 163498 71040 163504 71052
rect 89680 71012 163504 71040
rect 89680 71000 89686 71012
rect 163498 71000 163504 71012
rect 163556 71000 163562 71052
rect 69198 70320 69204 70372
rect 69256 70360 69262 70372
rect 194686 70360 194692 70372
rect 69256 70332 194692 70360
rect 69256 70320 69262 70332
rect 194686 70320 194692 70332
rect 194744 70320 194750 70372
rect 194686 69912 194692 69964
rect 194744 69952 194750 69964
rect 195330 69952 195336 69964
rect 194744 69924 195336 69952
rect 194744 69912 194750 69924
rect 195330 69912 195336 69924
rect 195388 69912 195394 69964
rect 216030 69640 216036 69692
rect 216088 69680 216094 69692
rect 266354 69680 266360 69692
rect 216088 69652 266360 69680
rect 216088 69640 216094 69652
rect 266354 69640 266360 69652
rect 266412 69640 266418 69692
rect 64690 68960 64696 69012
rect 64748 69000 64754 69012
rect 192570 69000 192576 69012
rect 64748 68972 192576 69000
rect 64748 68960 64754 68972
rect 192570 68960 192576 68972
rect 192628 69000 192634 69012
rect 193030 69000 193036 69012
rect 192628 68972 193036 69000
rect 192628 68960 192634 68972
rect 193030 68960 193036 68972
rect 193088 68960 193094 69012
rect 188430 68892 188436 68944
rect 188488 68932 188494 68944
rect 250530 68932 250536 68944
rect 188488 68904 250536 68932
rect 188488 68892 188494 68904
rect 250530 68892 250536 68904
rect 250588 68892 250594 68944
rect 86862 68280 86868 68332
rect 86920 68320 86926 68332
rect 164878 68320 164884 68332
rect 86920 68292 164884 68320
rect 86920 68280 86926 68292
rect 164878 68280 164884 68292
rect 164936 68280 164942 68332
rect 193122 68280 193128 68332
rect 193180 68320 193186 68332
rect 309134 68320 309140 68332
rect 193180 68292 309140 68320
rect 193180 68280 193186 68292
rect 309134 68280 309140 68292
rect 309192 68280 309198 68332
rect 61838 67532 61844 67584
rect 61896 67572 61902 67584
rect 191098 67572 191104 67584
rect 61896 67544 191104 67572
rect 61896 67532 61902 67544
rect 191098 67532 191104 67544
rect 191156 67532 191162 67584
rect 196158 67532 196164 67584
rect 196216 67572 196222 67584
rect 285766 67572 285772 67584
rect 196216 67544 285772 67572
rect 196216 67532 196222 67544
rect 285766 67532 285772 67544
rect 285824 67532 285830 67584
rect 94498 67464 94504 67516
rect 94556 67504 94562 67516
rect 222194 67504 222200 67516
rect 94556 67476 222200 67504
rect 94556 67464 94562 67476
rect 222194 67464 222200 67476
rect 222252 67504 222258 67516
rect 222838 67504 222844 67516
rect 222252 67476 222844 67504
rect 222252 67464 222258 67476
rect 222838 67464 222844 67476
rect 222896 67464 222902 67516
rect 285766 66852 285772 66904
rect 285824 66892 285830 66904
rect 320174 66892 320180 66904
rect 285824 66864 320180 66892
rect 285824 66852 285830 66864
rect 320174 66852 320180 66864
rect 320232 66852 320238 66904
rect 86954 66172 86960 66224
rect 87012 66212 87018 66224
rect 219710 66212 219716 66224
rect 87012 66184 219716 66212
rect 87012 66172 87018 66184
rect 219710 66172 219716 66184
rect 219768 66212 219774 66224
rect 220078 66212 220084 66224
rect 219768 66184 220084 66212
rect 219768 66172 219774 66184
rect 220078 66172 220084 66184
rect 220136 66172 220142 66224
rect 66162 66104 66168 66156
rect 66220 66144 66226 66156
rect 185670 66144 185676 66156
rect 66220 66116 185676 66144
rect 66220 66104 66226 66116
rect 185670 66104 185676 66116
rect 185728 66104 185734 66156
rect 93762 64812 93768 64864
rect 93820 64852 93826 64864
rect 226334 64852 226340 64864
rect 93820 64824 226340 64852
rect 93820 64812 93826 64824
rect 226334 64812 226340 64824
rect 226392 64812 226398 64864
rect 68278 64744 68284 64796
rect 68336 64784 68342 64796
rect 193858 64784 193864 64796
rect 68336 64756 193864 64784
rect 68336 64744 68342 64756
rect 193858 64744 193864 64756
rect 193916 64744 193922 64796
rect 195330 64744 195336 64796
rect 195388 64784 195394 64796
rect 289814 64784 289820 64796
rect 195388 64756 289820 64784
rect 195388 64744 195394 64756
rect 289814 64744 289820 64756
rect 289872 64744 289878 64796
rect 289814 64132 289820 64184
rect 289872 64172 289878 64184
rect 345014 64172 345020 64184
rect 289872 64144 345020 64172
rect 289872 64132 289878 64144
rect 345014 64132 345020 64144
rect 345072 64132 345078 64184
rect 226334 63520 226340 63572
rect 226392 63560 226398 63572
rect 226978 63560 226984 63572
rect 226392 63532 226984 63560
rect 226392 63520 226398 63532
rect 226978 63520 226984 63532
rect 227036 63520 227042 63572
rect 142982 62772 142988 62824
rect 143040 62812 143046 62824
rect 180150 62812 180156 62824
rect 143040 62784 180156 62812
rect 143040 62772 143046 62784
rect 180150 62772 180156 62784
rect 180208 62772 180214 62824
rect 192478 62772 192484 62824
rect 192536 62812 192542 62824
rect 242986 62812 242992 62824
rect 192536 62784 242992 62812
rect 192536 62772 192542 62784
rect 242986 62772 242992 62784
rect 243044 62772 243050 62824
rect 89530 62024 89536 62076
rect 89588 62064 89594 62076
rect 217318 62064 217324 62076
rect 89588 62036 217324 62064
rect 89588 62024 89594 62036
rect 217318 62024 217324 62036
rect 217376 62024 217382 62076
rect 73338 60664 73344 60716
rect 73396 60704 73402 60716
rect 199378 60704 199384 60716
rect 73396 60676 199384 60704
rect 73396 60664 73402 60676
rect 199378 60664 199384 60676
rect 199436 60664 199442 60716
rect 66898 59984 66904 60036
rect 66956 60024 66962 60036
rect 131758 60024 131764 60036
rect 66956 59996 131764 60024
rect 66956 59984 66962 59996
rect 131758 59984 131764 59996
rect 131816 59984 131822 60036
rect 286410 59984 286416 60036
rect 286468 60024 286474 60036
rect 292666 60024 292672 60036
rect 286468 59996 292672 60024
rect 286468 59984 286474 59996
rect 292666 59984 292672 59996
rect 292724 59984 292730 60036
rect 2958 59304 2964 59356
rect 3016 59344 3022 59356
rect 57238 59344 57244 59356
rect 3016 59316 57244 59344
rect 3016 59304 3022 59316
rect 57238 59304 57244 59316
rect 57296 59304 57302 59356
rect 101398 59304 101404 59356
rect 101456 59344 101462 59356
rect 200114 59344 200120 59356
rect 101456 59316 200120 59344
rect 101456 59304 101462 59316
rect 200114 59304 200120 59316
rect 200172 59344 200178 59356
rect 201402 59344 201408 59356
rect 200172 59316 201408 59344
rect 200172 59304 200178 59316
rect 201402 59304 201408 59316
rect 201460 59304 201466 59356
rect 57882 58624 57888 58676
rect 57940 58664 57946 58676
rect 181438 58664 181444 58676
rect 57940 58636 181444 58664
rect 57940 58624 57946 58636
rect 181438 58624 181444 58636
rect 181496 58624 181502 58676
rect 187050 58624 187056 58676
rect 187108 58664 187114 58676
rect 269114 58664 269120 58676
rect 187108 58636 269120 58664
rect 187108 58624 187114 58636
rect 269114 58624 269120 58636
rect 269172 58624 269178 58676
rect 68922 57876 68928 57928
rect 68980 57916 68986 57928
rect 195238 57916 195244 57928
rect 68980 57888 195244 57916
rect 68980 57876 68986 57888
rect 195238 57876 195244 57888
rect 195296 57876 195302 57928
rect 111058 57808 111064 57860
rect 111116 57848 111122 57860
rect 206278 57848 206284 57860
rect 111116 57820 206284 57848
rect 111116 57808 111122 57820
rect 206278 57808 206284 57820
rect 206336 57808 206342 57860
rect 206922 57196 206928 57248
rect 206980 57236 206986 57248
rect 213178 57236 213184 57248
rect 206980 57208 213184 57236
rect 206980 57196 206986 57208
rect 213178 57196 213184 57208
rect 213236 57196 213242 57248
rect 213270 57196 213276 57248
rect 213328 57236 213334 57248
rect 280798 57236 280804 57248
rect 213328 57208 280804 57236
rect 213328 57196 213334 57208
rect 280798 57196 280804 57208
rect 280856 57196 280862 57248
rect 70394 56516 70400 56568
rect 70452 56556 70458 56568
rect 196618 56556 196624 56568
rect 70452 56528 196624 56556
rect 70452 56516 70458 56528
rect 196618 56516 196624 56528
rect 196676 56516 196682 56568
rect 201402 56516 201408 56568
rect 201460 56556 201466 56568
rect 273254 56556 273260 56568
rect 201460 56528 273260 56556
rect 201460 56516 201466 56528
rect 273254 56516 273260 56528
rect 273312 56516 273318 56568
rect 273254 55836 273260 55888
rect 273312 55876 273318 55888
rect 340966 55876 340972 55888
rect 273312 55848 340972 55876
rect 273312 55836 273318 55848
rect 340966 55836 340972 55848
rect 341024 55836 341030 55888
rect 73062 53048 73068 53100
rect 73120 53088 73126 53100
rect 138658 53088 138664 53100
rect 73120 53060 138664 53088
rect 73120 53048 73126 53060
rect 138658 53048 138664 53060
rect 138716 53048 138722 53100
rect 189718 53048 189724 53100
rect 189776 53088 189782 53100
rect 270494 53088 270500 53100
rect 189776 53060 270500 53088
rect 189776 53048 189782 53060
rect 270494 53048 270500 53060
rect 270552 53048 270558 53100
rect 101398 51688 101404 51740
rect 101456 51728 101462 51740
rect 134610 51728 134616 51740
rect 101456 51700 134616 51728
rect 101456 51688 101462 51700
rect 134610 51688 134616 51700
rect 134668 51688 134674 51740
rect 207658 51688 207664 51740
rect 207716 51728 207722 51740
rect 274634 51728 274640 51740
rect 207716 51700 274640 51728
rect 207716 51688 207722 51700
rect 274634 51688 274640 51700
rect 274692 51688 274698 51740
rect 185578 50328 185584 50380
rect 185636 50368 185642 50380
rect 248414 50368 248420 50380
rect 185636 50340 248420 50368
rect 185636 50328 185642 50340
rect 248414 50328 248420 50340
rect 248472 50328 248478 50380
rect 53650 47540 53656 47592
rect 53708 47580 53714 47592
rect 146938 47580 146944 47592
rect 53708 47552 146944 47580
rect 53708 47540 53714 47552
rect 146938 47540 146944 47552
rect 146996 47540 147002 47592
rect 183002 47540 183008 47592
rect 183060 47580 183066 47592
rect 338114 47580 338120 47592
rect 183060 47552 338120 47580
rect 183060 47540 183066 47552
rect 338114 47540 338120 47552
rect 338172 47540 338178 47592
rect 188338 46860 188344 46912
rect 188396 46900 188402 46912
rect 580166 46900 580172 46912
rect 188396 46872 580172 46900
rect 188396 46860 188402 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 115842 46248 115848 46300
rect 115900 46288 115906 46300
rect 142890 46288 142896 46300
rect 115900 46260 142896 46288
rect 115900 46248 115906 46260
rect 142890 46248 142896 46260
rect 142948 46248 142954 46300
rect 59262 46180 59268 46232
rect 59320 46220 59326 46232
rect 135898 46220 135904 46232
rect 59320 46192 135904 46220
rect 59320 46180 59326 46192
rect 135898 46180 135904 46192
rect 135956 46180 135962 46232
rect 3418 45500 3424 45552
rect 3476 45540 3482 45552
rect 65518 45540 65524 45552
rect 3476 45512 65524 45540
rect 3476 45500 3482 45512
rect 65518 45500 65524 45512
rect 65576 45500 65582 45552
rect 66162 44820 66168 44872
rect 66220 44860 66226 44872
rect 140038 44860 140044 44872
rect 66220 44832 140044 44860
rect 66220 44820 66226 44832
rect 140038 44820 140044 44832
rect 140096 44820 140102 44872
rect 184198 44820 184204 44872
rect 184256 44860 184262 44872
rect 253198 44860 253204 44872
rect 184256 44832 253204 44860
rect 184256 44820 184262 44832
rect 253198 44820 253204 44832
rect 253256 44820 253262 44872
rect 62022 43392 62028 43444
rect 62080 43432 62086 43444
rect 137370 43432 137376 43444
rect 62080 43404 137376 43432
rect 62080 43392 62086 43404
rect 137370 43392 137376 43404
rect 137428 43392 137434 43444
rect 251818 43392 251824 43444
rect 251876 43432 251882 43444
rect 349798 43432 349804 43444
rect 251876 43404 349804 43432
rect 251876 43392 251882 43404
rect 349798 43392 349804 43404
rect 349856 43392 349862 43444
rect 79962 42032 79968 42084
rect 80020 42072 80026 42084
rect 151170 42072 151176 42084
rect 80020 42044 151176 42072
rect 80020 42032 80026 42044
rect 151170 42032 151176 42044
rect 151228 42032 151234 42084
rect 199378 42032 199384 42084
rect 199436 42072 199442 42084
rect 233878 42072 233884 42084
rect 199436 42044 233884 42072
rect 199436 42032 199442 42044
rect 233878 42032 233884 42044
rect 233936 42032 233942 42084
rect 236638 42032 236644 42084
rect 236696 42072 236702 42084
rect 289814 42072 289820 42084
rect 236696 42044 289820 42072
rect 236696 42032 236702 42044
rect 289814 42032 289820 42044
rect 289872 42032 289878 42084
rect 77202 40672 77208 40724
rect 77260 40712 77266 40724
rect 142798 40712 142804 40724
rect 77260 40684 142804 40712
rect 77260 40672 77266 40684
rect 142798 40672 142804 40684
rect 142856 40672 142862 40724
rect 186958 40672 186964 40724
rect 187016 40712 187022 40724
rect 249794 40712 249800 40724
rect 187016 40684 249800 40712
rect 187016 40672 187022 40684
rect 249794 40672 249800 40684
rect 249852 40672 249858 40724
rect 250438 40672 250444 40724
rect 250496 40712 250502 40724
rect 285674 40712 285680 40724
rect 250496 40684 285680 40712
rect 250496 40672 250502 40684
rect 285674 40672 285680 40684
rect 285732 40672 285738 40724
rect 119890 39312 119896 39364
rect 119948 39352 119954 39364
rect 151078 39352 151084 39364
rect 119948 39324 151084 39352
rect 119948 39312 119954 39324
rect 151078 39312 151084 39324
rect 151136 39312 151142 39364
rect 179322 39312 179328 39364
rect 179380 39352 179386 39364
rect 305730 39352 305736 39364
rect 179380 39324 305736 39352
rect 179380 39312 179386 39324
rect 305730 39312 305736 39324
rect 305788 39312 305794 39364
rect 55030 37884 55036 37936
rect 55088 37924 55094 37936
rect 145558 37924 145564 37936
rect 55088 37896 145564 37924
rect 55088 37884 55094 37896
rect 145558 37884 145564 37896
rect 145616 37884 145622 37936
rect 180610 37884 180616 37936
rect 180668 37924 180674 37936
rect 332686 37924 332692 37936
rect 180668 37896 332692 37924
rect 180668 37884 180674 37896
rect 332686 37884 332692 37896
rect 332744 37884 332750 37936
rect 111702 36524 111708 36576
rect 111760 36564 111766 36576
rect 141510 36564 141516 36576
rect 111760 36536 141516 36564
rect 111760 36524 111766 36536
rect 141510 36524 141516 36536
rect 141568 36524 141574 36576
rect 193858 36524 193864 36576
rect 193916 36564 193922 36576
rect 291194 36564 291200 36576
rect 193916 36536 291200 36564
rect 193916 36524 193922 36536
rect 291194 36524 291200 36536
rect 291252 36524 291258 36576
rect 61654 35164 61660 35216
rect 61712 35204 61718 35216
rect 125594 35204 125600 35216
rect 61712 35176 125600 35204
rect 61712 35164 61718 35176
rect 125594 35164 125600 35176
rect 125652 35164 125658 35216
rect 204898 35164 204904 35216
rect 204956 35204 204962 35216
rect 340230 35204 340236 35216
rect 204956 35176 340236 35204
rect 204956 35164 204962 35176
rect 340230 35164 340236 35176
rect 340288 35164 340294 35216
rect 108942 33736 108948 33788
rect 109000 33776 109006 33788
rect 155218 33776 155224 33788
rect 109000 33748 155224 33776
rect 109000 33736 109006 33748
rect 155218 33736 155224 33748
rect 155276 33736 155282 33788
rect 280890 33736 280896 33788
rect 280948 33776 280954 33788
rect 325694 33776 325700 33788
rect 280948 33748 325700 33776
rect 280948 33736 280954 33748
rect 325694 33736 325700 33748
rect 325752 33736 325758 33788
rect 3510 33056 3516 33108
rect 3568 33096 3574 33108
rect 58618 33096 58624 33108
rect 3568 33068 58624 33096
rect 3568 33056 3574 33068
rect 58618 33056 58624 33068
rect 58676 33056 58682 33108
rect 70210 32376 70216 32428
rect 70268 32416 70274 32428
rect 133138 32416 133144 32428
rect 70268 32388 133144 32416
rect 70268 32376 70274 32388
rect 133138 32376 133144 32388
rect 133196 32376 133202 32428
rect 46842 31016 46848 31068
rect 46900 31056 46906 31068
rect 160830 31056 160836 31068
rect 46900 31028 160836 31056
rect 46900 31016 46906 31028
rect 160830 31016 160836 31028
rect 160888 31016 160894 31068
rect 197354 31016 197360 31068
rect 197412 31056 197418 31068
rect 342254 31056 342260 31068
rect 197412 31028 342260 31056
rect 197412 31016 197418 31028
rect 342254 31016 342260 31028
rect 342312 31016 342318 31068
rect 43990 29588 43996 29640
rect 44048 29628 44054 29640
rect 166258 29628 166264 29640
rect 44048 29600 166264 29628
rect 44048 29588 44054 29600
rect 166258 29588 166264 29600
rect 166316 29588 166322 29640
rect 209682 29588 209688 29640
rect 209740 29628 209746 29640
rect 278774 29628 278780 29640
rect 209740 29600 278780 29628
rect 209740 29588 209746 29600
rect 278774 29588 278780 29600
rect 278832 29588 278838 29640
rect 121362 28228 121368 28280
rect 121420 28268 121426 28280
rect 175918 28268 175924 28280
rect 121420 28240 175924 28268
rect 121420 28228 121426 28240
rect 175918 28228 175924 28240
rect 175976 28228 175982 28280
rect 192570 28228 192576 28280
rect 192628 28268 192634 28280
rect 328454 28268 328460 28280
rect 192628 28240 328460 28268
rect 192628 28228 192634 28240
rect 328454 28228 328460 28240
rect 328512 28228 328518 28280
rect 61930 26868 61936 26920
rect 61988 26908 61994 26920
rect 160738 26908 160744 26920
rect 61988 26880 160744 26908
rect 61988 26868 61994 26880
rect 160738 26868 160744 26880
rect 160796 26868 160802 26920
rect 229830 26868 229836 26920
rect 229888 26908 229894 26920
rect 260834 26908 260840 26920
rect 229888 26880 260840 26908
rect 229888 26868 229894 26880
rect 260834 26868 260840 26880
rect 260892 26868 260898 26920
rect 100662 25508 100668 25560
rect 100720 25548 100726 25560
rect 162118 25548 162124 25560
rect 100720 25520 162124 25548
rect 100720 25508 100726 25520
rect 162118 25508 162124 25520
rect 162176 25508 162182 25560
rect 204162 25508 204168 25560
rect 204220 25548 204226 25560
rect 324406 25548 324412 25560
rect 204220 25520 324412 25548
rect 204220 25508 204226 25520
rect 324406 25508 324412 25520
rect 324464 25508 324470 25560
rect 84010 24080 84016 24132
rect 84068 24120 84074 24132
rect 152458 24120 152464 24132
rect 84068 24092 152464 24120
rect 84068 24080 84074 24092
rect 152458 24080 152464 24092
rect 152516 24080 152522 24132
rect 206278 24080 206284 24132
rect 206336 24120 206342 24132
rect 247034 24120 247040 24132
rect 206336 24092 247040 24120
rect 206336 24080 206342 24092
rect 247034 24080 247040 24092
rect 247092 24080 247098 24132
rect 250530 24080 250536 24132
rect 250588 24120 250594 24132
rect 331214 24120 331220 24132
rect 250588 24092 331220 24120
rect 250588 24080 250594 24092
rect 331214 24080 331220 24092
rect 331272 24080 331278 24132
rect 102042 22720 102048 22772
rect 102100 22760 102106 22772
rect 141418 22760 141424 22772
rect 102100 22732 141424 22760
rect 102100 22720 102106 22732
rect 141418 22720 141424 22732
rect 141476 22720 141482 22772
rect 214558 22720 214564 22772
rect 214616 22760 214622 22772
rect 347038 22760 347044 22772
rect 214616 22732 347044 22760
rect 214616 22720 214622 22732
rect 347038 22720 347044 22732
rect 347096 22720 347102 22772
rect 86770 21360 86776 21412
rect 86828 21400 86834 21412
rect 137278 21400 137284 21412
rect 86828 21372 137284 21400
rect 86828 21360 86834 21372
rect 137278 21360 137284 21372
rect 137336 21360 137342 21412
rect 191742 21360 191748 21412
rect 191800 21400 191806 21412
rect 264974 21400 264980 21412
rect 191800 21372 264980 21400
rect 191800 21360 191806 21372
rect 264974 21360 264980 21372
rect 265032 21360 265038 21412
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 93118 20652 93124 20664
rect 3476 20624 93124 20652
rect 3476 20612 3482 20624
rect 93118 20612 93124 20624
rect 93176 20612 93182 20664
rect 93762 19932 93768 19984
rect 93820 19972 93826 19984
rect 169018 19972 169024 19984
rect 93820 19944 169024 19972
rect 93820 19932 93826 19944
rect 169018 19932 169024 19944
rect 169076 19932 169082 19984
rect 220078 19932 220084 19984
rect 220136 19972 220142 19984
rect 284386 19972 284392 19984
rect 220136 19944 284392 19972
rect 220136 19932 220142 19944
rect 284386 19932 284392 19944
rect 284444 19932 284450 19984
rect 95050 18572 95056 18624
rect 95108 18612 95114 18624
rect 130378 18612 130384 18624
rect 95108 18584 130384 18612
rect 95108 18572 95114 18584
rect 130378 18572 130384 18584
rect 130436 18572 130442 18624
rect 253290 18572 253296 18624
rect 253348 18612 253354 18624
rect 344278 18612 344284 18624
rect 253348 18584 344284 18612
rect 253348 18572 253354 18584
rect 344278 18572 344284 18584
rect 344336 18572 344342 18624
rect 99282 17280 99288 17332
rect 99340 17320 99346 17332
rect 215938 17320 215944 17332
rect 99340 17292 215944 17320
rect 99340 17280 99346 17292
rect 215938 17280 215944 17292
rect 215996 17280 216002 17332
rect 240778 17280 240784 17332
rect 240836 17320 240842 17332
rect 256694 17320 256700 17332
rect 240836 17292 256700 17320
rect 240836 17280 240842 17292
rect 256694 17280 256700 17292
rect 256752 17280 256758 17332
rect 78582 17212 78588 17264
rect 78640 17252 78646 17264
rect 126238 17252 126244 17264
rect 78640 17224 126244 17252
rect 78640 17212 78646 17224
rect 126238 17212 126244 17224
rect 126296 17212 126302 17264
rect 202782 17212 202788 17264
rect 202840 17252 202846 17264
rect 321554 17252 321560 17264
rect 202840 17224 321560 17252
rect 202840 17212 202846 17224
rect 321554 17212 321560 17224
rect 321612 17212 321618 17264
rect 68922 15852 68928 15904
rect 68980 15892 68986 15904
rect 174538 15892 174544 15904
rect 68980 15864 174544 15892
rect 68980 15852 68986 15864
rect 174538 15852 174544 15864
rect 174596 15852 174602 15904
rect 184842 15852 184848 15904
rect 184900 15892 184906 15904
rect 280706 15892 280712 15904
rect 184900 15864 280712 15892
rect 184900 15852 184906 15864
rect 280706 15852 280712 15864
rect 280764 15852 280770 15904
rect 226978 14424 226984 14476
rect 227036 14464 227042 14476
rect 303154 14464 303160 14476
rect 227036 14436 303160 14464
rect 227036 14424 227042 14436
rect 303154 14424 303160 14436
rect 303212 14424 303218 14476
rect 64782 13064 64788 13116
rect 64840 13104 64846 13116
rect 177298 13104 177304 13116
rect 64840 13076 177304 13104
rect 64840 13064 64846 13076
rect 177298 13064 177304 13076
rect 177356 13064 177362 13116
rect 181530 13064 181536 13116
rect 181588 13104 181594 13116
rect 281534 13104 281540 13116
rect 181588 13076 281540 13104
rect 181588 13064 181594 13076
rect 281534 13064 281540 13076
rect 281592 13064 281598 13116
rect 251174 11772 251180 11824
rect 251232 11812 251238 11824
rect 252370 11812 252376 11824
rect 251232 11784 252376 11812
rect 251232 11772 251238 11784
rect 252370 11772 252376 11784
rect 252428 11772 252434 11824
rect 90910 11704 90916 11756
rect 90968 11744 90974 11756
rect 153838 11744 153844 11756
rect 90968 11716 153844 11744
rect 90968 11704 90974 11716
rect 153838 11704 153844 11716
rect 153896 11704 153902 11756
rect 195238 11704 195244 11756
rect 195296 11744 195302 11756
rect 312170 11744 312176 11756
rect 195296 11716 312176 11744
rect 195296 11704 195302 11716
rect 312170 11704 312176 11716
rect 312228 11704 312234 11756
rect 332686 11704 332692 11756
rect 332744 11744 332750 11756
rect 333882 11744 333888 11756
rect 332744 11716 333888 11744
rect 332744 11704 332750 11716
rect 333882 11704 333888 11716
rect 333940 11704 333946 11756
rect 97902 10344 97908 10396
rect 97960 10384 97966 10396
rect 148318 10384 148324 10396
rect 97960 10356 148324 10384
rect 97960 10344 97966 10356
rect 148318 10344 148324 10356
rect 148376 10344 148382 10396
rect 2682 10276 2688 10328
rect 2740 10316 2746 10328
rect 101398 10316 101404 10328
rect 2740 10288 101404 10316
rect 2740 10276 2746 10288
rect 101398 10276 101404 10288
rect 101456 10276 101462 10328
rect 222838 10276 222844 10328
rect 222896 10316 222902 10328
rect 334710 10316 334716 10328
rect 222896 10288 334716 10316
rect 222896 10276 222902 10288
rect 334710 10276 334716 10288
rect 334768 10276 334774 10328
rect 271782 9596 271788 9648
rect 271840 9636 271846 9648
rect 276014 9636 276020 9648
rect 271840 9608 276020 9636
rect 271840 9596 271846 9608
rect 276014 9596 276020 9608
rect 276072 9596 276078 9648
rect 255958 8984 255964 9036
rect 256016 9024 256022 9036
rect 302418 9024 302424 9036
rect 256016 8996 302424 9024
rect 256016 8984 256022 8996
rect 302418 8984 302424 8996
rect 302476 8984 302482 9036
rect 82078 8916 82084 8968
rect 82136 8956 82142 8968
rect 170398 8956 170404 8968
rect 82136 8928 170404 8956
rect 82136 8916 82142 8928
rect 170398 8916 170404 8928
rect 170456 8916 170462 8968
rect 196618 8916 196624 8968
rect 196676 8956 196682 8968
rect 258258 8956 258264 8968
rect 196676 8928 258264 8956
rect 196676 8916 196682 8928
rect 258258 8916 258264 8928
rect 258316 8916 258322 8968
rect 100294 7556 100300 7608
rect 100352 7596 100358 7608
rect 159358 7596 159364 7608
rect 100352 7568 159364 7596
rect 100352 7556 100358 7568
rect 159358 7556 159364 7568
rect 159416 7556 159422 7608
rect 3418 6604 3424 6656
rect 3476 6644 3482 6656
rect 7558 6644 7564 6656
rect 3476 6616 7564 6644
rect 3476 6604 3482 6616
rect 7558 6604 7564 6616
rect 7616 6604 7622 6656
rect 251174 6196 251180 6248
rect 251232 6236 251238 6248
rect 263594 6236 263600 6248
rect 251232 6208 263600 6236
rect 251232 6196 251238 6208
rect 263594 6196 263600 6208
rect 263652 6196 263658 6248
rect 224862 6128 224868 6180
rect 224920 6168 224926 6180
rect 254670 6168 254676 6180
rect 224920 6140 254676 6168
rect 224920 6128 224926 6140
rect 254670 6128 254676 6140
rect 254728 6128 254734 6180
rect 256050 6128 256056 6180
rect 256108 6168 256114 6180
rect 292482 6168 292488 6180
rect 256108 6140 292488 6168
rect 256108 6128 256114 6140
rect 292482 6128 292488 6140
rect 292540 6128 292546 6180
rect 300118 5584 300124 5636
rect 300176 5624 300182 5636
rect 306742 5624 306748 5636
rect 300176 5596 306748 5624
rect 300176 5584 300182 5596
rect 306742 5584 306748 5596
rect 306800 5584 306806 5636
rect 305730 5516 305736 5568
rect 305788 5556 305794 5568
rect 309042 5556 309048 5568
rect 305788 5528 309048 5556
rect 305788 5516 305794 5528
rect 309042 5516 309048 5528
rect 309100 5516 309106 5568
rect 349798 5516 349804 5568
rect 349856 5556 349862 5568
rect 351638 5556 351644 5568
rect 349856 5528 351644 5556
rect 349856 5516 349862 5528
rect 351638 5516 351644 5528
rect 351696 5516 351702 5568
rect 96246 4836 96252 4888
rect 96304 4876 96310 4888
rect 173158 4876 173164 4888
rect 96304 4848 173164 4876
rect 96304 4836 96310 4848
rect 173158 4836 173164 4848
rect 173216 4836 173222 4888
rect 228358 4836 228364 4888
rect 228416 4876 228422 4888
rect 239306 4876 239312 4888
rect 228416 4848 239312 4876
rect 228416 4836 228422 4848
rect 239306 4836 239312 4848
rect 239364 4836 239370 4888
rect 566 4768 572 4820
rect 624 4808 630 4820
rect 97258 4808 97264 4820
rect 624 4780 97264 4808
rect 624 4768 630 4780
rect 97258 4768 97264 4780
rect 97316 4768 97322 4820
rect 238018 4768 238024 4820
rect 238076 4808 238082 4820
rect 270034 4808 270040 4820
rect 238076 4780 270040 4808
rect 238076 4768 238082 4780
rect 270034 4768 270040 4780
rect 270092 4768 270098 4820
rect 323578 4768 323584 4820
rect 323636 4808 323642 4820
rect 330386 4808 330392 4820
rect 323636 4780 330392 4808
rect 323636 4768 323642 4780
rect 330386 4768 330392 4780
rect 330444 4768 330450 4820
rect 331858 4496 331864 4548
rect 331916 4536 331922 4548
rect 337470 4536 337476 4548
rect 331916 4508 337476 4536
rect 331916 4496 331922 4508
rect 337470 4496 337476 4508
rect 337528 4496 337534 4548
rect 291838 4428 291844 4480
rect 291896 4468 291902 4480
rect 297266 4468 297272 4480
rect 291896 4440 297272 4468
rect 291896 4428 291902 4440
rect 297266 4428 297272 4440
rect 297324 4428 297330 4480
rect 134518 4156 134524 4208
rect 134576 4196 134582 4208
rect 136450 4196 136456 4208
rect 134576 4168 136456 4196
rect 134576 4156 134582 4168
rect 136450 4156 136456 4168
rect 136508 4156 136514 4208
rect 307018 4156 307024 4208
rect 307076 4196 307082 4208
rect 315022 4196 315028 4208
rect 307076 4168 315028 4196
rect 307076 4156 307082 4168
rect 315022 4156 315028 4168
rect 315080 4156 315086 4208
rect 342990 4088 342996 4140
rect 343048 4128 343054 4140
rect 346946 4128 346952 4140
rect 343048 4100 346952 4128
rect 343048 4088 343054 4100
rect 346946 4088 346952 4100
rect 347004 4088 347010 4140
rect 233878 4020 233884 4072
rect 233936 4060 233942 4072
rect 240502 4060 240508 4072
rect 233936 4032 240508 4060
rect 233936 4020 233942 4032
rect 240502 4020 240508 4032
rect 240560 4020 240566 4072
rect 8754 3544 8760 3596
rect 8812 3584 8818 3596
rect 22738 3584 22744 3596
rect 8812 3556 22744 3584
rect 8812 3544 8818 3556
rect 22738 3544 22744 3556
rect 22796 3544 22802 3596
rect 66714 3544 66720 3596
rect 66772 3584 66778 3596
rect 76558 3584 76564 3596
rect 66772 3556 76564 3584
rect 66772 3544 66778 3556
rect 76558 3544 76564 3556
rect 76616 3544 76622 3596
rect 85666 3544 85672 3596
rect 85724 3584 85730 3596
rect 86770 3584 86776 3596
rect 85724 3556 86776 3584
rect 85724 3544 85730 3556
rect 86770 3544 86776 3556
rect 86828 3544 86834 3596
rect 1670 3476 1676 3528
rect 1728 3516 1734 3528
rect 2682 3516 2688 3528
rect 1728 3488 2688 3516
rect 1728 3476 1734 3488
rect 2682 3476 2688 3488
rect 2740 3476 2746 3528
rect 2866 3476 2872 3528
rect 2924 3516 2930 3528
rect 3970 3516 3976 3528
rect 2924 3488 3976 3516
rect 2924 3476 2930 3488
rect 3970 3476 3976 3488
rect 4028 3476 4034 3528
rect 9950 3476 9956 3528
rect 10008 3516 10014 3528
rect 10962 3516 10968 3528
rect 10008 3488 10968 3516
rect 10008 3476 10014 3488
rect 10962 3476 10968 3488
rect 11020 3476 11026 3528
rect 11146 3476 11152 3528
rect 11204 3516 11210 3528
rect 12342 3516 12348 3528
rect 11204 3488 12348 3516
rect 11204 3476 11210 3488
rect 12342 3476 12348 3488
rect 12400 3476 12406 3528
rect 15930 3476 15936 3528
rect 15988 3516 15994 3528
rect 16482 3516 16488 3528
rect 15988 3488 16488 3516
rect 15988 3476 15994 3488
rect 16482 3476 16488 3488
rect 16540 3476 16546 3528
rect 17034 3476 17040 3528
rect 17092 3516 17098 3528
rect 17862 3516 17868 3528
rect 17092 3488 17868 3516
rect 17092 3476 17098 3488
rect 17862 3476 17868 3488
rect 17920 3476 17926 3528
rect 18230 3476 18236 3528
rect 18288 3516 18294 3528
rect 19242 3516 19248 3528
rect 18288 3488 19248 3516
rect 18288 3476 18294 3488
rect 19242 3476 19248 3488
rect 19300 3476 19306 3528
rect 24210 3476 24216 3528
rect 24268 3516 24274 3528
rect 24762 3516 24768 3528
rect 24268 3488 24768 3516
rect 24268 3476 24274 3488
rect 24762 3476 24768 3488
rect 24820 3476 24826 3528
rect 26510 3476 26516 3528
rect 26568 3516 26574 3528
rect 27522 3516 27528 3528
rect 26568 3488 27528 3516
rect 26568 3476 26574 3488
rect 27522 3476 27528 3488
rect 27580 3476 27586 3528
rect 32398 3476 32404 3528
rect 32456 3516 32462 3528
rect 33042 3516 33048 3528
rect 32456 3488 33048 3516
rect 32456 3476 32462 3488
rect 33042 3476 33048 3488
rect 33100 3476 33106 3528
rect 33594 3476 33600 3528
rect 33652 3516 33658 3528
rect 34422 3516 34428 3528
rect 33652 3488 34428 3516
rect 33652 3476 33658 3488
rect 34422 3476 34428 3488
rect 34480 3476 34486 3528
rect 34790 3476 34796 3528
rect 34848 3516 34854 3528
rect 35802 3516 35808 3528
rect 34848 3488 35808 3516
rect 34848 3476 34854 3488
rect 35802 3476 35808 3488
rect 35860 3476 35866 3528
rect 35986 3476 35992 3528
rect 36044 3516 36050 3528
rect 37090 3516 37096 3528
rect 36044 3488 37096 3516
rect 36044 3476 36050 3488
rect 37090 3476 37096 3488
rect 37148 3476 37154 3528
rect 40678 3476 40684 3528
rect 40736 3516 40742 3528
rect 41138 3516 41144 3528
rect 40736 3488 41144 3516
rect 40736 3476 40742 3488
rect 41138 3476 41144 3488
rect 41196 3476 41202 3528
rect 41874 3476 41880 3528
rect 41932 3516 41938 3528
rect 42702 3516 42708 3528
rect 41932 3488 42708 3516
rect 41932 3476 41938 3488
rect 42702 3476 42708 3488
rect 42760 3476 42766 3528
rect 43070 3476 43076 3528
rect 43128 3516 43134 3528
rect 43990 3516 43996 3528
rect 43128 3488 43996 3516
rect 43128 3476 43134 3488
rect 43990 3476 43996 3488
rect 44048 3476 44054 3528
rect 48958 3476 48964 3528
rect 49016 3516 49022 3528
rect 49602 3516 49608 3528
rect 49016 3488 49608 3516
rect 49016 3476 49022 3488
rect 49602 3476 49608 3488
rect 49660 3476 49666 3528
rect 50154 3476 50160 3528
rect 50212 3516 50218 3528
rect 50706 3516 50712 3528
rect 50212 3488 50712 3516
rect 50212 3476 50218 3488
rect 50706 3476 50712 3488
rect 50764 3476 50770 3528
rect 52546 3476 52552 3528
rect 52604 3516 52610 3528
rect 53650 3516 53656 3528
rect 52604 3488 53656 3516
rect 52604 3476 52610 3488
rect 53650 3476 53656 3488
rect 53708 3476 53714 3528
rect 57238 3476 57244 3528
rect 57296 3516 57302 3528
rect 57882 3516 57888 3528
rect 57296 3488 57888 3516
rect 57296 3476 57302 3488
rect 57882 3476 57888 3488
rect 57940 3476 57946 3528
rect 58434 3476 58440 3528
rect 58492 3516 58498 3528
rect 59262 3516 59268 3528
rect 58492 3488 59268 3516
rect 58492 3476 58498 3488
rect 59262 3476 59268 3488
rect 59320 3476 59326 3528
rect 59630 3476 59636 3528
rect 59688 3516 59694 3528
rect 60642 3516 60648 3528
rect 59688 3488 60648 3516
rect 59688 3476 59694 3488
rect 60642 3476 60648 3488
rect 60700 3476 60706 3528
rect 60826 3476 60832 3528
rect 60884 3516 60890 3528
rect 61930 3516 61936 3528
rect 60884 3488 61936 3516
rect 60884 3476 60890 3488
rect 61930 3476 61936 3488
rect 61988 3476 61994 3528
rect 64322 3476 64328 3528
rect 64380 3516 64386 3528
rect 64782 3516 64788 3528
rect 64380 3488 64788 3516
rect 64380 3476 64386 3488
rect 64782 3476 64788 3488
rect 64840 3476 64846 3528
rect 65518 3476 65524 3528
rect 65576 3516 65582 3528
rect 66162 3516 66168 3528
rect 65576 3488 66168 3516
rect 65576 3476 65582 3488
rect 66162 3476 66168 3488
rect 66220 3476 66226 3528
rect 67910 3476 67916 3528
rect 67968 3516 67974 3528
rect 68922 3516 68928 3528
rect 67968 3488 68928 3516
rect 67968 3476 67974 3488
rect 68922 3476 68928 3488
rect 68980 3476 68986 3528
rect 69106 3476 69112 3528
rect 69164 3516 69170 3528
rect 70210 3516 70216 3528
rect 69164 3488 70216 3516
rect 69164 3476 69170 3488
rect 70210 3476 70216 3488
rect 70268 3476 70274 3528
rect 72602 3476 72608 3528
rect 72660 3516 72666 3528
rect 73062 3516 73068 3528
rect 72660 3488 73068 3516
rect 72660 3476 72666 3488
rect 73062 3476 73068 3488
rect 73120 3476 73126 3528
rect 74994 3476 75000 3528
rect 75052 3516 75058 3528
rect 75822 3516 75828 3528
rect 75052 3488 75828 3516
rect 75052 3476 75058 3488
rect 75822 3476 75828 3488
rect 75880 3476 75886 3528
rect 76190 3476 76196 3528
rect 76248 3516 76254 3528
rect 77202 3516 77208 3528
rect 76248 3488 77208 3516
rect 76248 3476 76254 3488
rect 77202 3476 77208 3488
rect 77260 3476 77266 3528
rect 80882 3476 80888 3528
rect 80940 3516 80946 3528
rect 81342 3516 81348 3528
rect 80940 3488 81348 3516
rect 80940 3476 80946 3488
rect 81342 3476 81348 3488
rect 81400 3476 81406 3528
rect 89162 3476 89168 3528
rect 89220 3516 89226 3528
rect 89622 3516 89628 3528
rect 89220 3488 89628 3516
rect 89220 3476 89226 3488
rect 89622 3476 89628 3488
rect 89680 3476 89686 3528
rect 90358 3476 90364 3528
rect 90416 3516 90422 3528
rect 90910 3516 90916 3528
rect 90416 3488 90916 3516
rect 90416 3476 90422 3488
rect 90910 3476 90916 3488
rect 90968 3476 90974 3528
rect 91002 3476 91008 3528
rect 91060 3516 91066 3528
rect 91554 3516 91560 3528
rect 91060 3488 91560 3516
rect 91060 3476 91066 3488
rect 91554 3476 91560 3488
rect 91612 3476 91618 3528
rect 92750 3476 92756 3528
rect 92808 3516 92814 3528
rect 93762 3516 93768 3528
rect 92808 3488 93768 3516
rect 92808 3476 92814 3488
rect 93762 3476 93768 3488
rect 93820 3476 93826 3528
rect 93946 3476 93952 3528
rect 94004 3516 94010 3528
rect 95050 3516 95056 3528
rect 94004 3488 95056 3516
rect 94004 3476 94010 3488
rect 95050 3476 95056 3488
rect 95108 3476 95114 3528
rect 97442 3476 97448 3528
rect 97500 3516 97506 3528
rect 97902 3516 97908 3528
rect 97500 3488 97908 3516
rect 97500 3476 97506 3488
rect 97902 3476 97908 3488
rect 97960 3476 97966 3528
rect 98638 3476 98644 3528
rect 98696 3516 98702 3528
rect 99282 3516 99288 3528
rect 98696 3488 99288 3516
rect 98696 3476 98702 3488
rect 99282 3476 99288 3488
rect 99340 3476 99346 3528
rect 99834 3476 99840 3528
rect 99892 3516 99898 3528
rect 100662 3516 100668 3528
rect 99892 3488 100668 3516
rect 99892 3476 99898 3488
rect 100662 3476 100668 3488
rect 100720 3476 100726 3528
rect 101030 3476 101036 3528
rect 101088 3516 101094 3528
rect 102042 3516 102048 3528
rect 101088 3488 102048 3516
rect 101088 3476 101094 3488
rect 102042 3476 102048 3488
rect 102100 3476 102106 3528
rect 102226 3476 102232 3528
rect 102284 3516 102290 3528
rect 106826 3516 106832 3528
rect 102284 3488 106832 3516
rect 102284 3476 102290 3488
rect 106826 3476 106832 3488
rect 106884 3476 106890 3528
rect 106918 3476 106924 3528
rect 106976 3516 106982 3528
rect 107562 3516 107568 3528
rect 106976 3488 107568 3516
rect 106976 3476 106982 3488
rect 107562 3476 107568 3488
rect 107620 3476 107626 3528
rect 108114 3476 108120 3528
rect 108172 3516 108178 3528
rect 108942 3516 108948 3528
rect 108172 3488 108948 3516
rect 108172 3476 108178 3488
rect 108942 3476 108948 3488
rect 109000 3476 109006 3528
rect 109310 3476 109316 3528
rect 109368 3516 109374 3528
rect 110322 3516 110328 3528
rect 109368 3488 110328 3516
rect 109368 3476 109374 3488
rect 110322 3476 110328 3488
rect 110380 3476 110386 3528
rect 114002 3476 114008 3528
rect 114060 3516 114066 3528
rect 114462 3516 114468 3528
rect 114060 3488 114468 3516
rect 114060 3476 114066 3488
rect 114462 3476 114468 3488
rect 114520 3476 114526 3528
rect 115198 3476 115204 3528
rect 115256 3516 115262 3528
rect 115842 3516 115848 3528
rect 115256 3488 115848 3516
rect 115256 3476 115262 3488
rect 115842 3476 115848 3488
rect 115900 3476 115906 3528
rect 116394 3476 116400 3528
rect 116452 3516 116458 3528
rect 117222 3516 117228 3528
rect 116452 3488 117228 3516
rect 116452 3476 116458 3488
rect 117222 3476 117228 3488
rect 117280 3476 117286 3528
rect 117590 3476 117596 3528
rect 117648 3516 117654 3528
rect 118602 3516 118608 3528
rect 117648 3488 118608 3516
rect 117648 3476 117654 3488
rect 118602 3476 118608 3488
rect 118660 3476 118666 3528
rect 122282 3476 122288 3528
rect 122340 3516 122346 3528
rect 122742 3516 122748 3528
rect 122340 3488 122748 3516
rect 122340 3476 122346 3488
rect 122742 3476 122748 3488
rect 122800 3476 122806 3528
rect 123478 3476 123484 3528
rect 123536 3516 123542 3528
rect 124122 3516 124128 3528
rect 123536 3488 124128 3516
rect 123536 3476 123542 3488
rect 124122 3476 124128 3488
rect 124180 3476 124186 3528
rect 124674 3476 124680 3528
rect 124732 3516 124738 3528
rect 125502 3516 125508 3528
rect 124732 3488 125508 3516
rect 124732 3476 124738 3488
rect 125502 3476 125508 3488
rect 125560 3476 125566 3528
rect 143534 3476 143540 3528
rect 143592 3516 143598 3528
rect 144822 3516 144828 3528
rect 143592 3488 144828 3516
rect 143592 3476 143598 3488
rect 144822 3476 144828 3488
rect 144880 3476 144886 3528
rect 147122 3476 147128 3528
rect 147180 3516 147186 3528
rect 147582 3516 147588 3528
rect 147180 3488 147588 3516
rect 147180 3476 147186 3488
rect 147582 3476 147588 3488
rect 147640 3476 147646 3528
rect 249058 3476 249064 3528
rect 249116 3516 249122 3528
rect 255866 3516 255872 3528
rect 249116 3488 255872 3516
rect 249116 3476 249122 3488
rect 255866 3476 255872 3488
rect 255924 3476 255930 3528
rect 260098 3476 260104 3528
rect 260156 3516 260162 3528
rect 267734 3516 267740 3528
rect 260156 3488 267740 3516
rect 260156 3476 260162 3488
rect 267734 3476 267740 3488
rect 267792 3476 267798 3528
rect 280798 3476 280804 3528
rect 280856 3516 280862 3528
rect 287790 3516 287796 3528
rect 280856 3488 287796 3516
rect 280856 3476 280862 3488
rect 287790 3476 287796 3488
rect 287848 3476 287854 3528
rect 299474 3476 299480 3528
rect 299532 3516 299538 3528
rect 300762 3516 300768 3528
rect 299532 3488 300768 3516
rect 299532 3476 299538 3488
rect 300762 3476 300768 3488
rect 300820 3476 300826 3528
rect 302418 3476 302424 3528
rect 302476 3516 302482 3528
rect 305546 3516 305552 3528
rect 302476 3488 305552 3516
rect 302476 3476 302482 3488
rect 305546 3476 305552 3488
rect 305604 3476 305610 3528
rect 324314 3476 324320 3528
rect 324372 3516 324378 3528
rect 325602 3516 325608 3528
rect 324372 3488 325608 3516
rect 324372 3476 324378 3488
rect 325602 3476 325608 3488
rect 325660 3476 325666 3528
rect 340138 3476 340144 3528
rect 340196 3516 340202 3528
rect 342162 3516 342168 3528
rect 340196 3488 342168 3516
rect 340196 3476 340202 3488
rect 342162 3476 342168 3488
rect 342220 3476 342226 3528
rect 1302 3408 1308 3460
rect 1360 3448 1366 3460
rect 1360 3420 12388 3448
rect 1360 3408 1366 3420
rect 12360 3392 12388 3420
rect 13538 3408 13544 3460
rect 13596 3448 13602 3460
rect 32306 3448 32312 3460
rect 13596 3420 32312 3448
rect 13596 3408 13602 3420
rect 32306 3408 32312 3420
rect 32364 3408 32370 3460
rect 51350 3408 51356 3460
rect 51408 3448 51414 3460
rect 66898 3448 66904 3460
rect 51408 3420 66904 3448
rect 51408 3408 51414 3420
rect 66898 3408 66904 3420
rect 66956 3408 66962 3460
rect 83274 3408 83280 3460
rect 83332 3448 83338 3460
rect 84010 3448 84016 3460
rect 83332 3420 84016 3448
rect 83332 3408 83338 3420
rect 84010 3408 84016 3420
rect 84068 3408 84074 3460
rect 98546 3448 98552 3460
rect 84166 3420 98552 3448
rect 12342 3340 12348 3392
rect 12400 3340 12406 3392
rect 27706 3340 27712 3392
rect 27764 3380 27770 3392
rect 33778 3380 33784 3392
rect 27764 3352 33784 3380
rect 27764 3340 27770 3352
rect 33778 3340 33784 3352
rect 33836 3340 33842 3392
rect 77386 3340 77392 3392
rect 77444 3380 77450 3392
rect 84166 3380 84194 3420
rect 98546 3408 98552 3420
rect 98604 3408 98610 3460
rect 105722 3408 105728 3460
rect 105780 3448 105786 3460
rect 115106 3448 115112 3460
rect 105780 3420 115112 3448
rect 105780 3408 105786 3420
rect 115106 3408 115112 3420
rect 115164 3408 115170 3460
rect 213178 3408 213184 3460
rect 213236 3448 213242 3460
rect 242894 3448 242900 3460
rect 213236 3420 242900 3448
rect 213236 3408 213242 3420
rect 242894 3408 242900 3420
rect 242952 3408 242958 3460
rect 246298 3408 246304 3460
rect 246356 3448 246362 3460
rect 253474 3448 253480 3460
rect 246356 3420 253480 3448
rect 246356 3408 246362 3420
rect 253474 3408 253480 3420
rect 253532 3408 253538 3460
rect 266998 3408 267004 3460
rect 267056 3448 267062 3460
rect 273622 3448 273628 3460
rect 267056 3420 273628 3448
rect 267056 3408 267062 3420
rect 273622 3408 273628 3420
rect 273680 3408 273686 3460
rect 320818 3408 320824 3460
rect 320876 3448 320882 3460
rect 332686 3448 332692 3460
rect 320876 3420 332692 3448
rect 320876 3408 320882 3420
rect 332686 3408 332692 3420
rect 332744 3408 332750 3460
rect 334710 3408 334716 3460
rect 334768 3448 334774 3460
rect 339862 3448 339868 3460
rect 334768 3420 339868 3448
rect 334768 3408 334774 3420
rect 339862 3408 339868 3420
rect 339920 3408 339926 3460
rect 344278 3408 344284 3460
rect 344336 3448 344342 3460
rect 350442 3448 350448 3460
rect 344336 3420 350448 3448
rect 344336 3408 344342 3420
rect 350442 3408 350448 3420
rect 350500 3408 350506 3460
rect 574738 3408 574744 3460
rect 574796 3448 574802 3460
rect 582190 3448 582196 3460
rect 574796 3420 582196 3448
rect 574796 3408 574802 3420
rect 582190 3408 582196 3420
rect 582248 3408 582254 3460
rect 77444 3352 84194 3380
rect 77444 3340 77450 3352
rect 253198 3340 253204 3392
rect 253256 3380 253262 3392
rect 264146 3380 264152 3392
rect 253256 3352 264152 3380
rect 253256 3340 253262 3352
rect 264146 3340 264152 3352
rect 264204 3340 264210 3392
rect 309870 3340 309876 3392
rect 309928 3380 309934 3392
rect 311434 3380 311440 3392
rect 309928 3352 311440 3380
rect 309928 3340 309934 3352
rect 311434 3340 311440 3352
rect 311492 3340 311498 3392
rect 289078 3272 289084 3324
rect 289136 3312 289142 3324
rect 292574 3312 292580 3324
rect 289136 3284 292580 3312
rect 289136 3272 289142 3284
rect 292574 3272 292580 3284
rect 292632 3272 292638 3324
rect 340230 3272 340236 3324
rect 340288 3312 340294 3324
rect 344554 3312 344560 3324
rect 340288 3284 344560 3312
rect 340288 3272 340294 3284
rect 344554 3272 344560 3284
rect 344612 3272 344618 3324
rect 317322 3204 317328 3256
rect 317380 3244 317386 3256
rect 321646 3244 321652 3256
rect 317380 3216 321652 3244
rect 317380 3204 317386 3216
rect 321646 3204 321652 3216
rect 321704 3204 321710 3256
rect 580994 3204 581000 3256
rect 581052 3244 581058 3256
rect 582466 3244 582472 3256
rect 581052 3216 582472 3244
rect 581052 3204 581058 3216
rect 582466 3204 582472 3216
rect 582524 3204 582530 3256
rect 25314 3136 25320 3188
rect 25372 3176 25378 3188
rect 26142 3176 26148 3188
rect 25372 3148 26148 3176
rect 25372 3136 25378 3148
rect 26142 3136 26148 3148
rect 26200 3136 26206 3188
rect 118786 3068 118792 3120
rect 118844 3108 118850 3120
rect 119798 3108 119804 3120
rect 118844 3080 119804 3108
rect 118844 3068 118850 3080
rect 119798 3068 119804 3080
rect 119856 3068 119862 3120
rect 299658 3068 299664 3120
rect 299716 3108 299722 3120
rect 302234 3108 302240 3120
rect 299716 3080 302240 3108
rect 299716 3068 299722 3080
rect 302234 3068 302240 3080
rect 302292 3068 302298 3120
rect 347038 3068 347044 3120
rect 347096 3108 347102 3120
rect 349246 3108 349252 3120
rect 347096 3080 349252 3108
rect 347096 3068 347102 3080
rect 349246 3068 349252 3080
rect 349304 3068 349310 3120
rect 55122 3000 55128 3052
rect 55180 3040 55186 3052
rect 56042 3040 56048 3052
rect 55180 3012 56048 3040
rect 55180 3000 55186 3012
rect 56042 3000 56048 3012
rect 56100 3000 56106 3052
rect 258718 3000 258724 3052
rect 258776 3040 258782 3052
rect 260650 3040 260656 3052
rect 258776 3012 260656 3040
rect 258776 3000 258782 3012
rect 260650 3000 260656 3012
rect 260708 3000 260714 3052
rect 304258 3000 304264 3052
rect 304316 3040 304322 3052
rect 307938 3040 307944 3052
rect 304316 3012 307944 3040
rect 304316 3000 304322 3012
rect 307938 3000 307944 3012
rect 307996 3000 308002 3052
rect 282178 2932 282184 2984
rect 282236 2972 282242 2984
rect 283098 2972 283104 2984
rect 282236 2944 283104 2972
rect 282236 2932 282242 2944
rect 283098 2932 283104 2944
rect 283156 2932 283162 2984
rect 292482 2932 292488 2984
rect 292540 2972 292546 2984
rect 294874 2972 294880 2984
rect 292540 2944 294880 2972
rect 292540 2932 292546 2944
rect 294874 2932 294880 2944
rect 294932 2932 294938 2984
rect 270034 2796 270040 2848
rect 270092 2836 270098 2848
rect 272426 2836 272432 2848
rect 270092 2808 272432 2836
rect 270092 2796 270098 2808
rect 272426 2796 272432 2808
rect 272484 2796 272490 2848
rect 140038 2728 140044 2780
rect 140096 2768 140102 2780
rect 142982 2768 142988 2780
rect 140096 2740 142988 2768
rect 140096 2728 140102 2740
rect 142982 2728 142988 2740
rect 143040 2728 143046 2780
rect 7650 2048 7656 2100
rect 7708 2088 7714 2100
rect 17218 2088 17224 2100
rect 7708 2060 17224 2088
rect 7708 2048 7714 2060
rect 17218 2048 17224 2060
rect 17276 2048 17282 2100
rect 19426 2048 19432 2100
rect 19484 2088 19490 2100
rect 178678 2088 178684 2100
rect 19484 2060 178684 2088
rect 19484 2048 19490 2060
rect 178678 2048 178684 2060
rect 178736 2048 178742 2100
<< via1 >>
rect 191748 703332 191800 703384
rect 283840 703332 283892 703384
rect 273904 703264 273956 703316
rect 348792 703264 348844 703316
rect 215208 703196 215260 703248
rect 364984 703196 365036 703248
rect 240784 703128 240836 703180
rect 332508 703128 332560 703180
rect 249708 703060 249760 703112
rect 413652 703060 413704 703112
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 220084 702992 220136 703044
rect 267648 702992 267700 703044
rect 282184 702992 282236 703044
rect 462320 702992 462372 703044
rect 104808 702924 104860 702976
rect 300124 702924 300176 702976
rect 24308 702856 24360 702908
rect 86224 702856 86276 702908
rect 90364 702856 90416 702908
rect 235172 702856 235224 702908
rect 271144 702856 271196 702908
rect 478512 702856 478564 702908
rect 70308 702788 70360 702840
rect 154120 702788 154172 702840
rect 213184 702788 213236 702840
rect 429844 702788 429896 702840
rect 40500 702720 40552 702772
rect 94688 702720 94740 702772
rect 173808 702720 173860 702772
rect 397460 702720 397512 702772
rect 8116 702652 8168 702704
rect 96620 702652 96672 702704
rect 280804 702652 280856 702704
rect 543464 702652 543516 702704
rect 84108 702584 84160 702636
rect 202788 702584 202840 702636
rect 215944 702584 215996 702636
rect 527088 702584 527140 702636
rect 66168 702516 66220 702568
rect 170312 702516 170364 702568
rect 177948 702516 178000 702568
rect 580908 702516 580960 702568
rect 77208 702448 77260 702500
rect 494796 702448 494848 702500
rect 79968 700272 80020 700324
rect 89168 700272 89220 700324
rect 218980 700272 219032 700324
rect 241520 700272 241572 700324
rect 3424 683136 3476 683188
rect 39304 683136 39356 683188
rect 3516 670692 3568 670744
rect 14464 670692 14516 670744
rect 3424 656888 3476 656940
rect 74540 656888 74592 656940
rect 68928 625812 68980 625864
rect 104900 625812 104952 625864
rect 3516 618264 3568 618316
rect 11704 618264 11756 618316
rect 2780 605888 2832 605940
rect 4804 605888 4856 605940
rect 79324 592016 79376 592068
rect 79968 592016 80020 592068
rect 112444 592016 112496 592068
rect 76472 590384 76524 590436
rect 77208 590384 77260 590436
rect 76472 589296 76524 589348
rect 124404 589296 124456 589348
rect 67732 588344 67784 588396
rect 68928 588344 68980 588396
rect 68928 587868 68980 587920
rect 128360 587868 128412 587920
rect 81808 587188 81860 587240
rect 84108 587188 84160 587240
rect 143540 587188 143592 587240
rect 4804 587120 4856 587172
rect 96712 587120 96764 587172
rect 121460 585760 121512 585812
rect 582840 585760 582892 585812
rect 87512 585216 87564 585268
rect 121460 585216 121512 585268
rect 72424 585148 72476 585200
rect 116584 585148 116636 585200
rect 74264 583788 74316 583840
rect 98644 583788 98696 583840
rect 88248 583720 88300 583772
rect 115204 583720 115256 583772
rect 78128 582632 78180 582684
rect 79324 582632 79376 582684
rect 57888 582564 57940 582616
rect 90456 582564 90508 582616
rect 86224 582496 86276 582548
rect 100208 582496 100260 582548
rect 50988 582428 51040 582480
rect 69940 582428 69992 582480
rect 79048 582360 79100 582412
rect 86868 582360 86920 582412
rect 90272 582360 90324 582412
rect 95976 582360 96028 582412
rect 76288 581068 76340 581120
rect 108304 581068 108356 581120
rect 59268 581000 59320 581052
rect 83004 581000 83056 581052
rect 93768 581000 93820 581052
rect 148324 581000 148376 581052
rect 69020 580660 69072 580712
rect 86868 580660 86920 580712
rect 3516 580184 3568 580236
rect 8116 580184 8168 580236
rect 64788 579708 64840 579760
rect 66536 579708 66588 579760
rect 53564 579640 53616 579692
rect 94688 580456 94740 580508
rect 95884 580456 95936 580508
rect 102784 580252 102836 580304
rect 97172 578212 97224 578264
rect 134524 578212 134576 578264
rect 97172 576852 97224 576904
rect 122840 576852 122892 576904
rect 187608 576852 187660 576904
rect 580172 576852 580224 576904
rect 3424 576784 3476 576836
rect 67640 576784 67692 576836
rect 97908 576104 97960 576156
rect 104808 576104 104860 576156
rect 125600 576104 125652 576156
rect 95976 574744 96028 574796
rect 104164 574744 104216 574796
rect 95884 573316 95936 573368
rect 120080 573316 120132 573368
rect 63408 572704 63460 572756
rect 66536 572704 66588 572756
rect 41328 571344 41380 571396
rect 66536 571344 66588 571396
rect 96804 571344 96856 571396
rect 106924 571344 106976 571396
rect 61936 569984 61988 570036
rect 66904 569984 66956 570036
rect 97908 569916 97960 569968
rect 115296 569916 115348 569968
rect 97908 568624 97960 568676
rect 104440 568624 104492 568676
rect 62028 565836 62080 565888
rect 66168 565836 66220 565888
rect 56508 564408 56560 564460
rect 66536 564408 66588 564460
rect 52368 563048 52420 563100
rect 66536 563048 66588 563100
rect 107016 562912 107068 562964
rect 111064 562912 111116 562964
rect 96804 561688 96856 561740
rect 117320 561688 117372 561740
rect 48044 560260 48096 560312
rect 66720 560260 66772 560312
rect 48228 558900 48280 558952
rect 66720 558900 66772 558952
rect 96804 558900 96856 558952
rect 112720 558900 112772 558952
rect 44088 557540 44140 557592
rect 66720 557540 66772 557592
rect 96988 554752 97040 554804
rect 129740 554752 129792 554804
rect 3332 553392 3384 553444
rect 29644 553392 29696 553444
rect 57796 553392 57848 553444
rect 66536 553392 66588 553444
rect 96988 552032 97040 552084
rect 108488 552032 108540 552084
rect 97908 550604 97960 550656
rect 115940 550604 115992 550656
rect 55128 549244 55180 549296
rect 66536 549244 66588 549296
rect 64696 547884 64748 547936
rect 66812 547884 66864 547936
rect 63316 545096 63368 545148
rect 66720 545096 66772 545148
rect 97080 543736 97132 543788
rect 104348 543736 104400 543788
rect 39304 543668 39356 543720
rect 67272 543668 67324 543720
rect 97172 540948 97224 541000
rect 130384 540948 130436 541000
rect 11704 540200 11756 540252
rect 73160 539792 73212 539844
rect 91008 539792 91060 539844
rect 96712 539792 96764 539844
rect 59176 539588 59228 539640
rect 66444 539588 66496 539640
rect 86224 539588 86276 539640
rect 94320 539588 94372 539640
rect 67824 539044 67876 539096
rect 71872 539044 71924 539096
rect 82728 538840 82780 538892
rect 95516 538840 95568 538892
rect 4804 538228 4856 538280
rect 93952 538228 94004 538280
rect 29644 538160 29696 538212
rect 70676 538160 70728 538212
rect 90364 538160 90416 538212
rect 136640 538160 136692 538212
rect 75828 537480 75880 537532
rect 96896 537480 96948 537532
rect 3424 536732 3476 536784
rect 69020 536732 69072 536784
rect 73436 536732 73488 536784
rect 76564 536732 76616 536784
rect 82176 536120 82228 536172
rect 95332 536120 95384 536172
rect 67732 536052 67784 536104
rect 83464 536052 83516 536104
rect 86684 535508 86736 535560
rect 87696 535508 87748 535560
rect 50804 534692 50856 534744
rect 87144 534692 87196 534744
rect 88340 533400 88392 533452
rect 88892 533400 88944 533452
rect 91100 533400 91152 533452
rect 91836 533400 91888 533452
rect 55036 533332 55088 533384
rect 96804 533332 96856 533384
rect 65892 531972 65944 532024
rect 107016 531972 107068 532024
rect 93768 531224 93820 531276
rect 94504 531224 94556 531276
rect 70676 530544 70728 530596
rect 141424 530544 141476 530596
rect 3424 529184 3476 529236
rect 93768 529184 93820 529236
rect 3516 527824 3568 527876
rect 122840 527824 122892 527876
rect 64604 526396 64656 526448
rect 84200 526396 84252 526448
rect 67364 525036 67416 525088
rect 113180 525036 113232 525088
rect 104348 521568 104400 521620
rect 108396 521568 108448 521620
rect 64696 520888 64748 520940
rect 69664 520888 69716 520940
rect 53656 518168 53708 518220
rect 98000 518168 98052 518220
rect 3516 514768 3568 514820
rect 7564 514768 7616 514820
rect 108488 506948 108540 507000
rect 112536 506948 112588 507000
rect 66076 501576 66128 501628
rect 125784 501576 125836 501628
rect 88432 498788 88484 498840
rect 124312 498788 124364 498840
rect 63316 496068 63368 496120
rect 123484 496068 123536 496120
rect 76564 493280 76616 493332
rect 102876 493280 102928 493332
rect 64788 490560 64840 490612
rect 92480 490560 92532 490612
rect 73804 487772 73856 487824
rect 99380 487772 99432 487824
rect 102140 487772 102192 487824
rect 102784 487772 102836 487824
rect 240784 487772 240836 487824
rect 77300 486412 77352 486464
rect 108488 486412 108540 486464
rect 77944 485052 77996 485104
rect 91192 485052 91244 485104
rect 188988 484372 189040 484424
rect 580172 484372 580224 484424
rect 112444 483624 112496 483676
rect 125692 483624 125744 483676
rect 87696 481584 87748 481636
rect 88248 481584 88300 481636
rect 241520 481584 241572 481636
rect 242164 481584 242216 481636
rect 88248 480904 88300 480956
rect 242164 480904 242216 480956
rect 67732 479476 67784 479528
rect 96988 479476 97040 479528
rect 90456 478864 90508 478916
rect 91008 478864 91060 478916
rect 218060 478864 218112 478916
rect 106924 478116 106976 478168
rect 128452 478116 128504 478168
rect 2780 476076 2832 476128
rect 3424 476076 3476 476128
rect 4804 476076 4856 476128
rect 104164 476076 104216 476128
rect 241520 476076 241572 476128
rect 78680 475396 78732 475448
rect 98736 475396 98788 475448
rect 98644 475328 98696 475380
rect 121552 475328 121604 475380
rect 104256 475192 104308 475244
rect 104808 475192 104860 475244
rect 104808 474716 104860 474768
rect 255412 474716 255464 474768
rect 93952 473832 94004 473884
rect 94688 473832 94740 473884
rect 94688 473356 94740 473408
rect 227812 473356 227864 473408
rect 88340 472608 88392 472660
rect 118700 472608 118752 472660
rect 118700 471996 118752 472048
rect 255596 471996 255648 472048
rect 108488 471248 108540 471300
rect 117412 471248 117464 471300
rect 117412 470568 117464 470620
rect 262220 470568 262272 470620
rect 82820 469820 82872 469872
rect 109684 469820 109736 469872
rect 159364 469276 159416 469328
rect 253940 469276 253992 469328
rect 112444 469208 112496 469260
rect 142896 469208 142948 469260
rect 252560 469208 252612 469260
rect 71688 468528 71740 468580
rect 91100 468528 91152 468580
rect 85580 468460 85632 468512
rect 113364 468460 113416 468512
rect 108396 467848 108448 467900
rect 245660 467848 245712 467900
rect 82728 466488 82780 466540
rect 211160 466488 211212 466540
rect 102416 466420 102468 466472
rect 102876 466420 102928 466472
rect 240876 466420 240928 466472
rect 87604 465672 87656 465724
rect 126980 465672 127032 465724
rect 188344 465128 188396 465180
rect 256700 465128 256752 465180
rect 137284 465060 137336 465112
rect 240140 465060 240192 465112
rect 57704 464992 57756 465044
rect 57888 464992 57940 465044
rect 86868 464312 86920 464364
rect 95240 464312 95292 464364
rect 141424 463768 141476 463820
rect 259552 463768 259604 463820
rect 57704 463700 57756 463752
rect 186964 463700 187016 463752
rect 191196 463700 191248 463752
rect 231124 463700 231176 463752
rect 77208 462952 77260 463004
rect 90364 462952 90416 463004
rect 92388 462408 92440 462460
rect 225604 462408 225656 462460
rect 3516 462340 3568 462392
rect 32404 462340 32456 462392
rect 223580 462340 223632 462392
rect 291200 462340 291252 462392
rect 80060 461592 80112 461644
rect 113272 461592 113324 461644
rect 285680 461592 285732 461644
rect 583208 461592 583260 461644
rect 166908 460980 166960 461032
rect 233240 460980 233292 461032
rect 75184 460912 75236 460964
rect 75828 460912 75880 460964
rect 195980 460912 196032 460964
rect 202144 460912 202196 460964
rect 285680 460912 285732 460964
rect 184848 459620 184900 459672
rect 233332 459620 233384 459672
rect 119344 459552 119396 459604
rect 258264 459552 258316 459604
rect 95240 458260 95292 458312
rect 197084 458260 197136 458312
rect 227720 458260 227772 458312
rect 85488 458192 85540 458244
rect 86224 458192 86276 458244
rect 148324 458192 148376 458244
rect 256792 458192 256844 458244
rect 192484 456900 192536 456952
rect 218888 456900 218940 456952
rect 72424 456832 72476 456884
rect 157340 456832 157392 456884
rect 197360 456832 197412 456884
rect 226432 456832 226484 456884
rect 260840 456832 260892 456884
rect 78680 456764 78732 456816
rect 175188 456764 175240 456816
rect 204444 456764 204496 456816
rect 247408 456764 247460 456816
rect 288348 456764 288400 456816
rect 580172 456764 580224 456816
rect 68928 456016 68980 456068
rect 80060 456016 80112 456068
rect 190368 455472 190420 455524
rect 204536 455472 204588 455524
rect 236000 455472 236052 455524
rect 260104 455472 260156 455524
rect 192576 455404 192628 455456
rect 213184 455404 213236 455456
rect 237380 455404 237432 455456
rect 273352 455404 273404 455456
rect 74540 455336 74592 455388
rect 75368 455336 75420 455388
rect 88248 454656 88300 454708
rect 104900 454656 104952 454708
rect 75368 454112 75420 454164
rect 151084 454112 151136 454164
rect 193404 454112 193456 454164
rect 237840 454112 237892 454164
rect 240784 454112 240836 454164
rect 276020 454112 276072 454164
rect 116676 454044 116728 454096
rect 245752 454044 245804 454096
rect 239220 453976 239272 454028
rect 240784 453976 240836 454028
rect 240140 453432 240192 453484
rect 240876 453432 240928 453484
rect 231676 453364 231728 453416
rect 237380 453364 237432 453416
rect 232596 452752 232648 452804
rect 82820 452684 82872 452736
rect 168288 452684 168340 452736
rect 200396 452684 200448 452736
rect 201592 452684 201644 452736
rect 205916 452684 205968 452736
rect 75276 452616 75328 452668
rect 201316 452616 201368 452668
rect 202788 452616 202840 452668
rect 209780 452616 209832 452668
rect 227720 452616 227772 452668
rect 229652 452616 229704 452668
rect 240140 452684 240192 452736
rect 259460 452684 259512 452736
rect 269120 452616 269172 452668
rect 111800 452548 111852 452600
rect 112444 452548 112496 452600
rect 191104 451868 191156 451920
rect 202788 451868 202840 451920
rect 104256 451324 104308 451376
rect 137284 451324 137336 451376
rect 248788 451324 248840 451376
rect 254032 451324 254084 451376
rect 39304 451256 39356 451308
rect 111800 451256 111852 451308
rect 122104 451256 122156 451308
rect 142068 451256 142120 451308
rect 184388 451256 184440 451308
rect 199292 451256 199344 451308
rect 204076 451256 204128 451308
rect 277400 451256 277452 451308
rect 87604 449964 87656 450016
rect 214196 449964 214248 450016
rect 218612 449964 218664 450016
rect 270500 449964 270552 450016
rect 67272 449896 67324 449948
rect 94780 449896 94832 449948
rect 95148 449896 95200 449948
rect 98644 449896 98696 449948
rect 232228 449896 232280 449948
rect 233148 449896 233200 449948
rect 244556 449896 244608 449948
rect 262864 449896 262916 449948
rect 191472 449828 191524 449880
rect 246028 449828 246080 449880
rect 251824 449692 251876 449744
rect 41328 449148 41380 449200
rect 106924 449148 106976 449200
rect 185584 449148 185636 449200
rect 193404 449148 193456 449200
rect 281632 448944 281684 448996
rect 3148 448536 3200 448588
rect 11704 448536 11756 448588
rect 61936 448536 61988 448588
rect 169024 448536 169076 448588
rect 176568 448536 176620 448588
rect 191656 448536 191708 448588
rect 67640 448332 67692 448384
rect 75368 448332 75420 448384
rect 73252 447788 73304 447840
rect 82820 447788 82872 447840
rect 95148 447788 95200 447840
rect 170404 447788 170456 447840
rect 178960 447788 179012 447840
rect 192576 447788 192628 447840
rect 82912 447108 82964 447160
rect 83464 447108 83516 447160
rect 178960 447108 179012 447160
rect 179236 447108 179288 447160
rect 172428 446360 172480 446412
rect 192484 446360 192536 446412
rect 253848 446360 253900 446412
rect 267740 446360 267792 446412
rect 37096 445816 37148 445868
rect 77300 445816 77352 445868
rect 77944 445816 77996 445868
rect 66168 445748 66220 445800
rect 191748 445748 191800 445800
rect 50988 445680 51040 445732
rect 95148 445680 95200 445732
rect 83464 444388 83516 444440
rect 176660 444388 176712 444440
rect 191748 444388 191800 444440
rect 188436 444320 188488 444372
rect 190460 444320 190512 444372
rect 69112 443640 69164 443692
rect 166264 443640 166316 443692
rect 255688 443640 255740 443692
rect 284300 443640 284352 443692
rect 33784 442960 33836 443012
rect 95332 442960 95384 443012
rect 255412 442960 255464 443012
rect 258816 442960 258868 443012
rect 88432 442892 88484 442944
rect 92572 442892 92624 442944
rect 48136 442212 48188 442264
rect 52368 442212 52420 442264
rect 88432 442212 88484 442264
rect 254676 442212 254728 442264
rect 271880 442212 271932 442264
rect 67456 441600 67508 441652
rect 162124 441600 162176 441652
rect 7564 441532 7616 441584
rect 104164 441532 104216 441584
rect 161388 440852 161440 440904
rect 191288 440852 191340 440904
rect 63316 440240 63368 440292
rect 191196 440240 191248 440292
rect 67180 439492 67232 439544
rect 83464 439492 83516 439544
rect 104808 439492 104860 439544
rect 114652 439492 114704 439544
rect 255412 439492 255464 439544
rect 258264 439492 258316 439544
rect 288624 439492 288676 439544
rect 582932 439492 582984 439544
rect 73988 438880 74040 438932
rect 75276 438880 75328 438932
rect 82912 438880 82964 438932
rect 180064 438880 180116 438932
rect 48044 438812 48096 438864
rect 74724 438812 74776 438864
rect 75368 438812 75420 438864
rect 94504 438812 94556 438864
rect 97356 438812 97408 438864
rect 255504 438812 255556 438864
rect 262220 438812 262272 438864
rect 70492 437452 70544 437504
rect 191748 437452 191800 437504
rect 262220 437452 262272 437504
rect 263692 437452 263744 437504
rect 82820 437384 82872 437436
rect 83924 437384 83976 437436
rect 87604 437384 87656 437436
rect 97356 437384 97408 437436
rect 98644 437384 98696 437436
rect 98736 437384 98788 437436
rect 103704 437384 103756 437436
rect 104256 437384 104308 437436
rect 108304 437384 108356 437436
rect 122104 437384 122156 437436
rect 255504 437384 255556 437436
rect 582380 437384 582432 437436
rect 107384 436704 107436 436756
rect 116676 436704 116728 436756
rect 87328 436432 87380 436484
rect 90456 436432 90508 436484
rect 53748 436160 53800 436212
rect 69848 436160 69900 436212
rect 17224 436092 17276 436144
rect 70860 436160 70912 436212
rect 75184 436160 75236 436212
rect 75644 436160 75696 436212
rect 78036 436160 78088 436212
rect 71688 436092 71740 436144
rect 72424 436092 72476 436144
rect 72516 436092 72568 436144
rect 77484 436092 77536 436144
rect 92388 436092 92440 436144
rect 94228 436092 94280 436144
rect 107568 435412 107620 435464
rect 116032 435412 116084 435464
rect 55036 435344 55088 435396
rect 191748 435344 191800 435396
rect 255412 435344 255464 435396
rect 259552 435344 259604 435396
rect 274640 435344 274692 435396
rect 137376 434868 137428 434920
rect 141424 434868 141476 434920
rect 64696 434732 64748 434784
rect 73988 434732 74040 434784
rect 115020 434664 115072 434716
rect 178684 434664 178736 434716
rect 188436 434664 188488 434716
rect 188896 434664 188948 434716
rect 191748 434664 191800 434716
rect 255412 434596 255464 434648
rect 258080 434596 258132 434648
rect 265072 434596 265124 434648
rect 100208 433984 100260 434036
rect 115388 433984 115440 434036
rect 64788 433304 64840 433356
rect 191656 433304 191708 433356
rect 68652 433236 68704 433288
rect 188896 433236 188948 433288
rect 255964 432624 256016 432676
rect 262220 432624 262272 432676
rect 254584 432556 254636 432608
rect 283012 432556 283064 432608
rect 187424 431944 187476 431996
rect 191104 431944 191156 431996
rect 115296 431264 115348 431316
rect 118700 431264 118752 431316
rect 171048 431196 171100 431248
rect 180156 431196 180208 431248
rect 115848 430244 115900 430296
rect 119436 430244 119488 430296
rect 255136 429836 255188 429888
rect 258724 429836 258776 429888
rect 258816 429836 258868 429888
rect 270592 429836 270644 429888
rect 61936 429088 61988 429140
rect 66812 429088 66864 429140
rect 151084 429088 151136 429140
rect 191564 429088 191616 429140
rect 115848 428408 115900 428460
rect 122932 428408 122984 428460
rect 123484 428408 123536 428460
rect 46848 427796 46900 427848
rect 66260 427796 66312 427848
rect 255412 427796 255464 427848
rect 264980 427796 265032 427848
rect 115848 427728 115900 427780
rect 159364 427728 159416 427780
rect 255504 427728 255556 427780
rect 260932 427728 260984 427780
rect 262128 427728 262180 427780
rect 169024 427048 169076 427100
rect 176752 427048 176804 427100
rect 262128 427048 262180 427100
rect 279332 427048 279384 427100
rect 50896 426436 50948 426488
rect 66904 426436 66956 426488
rect 176752 426436 176804 426488
rect 177856 426436 177908 426488
rect 191564 426436 191616 426488
rect 279332 426436 279384 426488
rect 582656 426436 582708 426488
rect 115296 426096 115348 426148
rect 119344 426096 119396 426148
rect 57888 425688 57940 425740
rect 66076 425688 66128 425740
rect 66628 425688 66680 425740
rect 181444 425076 181496 425128
rect 191012 425076 191064 425128
rect 115296 424940 115348 424992
rect 117412 424940 117464 424992
rect 157248 424328 157300 424380
rect 181536 424328 181588 424380
rect 256792 424328 256844 424380
rect 266360 424328 266412 424380
rect 114652 423716 114704 423768
rect 116032 423716 116084 423768
rect 55036 423648 55088 423700
rect 66812 423648 66864 423700
rect 3516 423580 3568 423632
rect 39304 423580 39356 423632
rect 52368 423580 52420 423632
rect 54944 423580 54996 423632
rect 66628 423580 66680 423632
rect 115848 423580 115900 423632
rect 137376 423580 137428 423632
rect 137928 422900 137980 422952
rect 148324 422900 148376 422952
rect 170404 422900 170456 422952
rect 170956 422900 171008 422952
rect 190828 422900 190880 422952
rect 255504 422288 255556 422340
rect 276112 422288 276164 422340
rect 64788 422220 64840 422272
rect 66812 422220 66864 422272
rect 48044 421540 48096 421592
rect 57704 421540 57756 421592
rect 255504 420928 255556 420980
rect 280160 420928 280212 420980
rect 173164 419568 173216 419620
rect 191564 419568 191616 419620
rect 63132 419500 63184 419552
rect 66904 419500 66956 419552
rect 115848 419500 115900 419552
rect 180156 419500 180208 419552
rect 255596 419500 255648 419552
rect 266452 419500 266504 419552
rect 63316 419432 63368 419484
rect 66812 419432 66864 419484
rect 286048 418752 286100 418804
rect 583024 418752 583076 418804
rect 184296 418140 184348 418192
rect 191564 418140 191616 418192
rect 255504 418140 255556 418192
rect 285680 418140 285732 418192
rect 286048 418140 286100 418192
rect 115204 418072 115256 418124
rect 188344 418072 188396 418124
rect 115848 418004 115900 418056
rect 133144 418004 133196 418056
rect 263784 417460 263836 417512
rect 271144 417460 271196 417512
rect 167644 417392 167696 417444
rect 184388 417392 184440 417444
rect 262128 417392 262180 417444
rect 583116 417392 583168 417444
rect 255596 416848 255648 416900
rect 260932 416848 260984 416900
rect 262128 416848 262180 416900
rect 187700 416780 187752 416832
rect 191564 416780 191616 416832
rect 255504 416780 255556 416832
rect 263784 416780 263836 416832
rect 179328 416100 179380 416152
rect 188988 416100 189040 416152
rect 191012 416100 191064 416152
rect 118700 416032 118752 416084
rect 137928 416032 137980 416084
rect 159456 416032 159508 416084
rect 187700 416032 187752 416084
rect 39948 415420 40000 415472
rect 57796 415420 57848 415472
rect 66904 415420 66956 415472
rect 115848 415420 115900 415472
rect 118700 415420 118752 415472
rect 130384 414672 130436 414724
rect 191564 414672 191616 414724
rect 64788 413992 64840 414044
rect 66720 413992 66772 414044
rect 115848 413788 115900 413840
rect 117320 413788 117372 413840
rect 49608 413244 49660 413296
rect 59268 413244 59320 413296
rect 66260 413244 66312 413296
rect 50804 412564 50856 412616
rect 66812 412564 66864 412616
rect 162124 412020 162176 412072
rect 162768 412020 162820 412072
rect 41328 411884 41380 411936
rect 50804 411884 50856 411936
rect 162768 411884 162820 411936
rect 191472 411884 191524 411936
rect 255504 411544 255556 411596
rect 258080 411544 258132 411596
rect 2964 411204 3016 411256
rect 33784 411204 33836 411256
rect 50988 410524 51040 410576
rect 62028 410524 62080 410576
rect 66904 410524 66956 410576
rect 255504 409912 255556 409964
rect 258264 409912 258316 409964
rect 115848 409844 115900 409896
rect 155224 409844 155276 409896
rect 187516 409844 187568 409896
rect 190828 409844 190880 409896
rect 52460 409776 52512 409828
rect 53656 409776 53708 409828
rect 66812 409776 66864 409828
rect 44088 409096 44140 409148
rect 52460 409096 52512 409148
rect 115848 409096 115900 409148
rect 124864 409096 124916 409148
rect 126888 408552 126940 408604
rect 143540 408552 143592 408604
rect 144184 408552 144236 408604
rect 115848 408484 115900 408536
rect 188344 408484 188396 408536
rect 255504 408484 255556 408536
rect 276204 408484 276256 408536
rect 255504 407192 255556 407244
rect 259552 407192 259604 407244
rect 52276 407124 52328 407176
rect 66812 407124 66864 407176
rect 115848 407124 115900 407176
rect 170404 407124 170456 407176
rect 162124 405764 162176 405816
rect 191472 405764 191524 405816
rect 115756 405696 115808 405748
rect 169024 405696 169076 405748
rect 255504 405696 255556 405748
rect 274732 405696 274784 405748
rect 115848 405628 115900 405680
rect 126888 405628 126940 405680
rect 62028 404336 62080 404388
rect 66904 404336 66956 404388
rect 182916 404336 182968 404388
rect 191380 404336 191432 404388
rect 255504 403384 255556 403436
rect 257344 403384 257396 403436
rect 159364 403044 159416 403096
rect 191472 403044 191524 403096
rect 54944 402976 54996 403028
rect 66812 402976 66864 403028
rect 115848 402976 115900 403028
rect 185768 402976 185820 403028
rect 114744 401344 114796 401396
rect 116676 401344 116728 401396
rect 118792 400868 118844 400920
rect 128360 400868 128412 400920
rect 187608 400732 187660 400784
rect 191472 400732 191524 400784
rect 53656 400188 53708 400240
rect 66720 400188 66772 400240
rect 115664 400188 115716 400240
rect 152464 400188 152516 400240
rect 184388 400188 184440 400240
rect 187608 400188 187660 400240
rect 255504 400188 255556 400240
rect 277492 400188 277544 400240
rect 289728 399440 289780 399492
rect 582748 399440 582800 399492
rect 115848 398828 115900 398880
rect 151084 398828 151136 398880
rect 174544 398828 174596 398880
rect 190828 398828 190880 398880
rect 255504 398828 255556 398880
rect 258356 398828 258408 398880
rect 288716 398828 288768 398880
rect 289728 398828 289780 398880
rect 291108 398080 291160 398132
rect 582472 398080 582524 398132
rect 115572 397536 115624 397588
rect 117964 397536 118016 397588
rect 118792 397536 118844 397588
rect 180248 397536 180300 397588
rect 191104 397536 191156 397588
rect 7564 397468 7616 397520
rect 67732 397468 67784 397520
rect 113824 397468 113876 397520
rect 188528 397468 188580 397520
rect 255504 397468 255556 397520
rect 289820 397468 289872 397520
rect 291108 397468 291160 397520
rect 176752 397400 176804 397452
rect 177948 397400 178000 397452
rect 191472 397400 191524 397452
rect 115848 396312 115900 396364
rect 122104 396312 122156 396364
rect 127624 396040 127676 396092
rect 191196 396040 191248 396092
rect 191380 396040 191432 396092
rect 64604 395428 64656 395480
rect 67180 395428 67232 395480
rect 115848 394680 115900 394732
rect 181536 394680 181588 394732
rect 60556 393388 60608 393440
rect 65892 393388 65944 393440
rect 129004 393388 129056 393440
rect 193404 393388 193456 393440
rect 59084 393320 59136 393372
rect 66812 393320 66864 393372
rect 115848 393320 115900 393372
rect 188436 393320 188488 393372
rect 255596 393320 255648 393372
rect 271972 393320 272024 393372
rect 115848 392572 115900 392624
rect 122840 392572 122892 392624
rect 123484 392572 123536 392624
rect 56416 391960 56468 392012
rect 66260 391960 66312 392012
rect 188528 391892 188580 391944
rect 191472 391892 191524 391944
rect 253572 391552 253624 391604
rect 254032 391552 254084 391604
rect 250536 390940 250588 390992
rect 258080 390940 258132 390992
rect 114836 390736 114888 390788
rect 116584 390736 116636 390788
rect 67364 390600 67416 390652
rect 73804 390600 73856 390652
rect 191012 390600 191064 390652
rect 203524 390600 203576 390652
rect 69664 390532 69716 390584
rect 163596 390532 163648 390584
rect 194140 390532 194192 390584
rect 96712 390464 96764 390516
rect 97540 390464 97592 390516
rect 67640 390124 67692 390176
rect 68790 390124 68842 390176
rect 56508 389784 56560 389836
rect 86776 389784 86828 389836
rect 87788 389784 87840 389836
rect 242164 389784 242216 389836
rect 254124 389784 254176 389836
rect 75092 389240 75144 389292
rect 164976 389240 165028 389292
rect 202052 389240 202104 389292
rect 249248 389240 249300 389292
rect 253664 389240 253716 389292
rect 94688 389172 94740 389224
rect 227720 389172 227772 389224
rect 228548 389172 228600 389224
rect 234896 389172 234948 389224
rect 249708 389172 249760 389224
rect 65984 389104 66036 389156
rect 71688 389104 71740 389156
rect 72608 389104 72660 389156
rect 111892 389104 111944 389156
rect 251824 389104 251876 389156
rect 241980 389036 242032 389088
rect 273904 389036 273956 389088
rect 234068 388696 234120 388748
rect 234528 388696 234580 388748
rect 239036 388696 239088 388748
rect 120724 388016 120776 388068
rect 121552 388016 121604 388068
rect 57704 387812 57756 387864
rect 66076 387812 66128 387864
rect 121460 387812 121512 387864
rect 129096 387812 129148 387864
rect 129740 387812 129792 387864
rect 214564 387812 214616 387864
rect 216220 387812 216272 387864
rect 232504 387812 232556 387864
rect 233332 387812 233384 387864
rect 241980 387812 242032 387864
rect 242808 387812 242860 387864
rect 3424 387744 3476 387796
rect 93952 387744 94004 387796
rect 94504 387744 94556 387796
rect 99472 387744 99524 387796
rect 104164 387744 104216 387796
rect 108948 387744 109000 387796
rect 114652 387744 114704 387796
rect 118792 387744 118844 387796
rect 218244 387744 218296 387796
rect 219256 387744 219308 387796
rect 101680 387676 101732 387728
rect 125600 387676 125652 387728
rect 126244 387676 126296 387728
rect 180156 387676 180208 387728
rect 255412 387676 255464 387728
rect 219256 387064 219308 387116
rect 232596 387064 232648 387116
rect 253388 387064 253440 387116
rect 267832 387064 267884 387116
rect 77300 386996 77352 387048
rect 78036 386996 78088 387048
rect 84200 386996 84252 387048
rect 85028 386996 85080 387048
rect 109040 386996 109092 387048
rect 109500 386996 109552 387048
rect 223580 386996 223632 387048
rect 224500 386996 224552 387048
rect 67824 386316 67876 386368
rect 174544 386316 174596 386368
rect 186964 386316 187016 386368
rect 208492 386316 208544 386368
rect 231124 386316 231176 386368
rect 234252 386316 234304 386368
rect 103152 385636 103204 385688
rect 187608 385636 187660 385688
rect 89628 385024 89680 385076
rect 94320 385024 94372 385076
rect 231860 385024 231912 385076
rect 281724 385024 281776 385076
rect 86868 384956 86920 385008
rect 118792 384956 118844 385008
rect 190276 384956 190328 385008
rect 216404 384956 216456 385008
rect 100392 384888 100444 384940
rect 126888 384888 126940 384940
rect 119988 384276 120040 384328
rect 186320 384276 186372 384328
rect 221004 384276 221056 384328
rect 244924 384276 244976 384328
rect 259552 384276 259604 384328
rect 216404 383664 216456 383716
rect 240232 383664 240284 383716
rect 242992 383664 243044 383716
rect 243820 383664 243872 383716
rect 244004 383664 244056 383716
rect 247684 383664 247736 383716
rect 98000 383596 98052 383648
rect 120724 383596 120776 383648
rect 67732 382984 67784 383036
rect 83464 382984 83516 383036
rect 80060 382916 80112 382968
rect 106372 382916 106424 382968
rect 115940 382916 115992 382968
rect 125508 382916 125560 382968
rect 231860 382916 231912 382968
rect 282920 382916 282972 382968
rect 283104 382916 283156 382968
rect 582840 382916 582892 382968
rect 239404 382304 239456 382356
rect 244280 382304 244332 382356
rect 226984 382236 227036 382288
rect 273536 382236 273588 382288
rect 97724 382168 97776 382220
rect 124220 382168 124272 382220
rect 125508 382168 125560 382220
rect 187608 382168 187660 382220
rect 239128 382168 239180 382220
rect 111892 381692 111944 381744
rect 112720 381692 112772 381744
rect 65984 381488 66036 381540
rect 77392 381488 77444 381540
rect 188436 381488 188488 381540
rect 223488 381488 223540 381540
rect 3424 380876 3476 380928
rect 111892 380876 111944 380928
rect 230756 380876 230808 380928
rect 273444 380876 273496 380928
rect 50988 380808 51040 380860
rect 184296 380808 184348 380860
rect 189080 380808 189132 380860
rect 189724 380808 189776 380860
rect 221280 380808 221332 380860
rect 223488 380808 223540 380860
rect 251916 380808 251968 380860
rect 109132 380128 109184 380180
rect 163504 380128 163556 380180
rect 246396 380128 246448 380180
rect 254216 380128 254268 380180
rect 50712 379516 50764 379568
rect 50988 379516 51040 379568
rect 52276 379448 52328 379500
rect 130384 379448 130436 379500
rect 240232 379448 240284 379500
rect 582932 379448 582984 379500
rect 92480 379380 92532 379432
rect 125692 379380 125744 379432
rect 126428 379380 126480 379432
rect 129096 379380 129148 379432
rect 204260 379380 204312 379432
rect 185768 379312 185820 379364
rect 244924 379312 244976 379364
rect 245752 378156 245804 378208
rect 246304 378156 246356 378208
rect 269304 378156 269356 378208
rect 67272 378088 67324 378140
rect 162124 378088 162176 378140
rect 188344 378088 188396 378140
rect 188896 378088 188948 378140
rect 256700 378088 256752 378140
rect 84292 377408 84344 377460
rect 97264 377408 97316 377460
rect 97632 377408 97684 377460
rect 118700 377408 118752 377460
rect 230756 377408 230808 377460
rect 256700 376728 256752 376780
rect 257344 376728 257396 376780
rect 291292 376728 291344 376780
rect 73804 376592 73856 376644
rect 159364 376592 159416 376644
rect 117964 376524 118016 376576
rect 277492 376524 277544 376576
rect 58900 375980 58952 376032
rect 76564 375980 76616 376032
rect 105544 375980 105596 376032
rect 117964 375980 118016 376032
rect 88248 375300 88300 375352
rect 91928 375300 91980 375352
rect 224960 375300 225012 375352
rect 72976 375232 73028 375284
rect 168380 375232 168432 375284
rect 181536 375232 181588 375284
rect 255504 375232 255556 375284
rect 170404 373940 170456 373992
rect 242164 373940 242216 373992
rect 94504 373260 94556 373312
rect 121460 373260 121512 373312
rect 226984 373260 227036 373312
rect 240784 373260 240836 373312
rect 262220 373260 262272 373312
rect 106096 372512 106148 372564
rect 242900 372512 242952 372564
rect 163504 372444 163556 372496
rect 248420 372444 248472 372496
rect 250444 372444 250496 372496
rect 81440 371832 81492 371884
rect 115940 371832 115992 371884
rect 117228 371832 117280 371884
rect 242900 371220 242952 371272
rect 243544 371220 243596 371272
rect 102048 371152 102100 371204
rect 236000 371152 236052 371204
rect 81256 370472 81308 370524
rect 129096 370472 129148 370524
rect 187424 370472 187476 370524
rect 198004 370472 198056 370524
rect 236000 369860 236052 369912
rect 236644 369860 236696 369912
rect 111892 369792 111944 369844
rect 274732 369792 274784 369844
rect 151084 369724 151136 369776
rect 245844 369724 245896 369776
rect 245844 369316 245896 369368
rect 246396 369316 246448 369368
rect 101404 369112 101456 369164
rect 111892 369112 111944 369164
rect 126428 368432 126480 368484
rect 226340 368432 226392 368484
rect 226984 368432 227036 368484
rect 67640 368364 67692 368416
rect 129004 368364 129056 368416
rect 152464 368364 152516 368416
rect 252560 368364 252612 368416
rect 59084 367004 59136 367056
rect 88984 366936 89036 366988
rect 183560 367004 183612 367056
rect 184388 367004 184440 367056
rect 189080 366936 189132 366988
rect 183560 366800 183612 366852
rect 188804 366324 188856 366376
rect 207112 366324 207164 366376
rect 108856 365644 108908 365696
rect 246304 365644 246356 365696
rect 86776 364964 86828 365016
rect 129004 364964 129056 365016
rect 170496 364352 170548 364404
rect 213828 364352 213880 364404
rect 116584 364284 116636 364336
rect 254032 364284 254084 364336
rect 71688 363604 71740 363656
rect 195888 363604 195940 363656
rect 254032 362924 254084 362976
rect 259552 362924 259604 362976
rect 77300 362856 77352 362908
rect 205732 362856 205784 362908
rect 213828 362856 213880 362908
rect 231124 362856 231176 362908
rect 195888 362788 195940 362840
rect 198740 362788 198792 362840
rect 86868 362176 86920 362228
rect 187700 362176 187752 362228
rect 198740 362176 198792 362228
rect 293960 362176 294012 362228
rect 69020 361496 69072 361548
rect 194600 361496 194652 361548
rect 123484 360816 123536 360868
rect 271972 360816 272024 360868
rect 69020 360476 69072 360528
rect 69756 360476 69808 360528
rect 124864 360136 124916 360188
rect 245660 360136 245712 360188
rect 97264 360068 97316 360120
rect 215392 360068 215444 360120
rect 215392 359660 215444 359712
rect 215944 359660 215996 359712
rect 245660 359660 245712 359712
rect 246304 359660 246356 359712
rect 82820 359456 82872 359508
rect 103520 359456 103572 359508
rect 243544 359456 243596 359508
rect 260932 359456 260984 359508
rect 104164 358708 104216 358760
rect 234620 358708 234672 358760
rect 235264 358708 235316 358760
rect 3240 358640 3292 358692
rect 7564 358640 7616 358692
rect 104716 357348 104768 357400
rect 242808 357348 242860 357400
rect 242808 356668 242860 356720
rect 254584 356668 254636 356720
rect 129096 355988 129148 356040
rect 211160 355988 211212 356040
rect 211804 355988 211856 356040
rect 129004 354016 129056 354068
rect 152556 354016 152608 354068
rect 216680 354016 216732 354068
rect 84200 353948 84252 354000
rect 164884 353948 164936 354000
rect 214564 353948 214616 354000
rect 115388 353200 115440 353252
rect 249248 353200 249300 353252
rect 218060 352520 218112 352572
rect 249156 352520 249208 352572
rect 193036 351228 193088 351280
rect 242992 351228 243044 351280
rect 169668 351160 169720 351212
rect 178684 351160 178736 351212
rect 187424 351160 187476 351212
rect 258172 351160 258224 351212
rect 169576 349800 169628 349852
rect 253480 349800 253532 349852
rect 115204 349052 115256 349104
rect 250536 349052 250588 349104
rect 202880 348372 202932 348424
rect 252744 348372 252796 348424
rect 192852 347012 192904 347064
rect 238116 347012 238168 347064
rect 177948 345652 178000 345704
rect 239404 345652 239456 345704
rect 3424 345312 3476 345364
rect 7564 345312 7616 345364
rect 198096 344292 198148 344344
rect 250536 344292 250588 344344
rect 209780 342864 209832 342916
rect 281816 342864 281868 342916
rect 247684 341572 247736 341624
rect 258172 341572 258224 341624
rect 196624 341504 196676 341556
rect 251916 341504 251968 341556
rect 173348 340892 173400 340944
rect 244280 340892 244332 340944
rect 187516 340144 187568 340196
rect 240876 340144 240928 340196
rect 92480 339464 92532 339516
rect 266452 339464 266504 339516
rect 73068 338104 73120 338156
rect 270684 338104 270736 338156
rect 236644 337356 236696 337408
rect 262312 337356 262364 337408
rect 130476 336744 130528 336796
rect 252560 336744 252612 336796
rect 169668 335996 169720 336048
rect 205640 335996 205692 336048
rect 236644 335996 236696 336048
rect 137284 335316 137336 335368
rect 253296 335316 253348 335368
rect 193404 334568 193456 334620
rect 229100 334568 229152 334620
rect 252468 334568 252520 334620
rect 260840 334568 260892 334620
rect 35808 333956 35860 334008
rect 220084 333956 220136 334008
rect 223672 333208 223724 333260
rect 238116 333208 238168 333260
rect 189908 332664 189960 332716
rect 190368 332664 190420 332716
rect 274824 332664 274876 332716
rect 12348 332596 12400 332648
rect 197360 332596 197412 332648
rect 193036 331848 193088 331900
rect 233884 331848 233936 331900
rect 238024 331848 238076 331900
rect 291384 331848 291436 331900
rect 138664 331236 138716 331288
rect 211252 331236 211304 331288
rect 142804 329876 142856 329928
rect 209044 329876 209096 329928
rect 223488 329876 223540 329928
rect 259644 329876 259696 329928
rect 102876 329808 102928 329860
rect 240232 329808 240284 329860
rect 240784 329808 240836 329860
rect 180156 329128 180208 329180
rect 265164 329128 265216 329180
rect 129004 329060 129056 329112
rect 255412 329060 255464 329112
rect 258264 329060 258316 329112
rect 226984 327700 227036 327752
rect 254768 327700 254820 327752
rect 174544 327156 174596 327208
rect 256700 327156 256752 327208
rect 37188 327088 37240 327140
rect 204260 327088 204312 327140
rect 251824 326408 251876 326460
rect 266452 326408 266504 326460
rect 68652 326340 68704 326392
rect 167644 326340 167696 326392
rect 234528 326340 234580 326392
rect 252008 326340 252060 326392
rect 126888 325660 126940 325712
rect 250628 325660 250680 325712
rect 144276 324912 144328 324964
rect 215944 324912 215996 324964
rect 228364 324912 228416 324964
rect 278872 324912 278924 324964
rect 174636 324300 174688 324352
rect 175188 324300 175240 324352
rect 280436 324300 280488 324352
rect 79324 323552 79376 323604
rect 159364 323552 159416 323604
rect 198740 323552 198792 323604
rect 255688 323552 255740 323604
rect 151176 323008 151228 323060
rect 198740 323008 198792 323060
rect 161940 322940 161992 322992
rect 162124 322940 162176 322992
rect 261024 322940 261076 322992
rect 116584 322192 116636 322244
rect 158720 322192 158772 322244
rect 263876 322192 263928 322244
rect 107568 322124 107620 322176
rect 115296 322124 115348 322176
rect 141516 321580 141568 321632
rect 142068 321580 142120 321632
rect 265256 321580 265308 321632
rect 116032 321512 116084 321564
rect 276112 321512 276164 321564
rect 104164 320832 104216 320884
rect 137284 320832 137336 320884
rect 98000 320152 98052 320204
rect 180156 320152 180208 320204
rect 270500 320152 270552 320204
rect 142896 320084 142948 320136
rect 143448 320084 143500 320136
rect 100760 320016 100812 320068
rect 102692 320016 102744 320068
rect 126888 320016 126940 320068
rect 127624 320016 127676 320068
rect 4068 319404 4120 319456
rect 17224 319404 17276 319456
rect 143448 319404 143500 319456
rect 211804 319404 211856 319456
rect 231124 319404 231176 319456
rect 272524 319404 272576 319456
rect 178776 318792 178828 318844
rect 179236 318792 179288 318844
rect 229744 318792 229796 318844
rect 265072 318724 265124 318776
rect 265348 318724 265400 318776
rect 183008 317500 183060 317552
rect 265348 317500 265400 317552
rect 82728 317432 82780 317484
rect 233884 317432 233936 317484
rect 101588 316684 101640 316736
rect 113272 316684 113324 316736
rect 135996 316684 136048 316736
rect 259460 316684 259512 316736
rect 177856 316004 177908 316056
rect 277584 316004 277636 316056
rect 229744 315256 229796 315308
rect 256884 315256 256936 315308
rect 153844 314712 153896 314764
rect 214288 314712 214340 314764
rect 67456 314644 67508 314696
rect 268016 314644 268068 314696
rect 250536 314032 250588 314084
rect 256976 314032 257028 314084
rect 171968 313352 172020 313404
rect 174544 313352 174596 313404
rect 192484 313352 192536 313404
rect 200120 313352 200172 313404
rect 201408 313352 201460 313404
rect 87604 313284 87656 313336
rect 88248 313284 88300 313336
rect 266544 313284 266596 313336
rect 167736 311924 167788 311976
rect 168288 311924 168340 311976
rect 226984 311924 227036 311976
rect 244556 311924 244608 311976
rect 244924 311924 244976 311976
rect 262404 311924 262456 311976
rect 181536 311856 181588 311908
rect 278964 311856 279016 311908
rect 193312 311108 193364 311160
rect 205732 311108 205784 311160
rect 281448 311108 281500 311160
rect 580264 311108 580316 311160
rect 266360 310972 266412 311024
rect 266636 310972 266688 311024
rect 210424 310564 210476 310616
rect 255412 310564 255464 310616
rect 174544 310496 174596 310548
rect 266636 310496 266688 310548
rect 201408 309816 201460 309868
rect 232504 309816 232556 309868
rect 41328 309748 41380 309800
rect 172612 309748 172664 309800
rect 173164 309748 173216 309800
rect 223580 309748 223632 309800
rect 255504 309748 255556 309800
rect 262864 309748 262916 309800
rect 264980 309748 265032 309800
rect 287336 309748 287388 309800
rect 155224 309136 155276 309188
rect 217416 309136 217468 309188
rect 240140 308456 240192 308508
rect 258356 308456 258408 308508
rect 230480 308388 230532 308440
rect 255596 308388 255648 308440
rect 171140 307844 171192 307896
rect 215300 307844 215352 307896
rect 151084 307776 151136 307828
rect 219716 307776 219768 307828
rect 220084 307708 220136 307760
rect 224776 307708 224828 307760
rect 63408 307028 63460 307080
rect 116584 307028 116636 307080
rect 236644 307028 236696 307080
rect 241796 307028 241848 307080
rect 244464 307028 244516 307080
rect 262220 307028 262272 307080
rect 148324 306416 148376 306468
rect 215944 306416 215996 306468
rect 117228 306348 117280 306400
rect 239312 306348 239364 306400
rect 242164 306348 242216 306400
rect 276296 306348 276348 306400
rect 226984 305600 227036 305652
rect 259460 305600 259512 305652
rect 141424 305056 141476 305108
rect 216588 305056 216640 305108
rect 3240 304988 3292 305040
rect 18604 304988 18656 305040
rect 77300 304988 77352 305040
rect 86224 304988 86276 305040
rect 142896 304988 142948 305040
rect 219072 304988 219124 305040
rect 250628 304988 250680 305040
rect 252928 304988 252980 305040
rect 209044 304512 209096 304564
rect 212172 304512 212224 304564
rect 86776 304308 86828 304360
rect 95332 304308 95384 304360
rect 130384 304308 130436 304360
rect 171140 304308 171192 304360
rect 232504 304308 232556 304360
rect 252652 304308 252704 304360
rect 253204 304308 253256 304360
rect 262864 304308 262916 304360
rect 60556 304240 60608 304292
rect 181536 304240 181588 304292
rect 247500 304240 247552 304292
rect 252468 304240 252520 304292
rect 295432 304240 295484 304292
rect 108856 303968 108908 304020
rect 115388 303968 115440 304020
rect 182824 303764 182876 303816
rect 231032 303764 231084 303816
rect 189816 303696 189868 303748
rect 196348 303696 196400 303748
rect 197360 303628 197412 303680
rect 198004 303628 198056 303680
rect 200212 303628 200264 303680
rect 201132 303628 201184 303680
rect 230112 303628 230164 303680
rect 238668 303628 238720 303680
rect 244280 303628 244332 303680
rect 244556 303628 244608 303680
rect 201408 303560 201460 303612
rect 210424 303560 210476 303612
rect 153108 302880 153160 302932
rect 192484 302880 192536 302932
rect 192760 302268 192812 302320
rect 198832 302268 198884 302320
rect 250628 302268 250680 302320
rect 260840 302268 260892 302320
rect 115296 302200 115348 302252
rect 118792 302200 118844 302252
rect 180248 302200 180300 302252
rect 218428 302200 218480 302252
rect 252008 302200 252060 302252
rect 253020 302200 253072 302252
rect 241060 302132 241112 302184
rect 253664 302132 253716 302184
rect 253296 301520 253348 301572
rect 254124 301520 254176 301572
rect 91192 301452 91244 301504
rect 135996 301452 136048 301504
rect 191472 301452 191524 301504
rect 191748 301452 191800 301504
rect 191748 301316 191800 301368
rect 196716 301316 196768 301368
rect 175924 300908 175976 300960
rect 191104 300976 191156 301028
rect 159456 300840 159508 300892
rect 240140 301316 240192 301368
rect 246488 301316 246540 301368
rect 249156 301316 249208 301368
rect 253112 301316 253164 301368
rect 178040 300772 178092 300824
rect 178776 300772 178828 300824
rect 192208 300772 192260 300824
rect 195060 300772 195112 300824
rect 93952 300160 94004 300212
rect 95056 300160 95108 300212
rect 186964 299888 187016 299940
rect 187608 299888 187660 299940
rect 191748 299888 191800 299940
rect 77944 299548 77996 299600
rect 178040 299548 178092 299600
rect 95056 299480 95108 299532
rect 147036 299480 147088 299532
rect 149796 299480 149848 299532
rect 206468 300772 206520 300824
rect 252836 300772 252888 300824
rect 256608 299548 256660 299600
rect 288532 299548 288584 299600
rect 256516 299480 256568 299532
rect 289820 299480 289872 299532
rect 105636 299412 105688 299464
rect 107568 299412 107620 299464
rect 190644 299412 190696 299464
rect 272524 299412 272576 299464
rect 580172 299412 580224 299464
rect 67548 298732 67600 298784
rect 167644 298732 167696 298784
rect 253112 298188 253164 298240
rect 262404 298188 262456 298240
rect 256608 298120 256660 298172
rect 285772 298120 285824 298172
rect 255872 297440 255924 297492
rect 266360 297440 266412 297492
rect 256516 297372 256568 297424
rect 259552 297372 259604 297424
rect 287244 297372 287296 297424
rect 119344 296692 119396 296744
rect 191748 296692 191800 296744
rect 259368 296624 259420 296676
rect 262496 296624 262548 296676
rect 76012 295944 76064 295996
rect 174636 295944 174688 295996
rect 256608 295944 256660 295996
rect 258264 295944 258316 295996
rect 276388 295944 276440 295996
rect 128360 295332 128412 295384
rect 187608 295332 187660 295384
rect 193036 295332 193088 295384
rect 256608 294992 256660 295044
rect 262496 294992 262548 295044
rect 96620 294584 96672 294636
rect 129096 294584 129148 294636
rect 140136 294584 140188 294636
rect 186964 294584 187016 294636
rect 258080 294584 258132 294636
rect 258264 294584 258316 294636
rect 184848 294108 184900 294160
rect 191748 294108 191800 294160
rect 102968 294040 103020 294092
rect 104164 294040 104216 294092
rect 256608 293972 256660 294024
rect 269120 293972 269172 294024
rect 102140 293904 102192 293956
rect 102784 293904 102836 293956
rect 128360 293904 128412 293956
rect 93124 293292 93176 293344
rect 102140 293292 102192 293344
rect 84200 293224 84252 293276
rect 177304 293224 177356 293276
rect 262404 293224 262456 293276
rect 281540 293224 281592 293276
rect 256608 292884 256660 292936
rect 259644 292884 259696 292936
rect 260748 292884 260800 292936
rect 99288 292476 99340 292528
rect 187424 292544 187476 292596
rect 191748 292544 191800 292596
rect 255412 292204 255464 292256
rect 259368 292204 259420 292256
rect 264888 291864 264940 291916
rect 280804 291864 280856 291916
rect 291200 291864 291252 291916
rect 53656 291796 53708 291848
rect 183468 291796 183520 291848
rect 191748 291796 191800 291848
rect 260748 291796 260800 291848
rect 291476 291796 291528 291848
rect 182916 291728 182968 291780
rect 72424 291184 72476 291236
rect 76012 291184 76064 291236
rect 98460 291184 98512 291236
rect 99288 291184 99340 291236
rect 255412 290504 255464 290556
rect 258448 290504 258500 290556
rect 262588 290504 262640 290556
rect 39856 290436 39908 290488
rect 61752 290436 61804 290488
rect 73252 290436 73304 290488
rect 77024 290436 77076 290488
rect 84844 290436 84896 290488
rect 88616 290436 88668 290488
rect 99564 290436 99616 290488
rect 258724 290436 258776 290488
rect 274824 290436 274876 290488
rect 184848 290300 184900 290352
rect 188896 290300 188948 290352
rect 191748 290300 191800 290352
rect 61844 290096 61896 290148
rect 62764 290096 62816 290148
rect 108396 289824 108448 289876
rect 184848 289824 184900 289876
rect 169760 289756 169812 289808
rect 171048 289756 171100 289808
rect 191564 289756 191616 289808
rect 255504 289756 255556 289808
rect 267832 289756 267884 289808
rect 274824 289756 274876 289808
rect 118976 289144 119028 289196
rect 151176 289144 151228 289196
rect 91008 289076 91060 289128
rect 185584 289076 185636 289128
rect 253664 288736 253716 288788
rect 254124 288736 254176 288788
rect 56324 288464 56376 288516
rect 72516 288464 72568 288516
rect 90272 288464 90324 288516
rect 91008 288464 91060 288516
rect 67364 288396 67416 288448
rect 118056 288396 118108 288448
rect 253848 288396 253900 288448
rect 269212 288396 269264 288448
rect 7564 288328 7616 288380
rect 37096 288328 37148 288380
rect 166540 288328 166592 288380
rect 166908 288328 166960 288380
rect 191748 288328 191800 288380
rect 255320 288328 255372 288380
rect 265256 288328 265308 288380
rect 171876 288260 171928 288312
rect 172428 288260 172480 288312
rect 190644 288260 190696 288312
rect 255504 288260 255556 288312
rect 261024 288260 261076 288312
rect 68652 287716 68704 287768
rect 78680 287716 78732 287768
rect 157984 287716 158036 287768
rect 166540 287716 166592 287768
rect 37096 287648 37148 287700
rect 70492 287648 70544 287700
rect 159364 287648 159416 287700
rect 171876 287648 171928 287700
rect 88064 287104 88116 287156
rect 93768 287104 93820 287156
rect 157984 287104 158036 287156
rect 75828 286968 75880 287020
rect 77944 286968 77996 287020
rect 79232 286968 79284 287020
rect 79968 286968 80020 287020
rect 159364 287036 159416 287088
rect 255504 286968 255556 287020
rect 276112 286968 276164 287020
rect 255412 286900 255464 286952
rect 262220 286900 262272 286952
rect 97448 286560 97500 286612
rect 97908 286560 97960 286612
rect 81992 286424 82044 286476
rect 83464 286424 83516 286476
rect 86868 286288 86920 286340
rect 88984 286288 89036 286340
rect 169760 286288 169812 286340
rect 170588 286288 170640 286340
rect 180156 286288 180208 286340
rect 50988 285744 51040 285796
rect 69112 285744 69164 285796
rect 69664 285744 69716 285796
rect 70308 285744 70360 285796
rect 76012 285744 76064 285796
rect 78588 285744 78640 285796
rect 45468 285540 45520 285592
rect 51724 285540 51776 285592
rect 73620 285676 73672 285728
rect 90824 285744 90876 285796
rect 112444 285744 112496 285796
rect 160928 285744 160980 285796
rect 191012 285744 191064 285796
rect 169760 285676 169812 285728
rect 48136 285472 48188 285524
rect 80152 285608 80204 285660
rect 177304 284928 177356 284980
rect 191748 284928 191800 284980
rect 96436 284384 96488 284436
rect 92388 284316 92440 284368
rect 99012 284316 99064 284368
rect 115848 284316 115900 284368
rect 176568 284316 176620 284368
rect 178040 284316 178092 284368
rect 263692 284316 263744 284368
rect 264888 284316 264940 284368
rect 152648 284248 152700 284300
rect 193036 284248 193088 284300
rect 255504 284248 255556 284300
rect 266452 284248 266504 284300
rect 267832 284248 267884 284300
rect 259092 284180 259144 284232
rect 266544 284180 266596 284232
rect 130568 283568 130620 283620
rect 152648 283568 152700 283620
rect 73252 283432 73304 283484
rect 74724 283364 74776 283416
rect 92480 283364 92532 283416
rect 92940 283364 92992 283416
rect 67548 283024 67600 283076
rect 99104 283228 99156 283280
rect 70952 283024 71004 283076
rect 98828 283024 98880 283076
rect 64696 282956 64748 283008
rect 66812 282956 66864 283008
rect 75368 282956 75420 283008
rect 81256 282956 81308 283008
rect 89536 282956 89588 283008
rect 65892 282208 65944 282260
rect 66168 282208 66220 282260
rect 57796 282140 57848 282192
rect 67088 282140 67140 282192
rect 67272 282140 67324 282192
rect 98000 282820 98052 282872
rect 168472 282820 168524 282872
rect 169576 282820 169628 282872
rect 191564 282820 191616 282872
rect 255504 282820 255556 282872
rect 268016 282820 268068 282872
rect 100760 282684 100812 282736
rect 102876 282684 102928 282736
rect 115848 282140 115900 282192
rect 149704 282140 149756 282192
rect 168472 282140 168524 282192
rect 255412 281868 255464 281920
rect 259460 281868 259512 281920
rect 98920 281596 98972 281648
rect 98000 281528 98052 281580
rect 173808 281528 173860 281580
rect 184296 281528 184348 281580
rect 191748 281528 191800 281580
rect 100760 281460 100812 281512
rect 118976 281460 119028 281512
rect 168288 281460 168340 281512
rect 171876 281460 171928 281512
rect 255412 281324 255464 281376
rect 259092 281324 259144 281376
rect 255412 281188 255464 281240
rect 259736 281188 259788 281240
rect 167736 280780 167788 280832
rect 175924 280780 175976 280832
rect 61752 280236 61804 280288
rect 66904 280236 66956 280288
rect 14464 280168 14516 280220
rect 66536 280168 66588 280220
rect 67180 280168 67232 280220
rect 100852 280168 100904 280220
rect 156696 280168 156748 280220
rect 100760 280100 100812 280152
rect 159548 280100 159600 280152
rect 168472 280100 168524 280152
rect 191564 280100 191616 280152
rect 255412 280100 255464 280152
rect 278964 280100 279016 280152
rect 255504 280032 255556 280084
rect 274732 280032 274784 280084
rect 4068 279420 4120 279472
rect 45376 279420 45428 279472
rect 60556 279420 60608 279472
rect 66628 279420 66680 279472
rect 98828 279420 98880 279472
rect 165528 279420 165580 279472
rect 189908 279420 189960 279472
rect 53564 278672 53616 278724
rect 53748 278672 53800 278724
rect 99104 278672 99156 278724
rect 157340 278672 157392 278724
rect 173808 278672 173860 278724
rect 174636 278672 174688 278724
rect 255412 278672 255464 278724
rect 261116 278672 261168 278724
rect 100760 278604 100812 278656
rect 130476 278604 130528 278656
rect 53564 277992 53616 278044
rect 66812 277992 66864 278044
rect 133236 277992 133288 278044
rect 174544 277992 174596 278044
rect 263692 277516 263744 277568
rect 269304 277516 269356 277568
rect 174636 277380 174688 277432
rect 192852 277380 192904 277432
rect 61660 277312 61712 277364
rect 66904 277312 66956 277364
rect 118056 277312 118108 277364
rect 100760 277244 100812 277296
rect 163504 277244 163556 277296
rect 185492 277312 185544 277364
rect 193220 277312 193272 277364
rect 255412 277312 255464 277364
rect 273536 277312 273588 277364
rect 190460 277244 190512 277296
rect 191288 277244 191340 277296
rect 255504 277244 255556 277296
rect 269396 277244 269448 277296
rect 269396 276020 269448 276072
rect 271880 276020 271932 276072
rect 99012 275952 99064 276004
rect 185584 275952 185636 276004
rect 255412 275952 255464 276004
rect 271972 275952 272024 276004
rect 108304 274660 108356 274712
rect 110420 274660 110472 274712
rect 255412 274660 255464 274712
rect 100760 274592 100812 274644
rect 177856 274592 177908 274644
rect 182180 274592 182232 274644
rect 255504 274592 255556 274644
rect 273444 274592 273496 274644
rect 183008 274524 183060 274576
rect 255412 274524 255464 274576
rect 265164 274524 265216 274576
rect 269304 274524 269356 274576
rect 273904 274524 273956 274576
rect 274640 274524 274692 274576
rect 53748 273912 53800 273964
rect 65892 273912 65944 273964
rect 66536 273912 66588 273964
rect 100760 273164 100812 273216
rect 108948 273164 109000 273216
rect 255504 273164 255556 273216
rect 281724 273164 281776 273216
rect 255412 273096 255464 273148
rect 259460 273096 259512 273148
rect 157340 272552 157392 272604
rect 172520 272552 172572 272604
rect 173808 272552 173860 272604
rect 50896 272484 50948 272536
rect 60464 272484 60516 272536
rect 108948 272484 109000 272536
rect 135996 272484 136048 272536
rect 162216 272484 162268 272536
rect 177304 272484 177356 272536
rect 177396 271940 177448 271992
rect 191748 271940 191800 271992
rect 43996 271872 44048 271924
rect 66628 271872 66680 271924
rect 173808 271872 173860 271924
rect 191656 271872 191708 271924
rect 100760 271804 100812 271856
rect 105636 271804 105688 271856
rect 164148 271804 164200 271856
rect 164884 271804 164936 271856
rect 184296 271804 184348 271856
rect 255412 271804 255464 271856
rect 270684 271804 270736 271856
rect 46848 271124 46900 271176
rect 60556 271124 60608 271176
rect 106188 271124 106240 271176
rect 115204 271124 115256 271176
rect 60556 270512 60608 270564
rect 66260 270512 66312 270564
rect 175924 270512 175976 270564
rect 191748 270512 191800 270564
rect 255412 270512 255464 270564
rect 258264 270512 258316 270564
rect 261024 270512 261076 270564
rect 59176 270444 59228 270496
rect 60648 270444 60700 270496
rect 100760 270444 100812 270496
rect 106096 270444 106148 270496
rect 255504 270444 255556 270496
rect 265072 270444 265124 270496
rect 291292 270444 291344 270496
rect 291660 270444 291712 270496
rect 580172 270444 580224 270496
rect 145656 269832 145708 269884
rect 162124 269832 162176 269884
rect 144828 269764 144880 269816
rect 188436 269764 188488 269816
rect 259368 269764 259420 269816
rect 277492 269764 277544 269816
rect 104256 269084 104308 269136
rect 123484 269084 123536 269136
rect 185768 269084 185820 269136
rect 190828 269084 190880 269136
rect 255412 269084 255464 269136
rect 57888 269016 57940 269068
rect 60648 269016 60700 269068
rect 100760 269016 100812 269068
rect 133236 269016 133288 269068
rect 258724 269016 258776 269068
rect 293960 269016 294012 269068
rect 255412 268948 255464 269000
rect 259368 268948 259420 269000
rect 255504 268880 255556 268932
rect 258816 268880 258868 268932
rect 60648 268404 60700 268456
rect 66904 268404 66956 268456
rect 54852 268336 54904 268388
rect 55036 268336 55088 268388
rect 66812 268336 66864 268388
rect 100760 268336 100812 268388
rect 111064 268336 111116 268388
rect 188436 267792 188488 267844
rect 191748 267792 191800 267844
rect 180156 267724 180208 267776
rect 191472 267724 191524 267776
rect 52368 266976 52420 267028
rect 63224 266976 63276 267028
rect 66628 266976 66680 267028
rect 100760 266976 100812 267028
rect 104808 266976 104860 267028
rect 156420 266976 156472 267028
rect 176016 266976 176068 267028
rect 255412 266976 255464 267028
rect 266820 266976 266872 267028
rect 267648 266976 267700 267028
rect 63316 266364 63368 266416
rect 66444 266364 66496 266416
rect 104808 266364 104860 266416
rect 109776 266364 109828 266416
rect 186964 266364 187016 266416
rect 191748 266364 191800 266416
rect 255504 266364 255556 266416
rect 260932 266364 260984 266416
rect 255412 266296 255464 266348
rect 291384 266296 291436 266348
rect 119436 265684 119488 265736
rect 144276 265684 144328 265736
rect 48044 265616 48096 265668
rect 57244 265616 57296 265668
rect 101496 265616 101548 265668
rect 151268 265616 151320 265668
rect 168288 265616 168340 265668
rect 184940 265616 184992 265668
rect 57244 264936 57296 264988
rect 57888 264936 57940 264988
rect 66812 264936 66864 264988
rect 100760 264936 100812 264988
rect 115204 264936 115256 264988
rect 184204 264936 184256 264988
rect 190828 264936 190880 264988
rect 255504 264936 255556 264988
rect 262496 264936 262548 264988
rect 39948 264188 40000 264240
rect 66260 264188 66312 264240
rect 255412 264188 255464 264240
rect 269856 264188 269908 264240
rect 100852 263644 100904 263696
rect 148508 263644 148560 263696
rect 173164 263644 173216 263696
rect 191748 263644 191800 263696
rect 59084 263576 59136 263628
rect 66812 263576 66864 263628
rect 100760 263576 100812 263628
rect 184296 263576 184348 263628
rect 255412 263576 255464 263628
rect 266544 263576 266596 263628
rect 267188 263576 267240 263628
rect 255044 263236 255096 263288
rect 259276 263236 259328 263288
rect 39304 262828 39356 262880
rect 67088 262828 67140 262880
rect 100760 262828 100812 262880
rect 108396 262828 108448 262880
rect 255596 262828 255648 262880
rect 265164 262828 265216 262880
rect 276020 262828 276072 262880
rect 169024 262284 169076 262336
rect 191012 262284 191064 262336
rect 100760 262216 100812 262268
rect 124864 262216 124916 262268
rect 163504 262216 163556 262268
rect 191748 262216 191800 262268
rect 278136 262216 278188 262268
rect 284392 262216 284444 262268
rect 100852 262148 100904 262200
rect 106188 262148 106240 262200
rect 126244 262148 126296 262200
rect 284668 262148 284720 262200
rect 288716 262148 288768 262200
rect 14556 260856 14608 260908
rect 66904 260856 66956 260908
rect 164884 260856 164936 260908
rect 191564 260856 191616 260908
rect 258816 260856 258868 260908
rect 284668 260856 284720 260908
rect 255412 260788 255464 260840
rect 280344 260788 280396 260840
rect 271788 260720 271840 260772
rect 289912 260720 289964 260772
rect 56508 260108 56560 260160
rect 66260 260108 66312 260160
rect 169116 259632 169168 259684
rect 170680 259632 170732 259684
rect 100760 259496 100812 259548
rect 133236 259496 133288 259548
rect 100852 259428 100904 259480
rect 145748 259428 145800 259480
rect 170404 259428 170456 259480
rect 191748 259428 191800 259480
rect 255504 259428 255556 259480
rect 270684 259428 270736 259480
rect 271788 259428 271840 259480
rect 255412 259360 255464 259412
rect 260748 259360 260800 259412
rect 278044 259360 278096 259412
rect 281632 259360 281684 259412
rect 580172 259360 580224 259412
rect 49608 258680 49660 258732
rect 64788 258680 64840 258732
rect 66444 258680 66496 258732
rect 101680 258680 101732 258732
rect 155408 258680 155460 258732
rect 167644 258136 167696 258188
rect 191748 258136 191800 258188
rect 126244 258068 126296 258120
rect 190644 258068 190696 258120
rect 258172 258068 258224 258120
rect 285956 258068 286008 258120
rect 287060 258068 287112 258120
rect 50712 258000 50764 258052
rect 66260 258000 66312 258052
rect 66444 258000 66496 258052
rect 68192 258000 68244 258052
rect 190736 258000 190788 258052
rect 193404 258000 193456 258052
rect 255412 257388 255464 257440
rect 258816 257388 258868 257440
rect 111156 257320 111208 257372
rect 171968 257320 172020 257372
rect 180616 257320 180668 257372
rect 183560 257320 183612 257372
rect 263784 257320 263836 257372
rect 285864 257320 285916 257372
rect 63408 256844 63460 256896
rect 66628 256844 66680 256896
rect 171784 256708 171836 256760
rect 191656 256708 191708 256760
rect 255412 256708 255464 256760
rect 261116 256708 261168 256760
rect 255504 256028 255556 256080
rect 263784 256028 263836 256080
rect 124128 255960 124180 256012
rect 159456 255960 159508 256012
rect 255412 255960 255464 256012
rect 287704 255960 287756 256012
rect 288624 255960 288676 256012
rect 100852 255348 100904 255400
rect 174820 255348 174872 255400
rect 177304 255348 177356 255400
rect 191012 255348 191064 255400
rect 174544 255280 174596 255332
rect 190828 255280 190880 255332
rect 3148 255212 3200 255264
rect 14464 255212 14516 255264
rect 255504 255212 255556 255264
rect 258172 255212 258224 255264
rect 100852 254940 100904 254992
rect 105544 254940 105596 254992
rect 53472 254532 53524 254584
rect 59268 254532 59320 254584
rect 66812 254532 66864 254584
rect 100852 253920 100904 253972
rect 153936 253920 153988 253972
rect 160744 253920 160796 253972
rect 191656 253920 191708 253972
rect 255412 253920 255464 253972
rect 266636 253920 266688 253972
rect 266912 253920 266964 253972
rect 270408 253852 270460 253904
rect 287152 253852 287204 253904
rect 255412 253240 255464 253292
rect 269396 253240 269448 253292
rect 270408 253240 270460 253292
rect 18604 253172 18656 253224
rect 66996 253172 67048 253224
rect 67272 253172 67324 253224
rect 108396 253172 108448 253224
rect 145656 253172 145708 253224
rect 161020 253172 161072 253224
rect 174728 253172 174780 253224
rect 258540 253172 258592 253224
rect 277584 253172 277636 253224
rect 278136 253172 278188 253224
rect 279424 253104 279476 253156
rect 281632 253104 281684 253156
rect 185676 252628 185728 252680
rect 191656 252628 191708 252680
rect 100852 252560 100904 252612
rect 105544 252560 105596 252612
rect 181444 252560 181496 252612
rect 191564 252560 191616 252612
rect 66904 252492 66956 252544
rect 68284 252492 68336 252544
rect 108488 252492 108540 252544
rect 108856 252492 108908 252544
rect 119344 252492 119396 252544
rect 176476 251880 176528 251932
rect 179420 251880 179472 251932
rect 54944 251812 54996 251864
rect 66812 251812 66864 251864
rect 106924 251812 106976 251864
rect 168380 251812 168432 251864
rect 177488 251812 177540 251864
rect 255412 251812 255464 251864
rect 258264 251812 258316 251864
rect 270408 251812 270460 251864
rect 582380 251812 582432 251864
rect 255504 251200 255556 251252
rect 269396 251200 269448 251252
rect 270408 251200 270460 251252
rect 53656 251132 53708 251184
rect 66812 251132 66864 251184
rect 107844 251132 107896 251184
rect 109684 251132 109736 251184
rect 160008 251132 160060 251184
rect 161112 251132 161164 251184
rect 100852 250996 100904 251048
rect 104256 250996 104308 251048
rect 101956 250452 102008 250504
rect 108488 250452 108540 250504
rect 262312 250452 262364 250504
rect 280252 250452 280304 250504
rect 255872 249908 255924 249960
rect 257344 249908 257396 249960
rect 41236 249772 41288 249824
rect 66444 249772 66496 249824
rect 112536 249772 112588 249824
rect 160008 249772 160060 249824
rect 160836 249772 160888 249824
rect 190644 249772 190696 249824
rect 255504 249772 255556 249824
rect 262312 249772 262364 249824
rect 99196 249704 99248 249756
rect 111800 249704 111852 249756
rect 254952 249704 255004 249756
rect 278044 249704 278096 249756
rect 55128 249024 55180 249076
rect 55864 249024 55916 249076
rect 66628 249024 66680 249076
rect 100852 249024 100904 249076
rect 103612 249024 103664 249076
rect 255412 249024 255464 249076
rect 269028 249024 269080 249076
rect 104808 248548 104860 248600
rect 106280 248548 106332 248600
rect 166264 248480 166316 248532
rect 190828 248480 190880 248532
rect 116676 248412 116728 248464
rect 192484 248412 192536 248464
rect 269028 248412 269080 248464
rect 582380 248412 582432 248464
rect 110972 247664 111024 247716
rect 115940 247664 115992 247716
rect 142988 247664 143040 247716
rect 189908 247664 189960 247716
rect 255504 247664 255556 247716
rect 262680 247664 262732 247716
rect 102784 247052 102836 247104
rect 110420 247052 110472 247104
rect 110972 247052 111024 247104
rect 183008 247052 183060 247104
rect 191656 247052 191708 247104
rect 252928 247052 252980 247104
rect 254032 247052 254084 247104
rect 254216 247052 254268 247104
rect 258172 247052 258224 247104
rect 100852 246304 100904 246356
rect 108304 246304 108356 246356
rect 184848 246304 184900 246356
rect 193680 246304 193732 246356
rect 255412 246304 255464 246356
rect 280160 246304 280212 246356
rect 255412 245760 255464 245812
rect 259644 245760 259696 245812
rect 100852 245624 100904 245676
rect 147128 245624 147180 245676
rect 58992 245556 59044 245608
rect 66812 245556 66864 245608
rect 255412 245556 255464 245608
rect 273352 245556 273404 245608
rect 100852 244944 100904 244996
rect 107752 244944 107804 244996
rect 151360 244944 151412 244996
rect 166356 244944 166408 244996
rect 184480 244944 184532 244996
rect 103612 244876 103664 244928
rect 129740 244876 129792 244928
rect 147036 244876 147088 244928
rect 192944 244876 192996 244928
rect 273352 244876 273404 244928
rect 291292 244876 291344 244928
rect 187148 244264 187200 244316
rect 191656 244264 191708 244316
rect 255504 244264 255556 244316
rect 273352 244264 273404 244316
rect 56416 244196 56468 244248
rect 66812 244196 66864 244248
rect 255412 244196 255464 244248
rect 281816 244196 281868 244248
rect 288624 244196 288676 244248
rect 98000 243516 98052 243568
rect 98276 243516 98328 243568
rect 140136 243516 140188 243568
rect 145748 243516 145800 243568
rect 184388 243516 184440 243568
rect 253204 243516 253256 243568
rect 262404 243516 262456 243568
rect 59268 242904 59320 242956
rect 66628 242904 66680 242956
rect 67640 242904 67692 242956
rect 68652 242904 68704 242956
rect 61752 242156 61804 242208
rect 100852 242904 100904 242956
rect 107016 242904 107068 242956
rect 178684 242904 178736 242956
rect 191656 242904 191708 242956
rect 75368 241748 75420 241800
rect 95976 241748 96028 241800
rect 82636 241612 82688 241664
rect 130568 241612 130620 241664
rect 93216 241544 93268 241596
rect 97724 241544 97776 241596
rect 102232 241544 102284 241596
rect 81440 241476 81492 241528
rect 82406 241476 82458 241528
rect 135996 241476 136048 241528
rect 214012 241476 214064 241528
rect 215208 241476 215260 241528
rect 257068 241544 257120 241596
rect 220084 241476 220136 241528
rect 249064 241476 249116 241528
rect 251916 241476 251968 241528
rect 252928 241476 252980 241528
rect 3516 241408 3568 241460
rect 14556 241408 14608 241460
rect 58532 241408 58584 241460
rect 58900 241408 58952 241460
rect 74678 241408 74730 241460
rect 151268 241408 151320 241460
rect 273444 241408 273496 241460
rect 273904 241408 273956 241460
rect 68928 241340 68980 241392
rect 77484 241340 77536 241392
rect 192944 241340 192996 241392
rect 205180 241340 205232 241392
rect 244280 240796 244332 240848
rect 255412 240796 255464 240848
rect 50896 240728 50948 240780
rect 58532 240728 58584 240780
rect 180248 240728 180300 240780
rect 186320 240728 186372 240780
rect 255596 240728 255648 240780
rect 582564 240728 582616 240780
rect 75920 240116 75972 240168
rect 76564 240116 76616 240168
rect 80060 240116 80112 240168
rect 80980 240116 81032 240168
rect 91100 240116 91152 240168
rect 92296 240116 92348 240168
rect 95240 240116 95292 240168
rect 95884 240116 95936 240168
rect 101404 240116 101456 240168
rect 172612 240116 172664 240168
rect 209044 240116 209096 240168
rect 69480 240048 69532 240100
rect 163596 240048 163648 240100
rect 164056 240048 164108 240100
rect 73896 239980 73948 240032
rect 164976 239980 165028 240032
rect 195244 240048 195296 240100
rect 251824 240048 251876 240100
rect 254032 240048 254084 240100
rect 256884 239980 256936 240032
rect 77484 239912 77536 239964
rect 77944 239912 77996 239964
rect 197360 239436 197412 239488
rect 231860 239436 231912 239488
rect 164056 239368 164108 239420
rect 171140 239368 171192 239420
rect 211896 239368 211948 239420
rect 256056 239232 256108 239284
rect 256792 239232 256844 239284
rect 284300 239368 284352 239420
rect 52368 238756 52420 238808
rect 69204 238756 69256 238808
rect 243544 238756 243596 238808
rect 248512 238756 248564 238808
rect 64604 238688 64656 238740
rect 77668 238688 77720 238740
rect 84292 238688 84344 238740
rect 111892 238688 111944 238740
rect 112536 238688 112588 238740
rect 82820 238620 82872 238672
rect 95148 238620 95200 238672
rect 125508 238076 125560 238128
rect 177396 238076 177448 238128
rect 246304 238076 246356 238128
rect 261116 238076 261168 238128
rect 174820 238008 174872 238060
rect 238852 238008 238904 238060
rect 248420 238008 248472 238060
rect 250352 238008 250404 238060
rect 270684 238008 270736 238060
rect 77668 237396 77720 237448
rect 78036 237396 78088 237448
rect 79968 237396 80020 237448
rect 80152 237396 80204 237448
rect 94688 237396 94740 237448
rect 95332 237396 95384 237448
rect 193220 237396 193272 237448
rect 195980 237396 196032 237448
rect 84200 237328 84252 237380
rect 180248 237328 180300 237380
rect 168288 237260 168340 237312
rect 262496 237260 262548 237312
rect 61844 236716 61896 236768
rect 73436 236716 73488 236768
rect 56324 236648 56376 236700
rect 74632 236648 74684 236700
rect 74816 236648 74868 236700
rect 84936 236648 84988 236700
rect 111064 236648 111116 236700
rect 126428 236648 126480 236700
rect 206284 236648 206336 236700
rect 209780 236648 209832 236700
rect 215944 236648 215996 236700
rect 265164 236648 265216 236700
rect 95148 235968 95200 236020
rect 98184 235968 98236 236020
rect 104624 235968 104676 236020
rect 104992 235968 105044 236020
rect 200764 235968 200816 236020
rect 201868 235968 201920 236020
rect 193680 235764 193732 235816
rect 194784 235764 194836 235816
rect 197360 235764 197412 235816
rect 245568 235288 245620 235340
rect 253204 235288 253256 235340
rect 3516 235220 3568 235272
rect 39304 235220 39356 235272
rect 91192 235220 91244 235272
rect 116584 235220 116636 235272
rect 124220 235220 124272 235272
rect 160008 235220 160060 235272
rect 195152 235220 195204 235272
rect 205180 235220 205232 235272
rect 219440 235220 219492 235272
rect 252468 235220 252520 235272
rect 272064 235220 272116 235272
rect 96528 234608 96580 234660
rect 100852 234608 100904 234660
rect 67456 234540 67508 234592
rect 111156 234540 111208 234592
rect 159548 234540 159600 234592
rect 268016 234540 268068 234592
rect 195152 234472 195204 234524
rect 209044 234472 209096 234524
rect 228364 233860 228416 233912
rect 255320 233860 255372 233912
rect 94780 233656 94832 233708
rect 101404 233656 101456 233708
rect 71780 233180 71832 233232
rect 73068 233180 73120 233232
rect 151360 233180 151412 233232
rect 176476 233180 176528 233232
rect 269396 233180 269448 233232
rect 76012 233112 76064 233164
rect 76564 233112 76616 233164
rect 116676 233112 116728 233164
rect 156696 233112 156748 233164
rect 230480 233112 230532 233164
rect 231768 233112 231820 233164
rect 176016 232976 176068 233028
rect 176476 232976 176528 233028
rect 254584 232500 254636 232552
rect 580172 232500 580224 232552
rect 97264 231752 97316 231804
rect 97908 231752 97960 231804
rect 184388 231752 184440 231804
rect 261024 231752 261076 231804
rect 68284 231072 68336 231124
rect 77484 231072 77536 231124
rect 240232 231072 240284 231124
rect 278964 231072 279016 231124
rect 18604 230528 18656 230580
rect 97264 230528 97316 230580
rect 77484 230460 77536 230512
rect 182180 230460 182232 230512
rect 182916 230460 182968 230512
rect 67272 230392 67324 230444
rect 108396 230392 108448 230444
rect 133236 230392 133288 230444
rect 277400 230392 277452 230444
rect 89720 229712 89772 229764
rect 111064 229712 111116 229764
rect 118700 229712 118752 229764
rect 218704 229712 218756 229764
rect 222200 229712 222252 229764
rect 253204 229712 253256 229764
rect 260840 229712 260892 229764
rect 112444 229032 112496 229084
rect 215300 229032 215352 229084
rect 215300 228692 215352 228744
rect 215944 228692 215996 228744
rect 80060 228352 80112 228404
rect 111800 228352 111852 228404
rect 119436 228352 119488 228404
rect 149888 228352 149940 228404
rect 238852 228352 238904 228404
rect 240048 228352 240100 228404
rect 262864 228352 262916 228404
rect 270776 228352 270828 228404
rect 3424 227672 3476 227724
rect 92480 227672 92532 227724
rect 148508 227060 148560 227112
rect 237380 227060 237432 227112
rect 258816 227060 258868 227112
rect 274824 227060 274876 227112
rect 65800 226992 65852 227044
rect 260932 226992 260984 227044
rect 92480 226312 92532 226364
rect 93124 226312 93176 226364
rect 236092 225632 236144 225684
rect 283012 225632 283064 225684
rect 65984 225564 66036 225616
rect 169116 225564 169168 225616
rect 213184 225564 213236 225616
rect 263876 225564 263928 225616
rect 580264 225564 580316 225616
rect 170772 224272 170824 224324
rect 53564 224204 53616 224256
rect 177396 224204 177448 224256
rect 240784 224272 240836 224324
rect 258172 224272 258224 224324
rect 213920 224204 213972 224256
rect 265624 224204 265676 224256
rect 88340 223524 88392 223576
rect 121460 223524 121512 223576
rect 152556 222912 152608 222964
rect 220820 222912 220872 222964
rect 222108 222912 222160 222964
rect 63224 222844 63276 222896
rect 159456 222844 159508 222896
rect 163688 222844 163740 222896
rect 237380 222844 237432 222896
rect 67364 222096 67416 222148
rect 269304 222096 269356 222148
rect 222844 221416 222896 221468
rect 254124 221416 254176 221468
rect 171048 220804 171100 220856
rect 173348 220804 173400 220856
rect 113824 220736 113876 220788
rect 236092 220736 236144 220788
rect 100116 220056 100168 220108
rect 277492 220056 277544 220108
rect 277676 220056 277728 220108
rect 288440 219376 288492 219428
rect 579896 219376 579948 219428
rect 77944 218764 77996 218816
rect 87604 218764 87656 218816
rect 103428 218764 103480 218816
rect 184204 218764 184256 218816
rect 60648 218696 60700 218748
rect 156696 218696 156748 218748
rect 254584 218696 254636 218748
rect 104256 217948 104308 218000
rect 240784 217948 240836 218000
rect 158628 217880 158680 217932
rect 272156 217880 272208 217932
rect 48136 217268 48188 217320
rect 77300 217268 77352 217320
rect 88248 217268 88300 217320
rect 154488 217268 154540 217320
rect 118608 215976 118660 216028
rect 185768 215976 185820 216028
rect 187056 215976 187108 216028
rect 251824 215976 251876 216028
rect 177396 215908 177448 215960
rect 250444 215908 250496 215960
rect 259644 215908 259696 215960
rect 91100 215228 91152 215280
rect 170496 215228 170548 215280
rect 227720 215228 227772 215280
rect 227720 214752 227772 214804
rect 228456 214752 228508 214804
rect 100208 214548 100260 214600
rect 267832 214548 267884 214600
rect 98092 213868 98144 213920
rect 98736 213868 98788 213920
rect 93860 213256 93912 213308
rect 121552 213256 121604 213308
rect 98736 213188 98788 213240
rect 206376 213188 206428 213240
rect 121552 212508 121604 212560
rect 259552 212508 259604 212560
rect 254584 211760 254636 211812
rect 267924 211760 267976 211812
rect 96620 211080 96672 211132
rect 102324 211080 102376 211132
rect 154488 211080 154540 211132
rect 224960 211080 225012 211132
rect 53564 210400 53616 210452
rect 73252 210400 73304 210452
rect 88248 210400 88300 210452
rect 102140 210400 102192 210452
rect 102324 209788 102376 209840
rect 270592 209788 270644 209840
rect 102232 209720 102284 209772
rect 263692 209720 263744 209772
rect 88156 209040 88208 209092
rect 120080 209040 120132 209092
rect 224224 209040 224276 209092
rect 253940 209040 253992 209092
rect 98644 208360 98696 208412
rect 102232 208360 102284 208412
rect 175188 208360 175240 208412
rect 180064 208360 180116 208412
rect 86960 207680 87012 207732
rect 110512 207680 110564 207732
rect 97264 207612 97316 207664
rect 266452 207612 266504 207664
rect 110512 207000 110564 207052
rect 256700 207000 256752 207052
rect 79968 206252 80020 206304
rect 91100 206252 91152 206304
rect 93124 206252 93176 206304
rect 274640 206252 274692 206304
rect 91100 205640 91152 205692
rect 92388 205640 92440 205692
rect 176016 205640 176068 205692
rect 95240 204892 95292 204944
rect 95884 204892 95936 204944
rect 262220 204892 262272 204944
rect 262588 204892 262640 204944
rect 3424 204212 3476 204264
rect 7564 204212 7616 204264
rect 158076 204212 158128 204264
rect 271972 204212 272024 204264
rect 169116 203532 169168 203584
rect 178868 203532 178920 203584
rect 99380 202784 99432 202836
rect 100208 202784 100260 202836
rect 147128 202784 147180 202836
rect 241520 202784 241572 202836
rect 3240 202104 3292 202156
rect 99380 202104 99432 202156
rect 188344 201424 188396 201476
rect 188896 201424 188948 201476
rect 257344 201424 257396 201476
rect 192944 199384 192996 199436
rect 249064 199384 249116 199436
rect 117964 197276 118016 197328
rect 223580 197276 223632 197328
rect 223580 196664 223632 196716
rect 224224 196664 224276 196716
rect 20628 196596 20680 196648
rect 120724 196596 120776 196648
rect 233884 196596 233936 196648
rect 244372 196596 244424 196648
rect 108304 195916 108356 195968
rect 220912 195916 220964 195968
rect 221832 195916 221884 195968
rect 84936 195236 84988 195288
rect 106280 195236 106332 195288
rect 240784 194556 240836 194608
rect 580172 194556 580224 194608
rect 44088 193808 44140 193860
rect 149796 193808 149848 193860
rect 188988 193808 189040 193860
rect 574744 193808 574796 193860
rect 84844 192516 84896 192568
rect 115388 192516 115440 192568
rect 3884 192448 3936 192500
rect 133144 192448 133196 192500
rect 229836 192448 229888 192500
rect 266544 192448 266596 192500
rect 221832 191768 221884 191820
rect 225144 191768 225196 191820
rect 59268 191088 59320 191140
rect 173256 191088 173308 191140
rect 190368 191088 190420 191140
rect 263784 191088 263836 191140
rect 3424 188980 3476 189032
rect 18604 188980 18656 189032
rect 27528 188300 27580 188352
rect 148416 188300 148468 188352
rect 193772 188300 193824 188352
rect 236000 188300 236052 188352
rect 87604 187008 87656 187060
rect 104164 187008 104216 187060
rect 5448 186940 5500 186992
rect 155316 186940 155368 186992
rect 184296 186940 184348 186992
rect 200764 186940 200816 186992
rect 240784 186940 240836 186992
rect 276296 186940 276348 186992
rect 17224 185580 17276 185632
rect 144184 185580 144236 185632
rect 213184 185580 213236 185632
rect 235264 185580 235316 185632
rect 86868 184220 86920 184272
rect 97356 184220 97408 184272
rect 28908 184152 28960 184204
rect 189724 184152 189776 184204
rect 88984 182792 89036 182844
rect 120172 182792 120224 182844
rect 133144 181432 133196 181484
rect 206284 181432 206336 181484
rect 91008 180072 91060 180124
rect 117320 180072 117372 180124
rect 99196 179392 99248 179444
rect 226432 179392 226484 179444
rect 92296 178644 92348 178696
rect 118700 178644 118752 178696
rect 238024 178644 238076 178696
rect 238668 178644 238720 178696
rect 580172 178644 580224 178696
rect 71044 178032 71096 178084
rect 159548 178032 159600 178084
rect 75368 177352 75420 177404
rect 129004 177352 129056 177404
rect 198004 177352 198056 177404
rect 226708 177352 226760 177404
rect 80796 177284 80848 177336
rect 106464 177284 106516 177336
rect 219532 177284 219584 177336
rect 219716 177284 219768 177336
rect 154028 175312 154080 175364
rect 204260 175312 204312 175364
rect 204904 175312 204956 175364
rect 89720 175244 89772 175296
rect 219440 175244 219492 175296
rect 220084 175244 220136 175296
rect 85580 174496 85632 174548
rect 195980 174496 196032 174548
rect 215944 174496 215996 174548
rect 153936 173884 153988 173936
rect 222200 173884 222252 173936
rect 222936 173884 222988 173936
rect 80704 173136 80756 173188
rect 160928 173136 160980 173188
rect 195244 173136 195296 173188
rect 206376 173136 206428 173188
rect 227812 173136 227864 173188
rect 75920 171776 75972 171828
rect 156604 171776 156656 171828
rect 202880 171776 202932 171828
rect 104624 171096 104676 171148
rect 210424 171096 210476 171148
rect 211160 171096 211212 171148
rect 317420 171096 317472 171148
rect 189724 170348 189776 170400
rect 250444 170348 250496 170400
rect 582748 170348 582800 170400
rect 67824 169736 67876 169788
rect 68560 169736 68612 169788
rect 194508 169736 194560 169788
rect 81532 168988 81584 169040
rect 154028 168988 154080 169040
rect 154488 168988 154540 169040
rect 162308 168988 162360 169040
rect 204996 168988 205048 169040
rect 193864 168376 193916 168428
rect 194508 168376 194560 168428
rect 166448 168308 166500 168360
rect 211160 168308 211212 168360
rect 234528 168308 234580 168360
rect 243544 168308 243596 168360
rect 82912 167628 82964 167680
rect 166448 167628 166500 167680
rect 141608 167016 141660 167068
rect 223580 167016 223632 167068
rect 200120 166336 200172 166388
rect 229836 166336 229888 166388
rect 84200 166268 84252 166320
rect 157984 166268 158036 166320
rect 213184 166268 213236 166320
rect 218060 166268 218112 166320
rect 267740 166268 267792 166320
rect 54944 165588 54996 165640
rect 190460 165588 190512 165640
rect 191196 165588 191248 165640
rect 92664 164840 92716 164892
rect 153936 164840 153988 164892
rect 202880 164296 202932 164348
rect 300124 164296 300176 164348
rect 100208 164228 100260 164280
rect 100668 164228 100720 164280
rect 237472 164228 237524 164280
rect 77392 163548 77444 163600
rect 154488 163548 154540 163600
rect 91744 163480 91796 163532
rect 129096 163480 129148 163532
rect 221004 163480 221056 163532
rect 3424 162868 3476 162920
rect 51816 162868 51868 162920
rect 153936 162868 153988 162920
rect 218060 162868 218112 162920
rect 84108 162120 84160 162172
rect 109040 162120 109092 162172
rect 243544 162120 243596 162172
rect 274640 162120 274692 162172
rect 148416 161508 148468 161560
rect 199384 161508 199436 161560
rect 233240 161508 233292 161560
rect 129188 161440 129240 161492
rect 241704 161440 241756 161492
rect 193036 160760 193088 160812
rect 245200 160760 245252 160812
rect 213276 160692 213328 160744
rect 277584 160692 277636 160744
rect 176568 160148 176620 160200
rect 196716 160148 196768 160200
rect 87604 160080 87656 160132
rect 88248 160080 88300 160132
rect 182088 160080 182140 160132
rect 72976 159332 73028 159384
rect 176568 159332 176620 159384
rect 229836 159332 229888 159384
rect 287704 159332 287756 159384
rect 194600 158788 194652 158840
rect 195244 158788 195296 158840
rect 250444 158788 250496 158840
rect 93860 158720 93912 158772
rect 95148 158720 95200 158772
rect 223672 158720 223724 158772
rect 210424 158652 210476 158704
rect 291292 158652 291344 158704
rect 45376 157972 45428 158024
rect 63500 157972 63552 158024
rect 186228 157972 186280 158024
rect 208400 157972 208452 158024
rect 291292 157972 291344 158024
rect 582932 157972 582984 158024
rect 209780 157428 209832 157480
rect 210424 157428 210476 157480
rect 63500 157360 63552 157412
rect 64604 157360 64656 157412
rect 189908 157360 189960 157412
rect 202144 157360 202196 157412
rect 202788 157360 202840 157412
rect 230572 157360 230624 157412
rect 206284 156680 206336 156732
rect 252468 156680 252520 156732
rect 255964 156680 256016 156732
rect 220820 156612 220872 156664
rect 582656 156612 582708 156664
rect 57704 156000 57756 156052
rect 162216 156000 162268 156052
rect 71780 155932 71832 155984
rect 72884 155932 72936 155984
rect 197452 155932 197504 155984
rect 70584 155252 70636 155304
rect 74632 155252 74684 155304
rect 183008 155252 183060 155304
rect 43996 155184 44048 155236
rect 178776 155184 178828 155236
rect 212724 154504 212776 154556
rect 213184 154504 213236 154556
rect 88340 153892 88392 153944
rect 153936 153892 153988 153944
rect 57888 153824 57940 153876
rect 187056 153824 187108 153876
rect 187148 153280 187200 153332
rect 224408 153280 224460 153332
rect 212724 153212 212776 153264
rect 295340 153212 295392 153264
rect 215392 153144 215444 153196
rect 259460 153144 259512 153196
rect 182088 152532 182140 152584
rect 216680 152532 216732 152584
rect 54852 152464 54904 152516
rect 184296 152464 184348 152516
rect 184204 151784 184256 151836
rect 202052 151784 202104 151836
rect 180248 150492 180300 150544
rect 214012 150492 214064 150544
rect 215484 150492 215536 150544
rect 215944 150492 215996 150544
rect 251180 150492 251232 150544
rect 127624 150424 127676 150476
rect 220912 150424 220964 150476
rect 208492 150356 208544 150408
rect 209136 150356 209188 150408
rect 281724 150356 281776 150408
rect 89628 149744 89680 149796
rect 127624 149744 127676 149796
rect 67732 149676 67784 149728
rect 77484 149676 77536 149728
rect 124864 149676 124916 149728
rect 240140 149676 240192 149728
rect 240784 149676 240836 149728
rect 77576 149132 77628 149184
rect 80796 149132 80848 149184
rect 86316 149132 86368 149184
rect 88984 149132 89036 149184
rect 67548 149064 67600 149116
rect 105636 149064 105688 149116
rect 212448 148996 212500 149048
rect 271880 148996 271932 149048
rect 183008 148384 183060 148436
rect 196072 148384 196124 148436
rect 162216 148316 162268 148368
rect 211804 148316 211856 148368
rect 61936 147704 61988 147756
rect 127624 147704 127676 147756
rect 76196 147636 76248 147688
rect 159456 147636 159508 147688
rect 205180 147636 205232 147688
rect 260104 147636 260156 147688
rect 194600 146956 194652 147008
rect 195060 146956 195112 147008
rect 200212 146956 200264 147008
rect 200948 146956 201000 147008
rect 223672 146956 223724 147008
rect 224592 146956 224644 147008
rect 60464 146888 60516 146940
rect 161020 146888 161072 146940
rect 214012 146888 214064 146940
rect 225052 146888 225104 146940
rect 226524 146888 226576 146940
rect 264980 146888 265032 146940
rect 165528 146344 165580 146396
rect 193772 146344 193824 146396
rect 98828 146276 98880 146328
rect 99288 146276 99340 146328
rect 230664 146276 230716 146328
rect 196716 146208 196768 146260
rect 199200 146208 199252 146260
rect 191656 145868 191708 145920
rect 193864 145868 193916 145920
rect 3332 145528 3384 145580
rect 95700 145528 95752 145580
rect 180156 145528 180208 145580
rect 188344 145528 188396 145580
rect 234528 145528 234580 145580
rect 340144 145528 340196 145580
rect 63132 144984 63184 145036
rect 63316 144984 63368 145036
rect 138756 144984 138808 145036
rect 206468 144984 206520 145036
rect 235264 144984 235316 145036
rect 95424 144916 95476 144968
rect 95700 144916 95752 144968
rect 226524 144916 226576 144968
rect 51816 144848 51868 144900
rect 87604 144848 87656 144900
rect 97448 144848 97500 144900
rect 100208 144848 100260 144900
rect 73804 144168 73856 144220
rect 165528 144168 165580 144220
rect 186872 143624 186924 143676
rect 225604 143624 225656 143676
rect 156604 143556 156656 143608
rect 211252 143556 211304 143608
rect 220084 143556 220136 143608
rect 246304 143556 246356 143608
rect 219532 143080 219584 143132
rect 220728 143080 220780 143132
rect 218244 142944 218296 142996
rect 218704 142944 218756 142996
rect 92572 142808 92624 142860
rect 149704 142808 149756 142860
rect 221924 142808 221976 142860
rect 60556 142196 60608 142248
rect 93216 142196 93268 142248
rect 223212 142196 223264 142248
rect 238024 142196 238076 142248
rect 46204 142128 46256 142180
rect 88708 142128 88760 142180
rect 204904 142128 204956 142180
rect 209780 142128 209832 142180
rect 218244 142128 218296 142180
rect 280896 142128 280948 142180
rect 63316 141516 63368 141568
rect 76564 141516 76616 141568
rect 76196 141448 76248 141500
rect 159364 141448 159416 141500
rect 203156 141448 203208 141500
rect 39856 141380 39908 141432
rect 72332 141380 72384 141432
rect 75828 141380 75880 141432
rect 170588 141380 170640 141432
rect 202604 141380 202656 141432
rect 219440 141380 219492 141432
rect 258724 141380 258776 141432
rect 203432 140768 203484 140820
rect 289084 140768 289136 140820
rect 188988 140428 189040 140480
rect 194784 140428 194836 140480
rect 64788 140020 64840 140072
rect 76656 140020 76708 140072
rect 85948 140020 86000 140072
rect 174636 140020 174688 140072
rect 59084 139408 59136 139460
rect 104256 139408 104308 139460
rect 174636 139408 174688 139460
rect 214656 140564 214708 140616
rect 213736 140496 213788 140548
rect 214840 140428 214892 140480
rect 224500 140428 224552 140480
rect 227904 140428 227956 140480
rect 249064 139408 249116 139460
rect 316040 138728 316092 138780
rect 51724 138660 51776 138712
rect 71228 138660 71280 138712
rect 88524 138660 88576 138712
rect 185584 138660 185636 138712
rect 226616 138660 226668 138712
rect 230480 138660 230532 138712
rect 582564 138660 582616 138712
rect 77392 138048 77444 138100
rect 77944 138048 77996 138100
rect 82912 138048 82964 138100
rect 83556 138048 83608 138100
rect 89720 138048 89772 138100
rect 90180 138048 90232 138100
rect 92388 138048 92440 138100
rect 92572 138048 92624 138100
rect 64512 137980 64564 138032
rect 81440 137980 81492 138032
rect 3240 137912 3292 137964
rect 72976 137912 73028 137964
rect 190092 137776 190144 137828
rect 192576 137776 192628 137828
rect 97356 137300 97408 137352
rect 100852 137300 100904 137352
rect 88708 137232 88760 137284
rect 96804 137232 96856 137284
rect 169208 137232 169260 137284
rect 187148 137232 187200 137284
rect 226616 137232 226668 137284
rect 233240 137232 233292 137284
rect 233884 137232 233936 137284
rect 72976 136688 73028 136740
rect 73160 136688 73212 136740
rect 74448 136688 74500 136740
rect 75184 136688 75236 136740
rect 81072 136688 81124 136740
rect 83464 136688 83516 136740
rect 85212 136688 85264 136740
rect 86316 136688 86368 136740
rect 66076 136620 66128 136672
rect 141700 136620 141752 136672
rect 88340 136552 88392 136604
rect 89628 136552 89680 136604
rect 91192 136552 91244 136604
rect 171876 136552 171928 136604
rect 191656 136552 191708 136604
rect 88616 136008 88668 136060
rect 89260 136008 89312 136060
rect 93768 135940 93820 135992
rect 141608 135940 141660 135992
rect 3424 135872 3476 135924
rect 88340 135872 88392 135924
rect 94228 135872 94280 135924
rect 151268 135872 151320 135924
rect 159364 135872 159416 135924
rect 169116 135872 169168 135924
rect 67272 135260 67324 135312
rect 94872 135260 94924 135312
rect 180156 135260 180208 135312
rect 191656 135260 191708 135312
rect 226800 135192 226852 135244
rect 278780 135192 278832 135244
rect 280068 135192 280120 135244
rect 69572 134988 69624 135040
rect 73804 134988 73856 135040
rect 68652 134784 68704 134836
rect 69664 134784 69716 134836
rect 93216 134580 93268 134632
rect 147128 134580 147180 134632
rect 94872 134512 94924 134564
rect 174636 134512 174688 134564
rect 280068 134512 280120 134564
rect 307024 134512 307076 134564
rect 173808 133832 173860 133884
rect 192484 133832 192536 133884
rect 226616 133696 226668 133748
rect 229192 133696 229244 133748
rect 96620 133152 96672 133204
rect 184388 133152 184440 133204
rect 225604 133152 225656 133204
rect 273444 133152 273496 133204
rect 50988 132404 51040 132456
rect 66260 132404 66312 132456
rect 138756 132404 138808 132456
rect 190460 132404 190512 132456
rect 191104 132404 191156 132456
rect 235264 132404 235316 132456
rect 280804 132404 280856 132456
rect 64696 132336 64748 132388
rect 66352 132336 66404 132388
rect 96712 132336 96764 132388
rect 148416 132336 148468 132388
rect 226340 132336 226392 132388
rect 238852 132336 238904 132388
rect 280804 131724 280856 131776
rect 305644 131724 305696 131776
rect 57796 131044 57848 131096
rect 66260 131044 66312 131096
rect 156696 131044 156748 131096
rect 190828 131044 190880 131096
rect 226340 131044 226392 131096
rect 266360 131044 266412 131096
rect 96620 130568 96672 130620
rect 102784 130568 102836 130620
rect 107016 130432 107068 130484
rect 152556 130432 152608 130484
rect 96712 130364 96764 130416
rect 188436 130364 188488 130416
rect 96712 129684 96764 129736
rect 181536 129684 181588 129736
rect 227076 129684 227128 129736
rect 227904 129684 227956 129736
rect 276388 129684 276440 129736
rect 278044 129684 278096 129736
rect 102784 129004 102836 129056
rect 156604 129004 156656 129056
rect 225328 128868 225380 128920
rect 228456 128868 228508 128920
rect 61660 128664 61712 128716
rect 66260 128664 66312 128716
rect 189080 128664 189132 128716
rect 191656 128664 191708 128716
rect 64604 128256 64656 128308
rect 66904 128256 66956 128308
rect 97632 128256 97684 128308
rect 147036 128256 147088 128308
rect 226800 128256 226852 128308
rect 237380 128256 237432 128308
rect 237380 127576 237432 127628
rect 331864 127576 331916 127628
rect 181536 126964 181588 127016
rect 191656 126964 191708 127016
rect 54944 126896 54996 126948
rect 66904 126896 66956 126948
rect 97908 126896 97960 126948
rect 152648 126896 152700 126948
rect 226616 126896 226668 126948
rect 229100 126896 229152 126948
rect 281632 126896 281684 126948
rect 61844 126828 61896 126880
rect 66812 126828 66864 126880
rect 226524 126828 226576 126880
rect 241704 126828 241756 126880
rect 287336 126828 287388 126880
rect 288348 126828 288400 126880
rect 176016 126216 176068 126268
rect 185584 126216 185636 126268
rect 288348 126216 288400 126268
rect 353300 126216 353352 126268
rect 97816 125536 97868 125588
rect 180248 125536 180300 125588
rect 190092 125740 190144 125792
rect 191012 125740 191064 125792
rect 190092 125604 190144 125656
rect 193128 125604 193180 125656
rect 97908 125468 97960 125520
rect 144184 125468 144236 125520
rect 147128 125468 147180 125520
rect 226800 125536 226852 125588
rect 231952 125536 232004 125588
rect 276204 125536 276256 125588
rect 63224 125332 63276 125384
rect 66812 125332 66864 125384
rect 53472 124856 53524 124908
rect 66812 124856 66864 124908
rect 246488 124856 246540 124908
rect 298100 124856 298152 124908
rect 97908 124108 97960 124160
rect 169208 124108 169260 124160
rect 226616 124108 226668 124160
rect 231860 124108 231912 124160
rect 280160 124108 280212 124160
rect 582840 124108 582892 124160
rect 110972 123428 111024 123480
rect 126336 123428 126388 123480
rect 141700 123428 141752 123480
rect 180616 123428 180668 123480
rect 189080 123428 189132 123480
rect 182364 122816 182416 122868
rect 193036 122816 193088 122868
rect 57704 122748 57756 122800
rect 66352 122748 66404 122800
rect 97908 122748 97960 122800
rect 129096 122748 129148 122800
rect 162308 122748 162360 122800
rect 181536 122748 181588 122800
rect 226616 122748 226668 122800
rect 237656 122748 237708 122800
rect 97448 122680 97500 122732
rect 124956 122680 125008 122732
rect 238116 122136 238168 122188
rect 246396 122136 246448 122188
rect 228456 122068 228508 122120
rect 267924 122068 267976 122120
rect 181628 121932 181680 121984
rect 187148 121932 187200 121984
rect 184296 121592 184348 121644
rect 184848 121592 184900 121644
rect 191564 121592 191616 121644
rect 43996 121388 44048 121440
rect 66812 121388 66864 121440
rect 97540 121388 97592 121440
rect 110972 121388 111024 121440
rect 178776 121388 178828 121440
rect 190092 121388 190144 121440
rect 226616 121388 226668 121440
rect 237564 121388 237616 121440
rect 60556 121320 60608 121372
rect 66904 121320 66956 121372
rect 97632 121048 97684 121100
rect 102784 121048 102836 121100
rect 104256 120708 104308 120760
rect 178040 120708 178092 120760
rect 233884 120708 233936 120760
rect 282184 120708 282236 120760
rect 187700 120096 187752 120148
rect 190828 120096 190880 120148
rect 60464 120028 60516 120080
rect 66812 120028 66864 120080
rect 97172 120028 97224 120080
rect 109684 120028 109736 120080
rect 160928 120028 160980 120080
rect 59176 119960 59228 120012
rect 66904 119960 66956 120012
rect 187056 120028 187108 120080
rect 191564 120028 191616 120080
rect 189724 119960 189776 120012
rect 226616 119620 226668 119672
rect 230572 119620 230624 119672
rect 229836 119348 229888 119400
rect 313280 119348 313332 119400
rect 54852 118600 54904 118652
rect 66812 118600 66864 118652
rect 97816 118600 97868 118652
rect 155316 118600 155368 118652
rect 184848 118600 184900 118652
rect 186964 118600 187016 118652
rect 56416 118532 56468 118584
rect 66904 118532 66956 118584
rect 97908 118532 97960 118584
rect 107016 118532 107068 118584
rect 226800 117988 226852 118040
rect 236000 117988 236052 118040
rect 178040 117920 178092 117972
rect 179328 117920 179380 117972
rect 190828 117920 190880 117972
rect 226616 117920 226668 117972
rect 240140 117920 240192 117972
rect 240784 117920 240836 117972
rect 186320 117308 186372 117360
rect 191564 117308 191616 117360
rect 63132 117240 63184 117292
rect 66628 117240 66680 117292
rect 97908 117240 97960 117292
rect 149796 117240 149848 117292
rect 159456 117240 159508 117292
rect 187700 117240 187752 117292
rect 182916 117172 182968 117224
rect 191380 117172 191432 117224
rect 226984 116628 227036 116680
rect 238760 116628 238812 116680
rect 231768 116560 231820 116612
rect 261024 116560 261076 116612
rect 188436 116016 188488 116068
rect 191564 116016 191616 116068
rect 226616 115948 226668 116000
rect 230480 115948 230532 116000
rect 231768 115948 231820 116000
rect 57888 115880 57940 115932
rect 66812 115880 66864 115932
rect 97540 115880 97592 115932
rect 124864 115880 124916 115932
rect 127624 115880 127676 115932
rect 170128 115880 170180 115932
rect 97172 115676 97224 115728
rect 100760 115676 100812 115728
rect 61936 115404 61988 115456
rect 66904 115404 66956 115456
rect 187608 115404 187660 115456
rect 191012 115404 191064 115456
rect 227996 115268 228048 115320
rect 277400 115268 277452 115320
rect 170128 115200 170180 115252
rect 171048 115200 171100 115252
rect 184848 115200 184900 115252
rect 186320 115200 186372 115252
rect 236000 115200 236052 115252
rect 304264 115200 304316 115252
rect 59084 114452 59136 114504
rect 66812 114452 66864 114504
rect 178868 114452 178920 114504
rect 191564 114452 191616 114504
rect 184480 114112 184532 114164
rect 186228 114112 186280 114164
rect 226524 113840 226576 113892
rect 230664 113840 230716 113892
rect 7564 113772 7616 113824
rect 63224 113772 63276 113824
rect 66904 113772 66956 113824
rect 244924 113772 244976 113824
rect 254584 113772 254636 113824
rect 97540 113160 97592 113212
rect 178776 113160 178828 113212
rect 186228 113160 186280 113212
rect 190828 113160 190880 113212
rect 227812 113160 227864 113212
rect 229836 113160 229888 113212
rect 157984 113092 158036 113144
rect 191564 113092 191616 113144
rect 226616 113092 226668 113144
rect 277492 113092 277544 113144
rect 278688 113092 278740 113144
rect 50804 112412 50856 112464
rect 67180 112412 67232 112464
rect 278688 112412 278740 112464
rect 324320 112412 324372 112464
rect 96712 111868 96764 111920
rect 98736 111868 98788 111920
rect 97908 111800 97960 111852
rect 184296 111800 184348 111852
rect 56508 111732 56560 111784
rect 66904 111732 66956 111784
rect 96712 111732 96764 111784
rect 98828 111732 98880 111784
rect 118700 111732 118752 111784
rect 167736 111732 167788 111784
rect 177396 111732 177448 111784
rect 191196 111732 191248 111784
rect 226708 111732 226760 111784
rect 244372 111732 244424 111784
rect 98736 111120 98788 111172
rect 118700 111120 118752 111172
rect 101404 111052 101456 111104
rect 188436 111052 188488 111104
rect 244372 111052 244424 111104
rect 291844 111052 291896 111104
rect 64512 110372 64564 110424
rect 66812 110372 66864 110424
rect 97908 110372 97960 110424
rect 184204 110372 184256 110424
rect 105636 110304 105688 110356
rect 191012 110304 191064 110356
rect 97080 110236 97132 110288
rect 100116 110236 100168 110288
rect 226984 109692 227036 109744
rect 263692 109692 263744 109744
rect 65524 109012 65576 109064
rect 65984 109012 66036 109064
rect 115388 108944 115440 108996
rect 164148 108944 164200 108996
rect 226616 108944 226668 108996
rect 229744 108944 229796 108996
rect 155316 108876 155368 108928
rect 158628 108876 158680 108928
rect 190276 108876 190328 108928
rect 164148 108264 164200 108316
rect 177396 108264 177448 108316
rect 236736 108264 236788 108316
rect 259552 108264 259604 108316
rect 240048 108128 240100 108180
rect 241520 108128 241572 108180
rect 98000 108060 98052 108112
rect 98920 108060 98972 108112
rect 98920 107652 98972 107704
rect 152556 107652 152608 107704
rect 166908 107584 166960 107636
rect 190644 107584 190696 107636
rect 226708 107584 226760 107636
rect 288532 107584 288584 107636
rect 289728 107584 289780 107636
rect 100116 106904 100168 106956
rect 110512 106904 110564 106956
rect 289728 106904 289780 106956
rect 342904 106904 342956 106956
rect 97908 106360 97960 106412
rect 157984 106360 158036 106412
rect 7564 106292 7616 106344
rect 66812 106292 66864 106344
rect 123576 106292 123628 106344
rect 185768 106292 185820 106344
rect 96804 106224 96856 106276
rect 100024 106224 100076 106276
rect 174636 106224 174688 106276
rect 191012 106224 191064 106276
rect 46848 105544 46900 105596
rect 66076 105544 66128 105596
rect 66628 105544 66680 105596
rect 98000 105544 98052 105596
rect 123576 105544 123628 105596
rect 271788 105544 271840 105596
rect 291476 105544 291528 105596
rect 188896 104864 188948 104916
rect 191564 104864 191616 104916
rect 226708 104864 226760 104916
rect 271788 104864 271840 104916
rect 53656 104796 53708 104848
rect 66812 104796 66864 104848
rect 227444 104116 227496 104168
rect 267832 104116 267884 104168
rect 102048 103504 102100 103556
rect 174636 103504 174688 103556
rect 187056 103504 187108 103556
rect 193220 103504 193272 103556
rect 226524 103504 226576 103556
rect 231860 103504 231912 103556
rect 323584 103504 323636 103556
rect 63408 103436 63460 103488
rect 67824 103436 67876 103488
rect 97908 103436 97960 103488
rect 129740 103436 129792 103488
rect 97816 103368 97868 103420
rect 102048 103368 102100 103420
rect 55036 102756 55088 102808
rect 61752 102756 61804 102808
rect 66812 102756 66864 102808
rect 129740 102756 129792 102808
rect 187240 102756 187292 102808
rect 227904 102756 227956 102808
rect 258816 102756 258868 102808
rect 278044 102756 278096 102808
rect 299480 102756 299532 102808
rect 188988 102212 189040 102264
rect 191472 102212 191524 102264
rect 188528 102144 188580 102196
rect 191564 102144 191616 102196
rect 226616 102144 226668 102196
rect 96712 102076 96764 102128
rect 98920 102076 98972 102128
rect 106280 102076 106332 102128
rect 169668 102076 169720 102128
rect 229744 102076 229796 102128
rect 287060 102076 287112 102128
rect 288348 102076 288400 102128
rect 96712 101804 96764 101856
rect 99380 101804 99432 101856
rect 41236 101396 41288 101448
rect 65984 101396 66036 101448
rect 66536 101396 66588 101448
rect 101496 101396 101548 101448
rect 106280 101396 106332 101448
rect 169668 101396 169720 101448
rect 182916 101396 182968 101448
rect 288348 101396 288400 101448
rect 321652 101396 321704 101448
rect 61844 100716 61896 100768
rect 66812 100716 66864 100768
rect 98828 100716 98880 100768
rect 190644 100716 190696 100768
rect 188344 100648 188396 100700
rect 191748 100648 191800 100700
rect 230388 99968 230440 100020
rect 240048 99968 240100 100020
rect 320824 99968 320876 100020
rect 185676 99560 185728 99612
rect 191564 99560 191616 99612
rect 55864 99424 55916 99476
rect 64604 99424 64656 99476
rect 66720 99424 66772 99476
rect 225144 99424 225196 99476
rect 242808 99424 242860 99476
rect 97908 99356 97960 99408
rect 185860 99356 185912 99408
rect 226432 99356 226484 99408
rect 229100 99356 229152 99408
rect 230388 99356 230440 99408
rect 97908 99016 97960 99068
rect 100760 99016 100812 99068
rect 97908 98132 97960 98184
rect 188436 98132 188488 98184
rect 101588 98064 101640 98116
rect 171048 98064 171100 98116
rect 187700 97996 187752 98048
rect 191748 97996 191800 98048
rect 226708 97996 226760 98048
rect 250536 97996 250588 98048
rect 3424 97928 3476 97980
rect 46204 97928 46256 97980
rect 187148 97928 187200 97980
rect 190644 97928 190696 97980
rect 253204 97928 253256 97980
rect 100024 97248 100076 97300
rect 187700 97248 187752 97300
rect 96712 96840 96764 96892
rect 98644 96840 98696 96892
rect 226340 96568 226392 96620
rect 240876 96568 240928 96620
rect 226892 95888 226944 95940
rect 266452 95888 266504 95940
rect 97816 95276 97868 95328
rect 187608 95276 187660 95328
rect 64696 95208 64748 95260
rect 66904 95208 66956 95260
rect 97908 95208 97960 95260
rect 190460 95208 190512 95260
rect 59268 95140 59320 95192
rect 66812 95140 66864 95192
rect 94872 94460 94924 94512
rect 117320 94460 117372 94512
rect 193404 94460 193456 94512
rect 242808 94460 242860 94512
rect 277400 94460 277452 94512
rect 97908 93644 97960 93696
rect 102324 93644 102376 93696
rect 94688 93508 94740 93560
rect 95884 93508 95936 93560
rect 171048 93168 171100 93220
rect 191748 93168 191800 93220
rect 193772 93168 193824 93220
rect 95148 93100 95200 93152
rect 120172 93100 120224 93152
rect 184388 93100 184440 93152
rect 185860 93100 185912 93152
rect 205088 93100 205140 93152
rect 67548 92828 67600 92880
rect 68376 92828 68428 92880
rect 68928 92692 68980 92744
rect 70262 92692 70314 92744
rect 88662 92692 88714 92744
rect 95240 92760 95292 92812
rect 81624 92556 81676 92608
rect 82590 92556 82642 92608
rect 89904 92556 89956 92608
rect 90686 92556 90738 92608
rect 62028 92488 62080 92540
rect 67548 92488 67600 92540
rect 222844 92488 222896 92540
rect 225236 92488 225288 92540
rect 52368 92420 52420 92472
rect 74724 92420 74776 92472
rect 95148 92420 95200 92472
rect 190460 92420 190512 92472
rect 226800 92420 226852 92472
rect 64788 92352 64840 92404
rect 76288 92352 76340 92404
rect 85580 92352 85632 92404
rect 88156 92352 88208 92404
rect 94872 92352 94924 92404
rect 179420 92352 179472 92404
rect 180708 92352 180760 92404
rect 210424 92352 210476 92404
rect 211068 92352 211120 92404
rect 95148 91060 95200 91112
rect 120080 91060 120132 91112
rect 220728 91060 220780 91112
rect 224960 91060 225012 91112
rect 84660 90992 84712 91044
rect 100852 90992 100904 91044
rect 212172 90992 212224 91044
rect 213276 90992 213328 91044
rect 228364 90992 228416 91044
rect 63316 90924 63368 90976
rect 78956 90924 79008 90976
rect 110420 90924 110472 90976
rect 75736 90856 75788 90908
rect 223764 90788 223816 90840
rect 224868 90788 224920 90840
rect 222476 90244 222528 90296
rect 226340 90244 226392 90296
rect 69204 89700 69256 89752
rect 71044 89700 71096 89752
rect 73068 89700 73120 89752
rect 74264 89700 74316 89752
rect 110420 89700 110472 89752
rect 111156 89700 111208 89752
rect 111248 89700 111300 89752
rect 111800 89700 111852 89752
rect 214656 89700 214708 89752
rect 218796 89700 218848 89752
rect 53564 89632 53616 89684
rect 73160 89632 73212 89684
rect 73712 89632 73764 89684
rect 89260 89632 89312 89684
rect 111064 89632 111116 89684
rect 217692 89632 217744 89684
rect 221372 89632 221424 89684
rect 236736 89632 236788 89684
rect 88708 89564 88760 89616
rect 89536 89564 89588 89616
rect 114376 89564 114428 89616
rect 204996 89564 205048 89616
rect 205088 89564 205140 89616
rect 229100 89564 229152 89616
rect 73160 89020 73212 89072
rect 77944 89020 77996 89072
rect 67456 88952 67508 89004
rect 87604 88952 87656 89004
rect 194692 88544 194744 88596
rect 194692 88340 194744 88392
rect 63224 88272 63276 88324
rect 101404 88272 101456 88324
rect 120080 88272 120132 88324
rect 214012 88272 214064 88324
rect 72332 88204 72384 88256
rect 96988 88204 97040 88256
rect 203708 88204 203760 88256
rect 204996 88204 205048 88256
rect 206284 88204 206336 88256
rect 207388 88204 207440 88256
rect 226800 87592 226852 87644
rect 241520 87592 241572 87644
rect 80980 86912 81032 86964
rect 115388 86912 115440 86964
rect 89812 86844 89864 86896
rect 116584 86844 116636 86896
rect 218244 86912 218296 86964
rect 185768 86844 185820 86896
rect 225052 86844 225104 86896
rect 3148 85484 3200 85536
rect 65524 85484 65576 85536
rect 87236 85484 87288 85536
rect 121460 85484 121512 85536
rect 215300 85484 215352 85536
rect 217324 85484 217376 85536
rect 244280 85484 244332 85536
rect 75460 85416 75512 85468
rect 101496 85416 101548 85468
rect 193220 85416 193272 85468
rect 216036 85416 216088 85468
rect 244280 84804 244332 84856
rect 245568 84804 245620 84856
rect 256056 84804 256108 84856
rect 71044 84124 71096 84176
rect 101588 84124 101640 84176
rect 80060 84056 80112 84108
rect 107660 84124 107712 84176
rect 205640 84124 205692 84176
rect 206928 84124 206980 84176
rect 191656 83512 191708 83564
rect 267004 83512 267056 83564
rect 210424 83444 210476 83496
rect 582840 83444 582892 83496
rect 65984 82764 66036 82816
rect 155500 82764 155552 82816
rect 187240 82764 187292 82816
rect 229744 82764 229796 82816
rect 76012 82696 76064 82748
rect 104164 82696 104216 82748
rect 200396 82084 200448 82136
rect 245660 82084 245712 82136
rect 281540 82084 281592 82136
rect 322940 82084 322992 82136
rect 65524 81404 65576 81456
rect 65984 81404 66036 81456
rect 87604 81336 87656 81388
rect 189908 81336 189960 81388
rect 80152 81268 80204 81320
rect 111248 81268 111300 81320
rect 167736 81268 167788 81320
rect 214564 81268 214616 81320
rect 198740 80044 198792 80096
rect 244280 80044 244332 80096
rect 67732 79976 67784 80028
rect 184204 79976 184256 80028
rect 184480 79976 184532 80028
rect 81716 79908 81768 79960
rect 115296 79908 115348 79960
rect 177396 79908 177448 79960
rect 207020 79908 207072 79960
rect 207020 79500 207072 79552
rect 207664 79500 207716 79552
rect 190368 79296 190420 79348
rect 284300 79296 284352 79348
rect 97448 78616 97500 78668
rect 225144 78616 225196 78668
rect 97356 78548 97408 78600
rect 222844 78548 222896 78600
rect 81624 77188 81676 77240
rect 109040 77188 109092 77240
rect 209780 77188 209832 77240
rect 206928 77120 206980 77172
rect 262864 77120 262916 77172
rect 71688 76508 71740 76560
rect 171784 76508 171836 76560
rect 77944 75828 77996 75880
rect 198740 75828 198792 75880
rect 152556 75760 152608 75812
rect 227904 75828 227956 75880
rect 228364 75828 228416 75880
rect 84200 74468 84252 74520
rect 115940 74468 115992 74520
rect 212540 74468 212592 74520
rect 215944 73788 215996 73840
rect 248420 73788 248472 73840
rect 69848 73108 69900 73160
rect 196164 73108 196216 73160
rect 212540 73108 212592 73160
rect 282920 73108 282972 73160
rect 174636 73040 174688 73092
rect 231860 73040 231912 73092
rect 282920 72428 282972 72480
rect 333980 72428 334032 72480
rect 67824 71680 67876 71732
rect 187700 71680 187752 71732
rect 196624 71680 196676 71732
rect 244924 71680 244976 71732
rect 195980 71340 196032 71392
rect 196624 71340 196676 71392
rect 89628 71000 89680 71052
rect 163504 71000 163556 71052
rect 69204 70320 69256 70372
rect 194692 70320 194744 70372
rect 194692 69912 194744 69964
rect 195336 69912 195388 69964
rect 216036 69640 216088 69692
rect 266360 69640 266412 69692
rect 64696 68960 64748 69012
rect 192576 68960 192628 69012
rect 193036 68960 193088 69012
rect 188436 68892 188488 68944
rect 250536 68892 250588 68944
rect 86868 68280 86920 68332
rect 164884 68280 164936 68332
rect 193128 68280 193180 68332
rect 309140 68280 309192 68332
rect 61844 67532 61896 67584
rect 191104 67532 191156 67584
rect 196164 67532 196216 67584
rect 285772 67532 285824 67584
rect 94504 67464 94556 67516
rect 222200 67464 222252 67516
rect 222844 67464 222896 67516
rect 285772 66852 285824 66904
rect 320180 66852 320232 66904
rect 86960 66172 87012 66224
rect 219716 66172 219768 66224
rect 220084 66172 220136 66224
rect 66168 66104 66220 66156
rect 185676 66104 185728 66156
rect 93768 64812 93820 64864
rect 226340 64812 226392 64864
rect 68284 64744 68336 64796
rect 193864 64744 193916 64796
rect 195336 64744 195388 64796
rect 289820 64744 289872 64796
rect 289820 64132 289872 64184
rect 345020 64132 345072 64184
rect 226340 63520 226392 63572
rect 226984 63520 227036 63572
rect 142988 62772 143040 62824
rect 180156 62772 180208 62824
rect 192484 62772 192536 62824
rect 242992 62772 243044 62824
rect 89536 62024 89588 62076
rect 217324 62024 217376 62076
rect 73344 60664 73396 60716
rect 199384 60664 199436 60716
rect 66904 59984 66956 60036
rect 131764 59984 131816 60036
rect 286416 59984 286468 60036
rect 292672 59984 292724 60036
rect 2964 59304 3016 59356
rect 57244 59304 57296 59356
rect 101404 59304 101456 59356
rect 200120 59304 200172 59356
rect 201408 59304 201460 59356
rect 57888 58624 57940 58676
rect 181444 58624 181496 58676
rect 187056 58624 187108 58676
rect 269120 58624 269172 58676
rect 68928 57876 68980 57928
rect 195244 57876 195296 57928
rect 111064 57808 111116 57860
rect 206284 57808 206336 57860
rect 206928 57196 206980 57248
rect 213184 57196 213236 57248
rect 213276 57196 213328 57248
rect 280804 57196 280856 57248
rect 70400 56516 70452 56568
rect 196624 56516 196676 56568
rect 201408 56516 201460 56568
rect 273260 56516 273312 56568
rect 273260 55836 273312 55888
rect 340972 55836 341024 55888
rect 73068 53048 73120 53100
rect 138664 53048 138716 53100
rect 189724 53048 189776 53100
rect 270500 53048 270552 53100
rect 101404 51688 101456 51740
rect 134616 51688 134668 51740
rect 207664 51688 207716 51740
rect 274640 51688 274692 51740
rect 185584 50328 185636 50380
rect 248420 50328 248472 50380
rect 53656 47540 53708 47592
rect 146944 47540 146996 47592
rect 183008 47540 183060 47592
rect 338120 47540 338172 47592
rect 188344 46860 188396 46912
rect 580172 46860 580224 46912
rect 115848 46248 115900 46300
rect 142896 46248 142948 46300
rect 59268 46180 59320 46232
rect 135904 46180 135956 46232
rect 3424 45500 3476 45552
rect 65524 45500 65576 45552
rect 66168 44820 66220 44872
rect 140044 44820 140096 44872
rect 184204 44820 184256 44872
rect 253204 44820 253256 44872
rect 62028 43392 62080 43444
rect 137376 43392 137428 43444
rect 251824 43392 251876 43444
rect 349804 43392 349856 43444
rect 79968 42032 80020 42084
rect 151176 42032 151228 42084
rect 199384 42032 199436 42084
rect 233884 42032 233936 42084
rect 236644 42032 236696 42084
rect 289820 42032 289872 42084
rect 77208 40672 77260 40724
rect 142804 40672 142856 40724
rect 186964 40672 187016 40724
rect 249800 40672 249852 40724
rect 250444 40672 250496 40724
rect 285680 40672 285732 40724
rect 119896 39312 119948 39364
rect 151084 39312 151136 39364
rect 179328 39312 179380 39364
rect 305736 39312 305788 39364
rect 55036 37884 55088 37936
rect 145564 37884 145616 37936
rect 180616 37884 180668 37936
rect 332692 37884 332744 37936
rect 111708 36524 111760 36576
rect 141516 36524 141568 36576
rect 193864 36524 193916 36576
rect 291200 36524 291252 36576
rect 61660 35164 61712 35216
rect 125600 35164 125652 35216
rect 204904 35164 204956 35216
rect 340236 35164 340288 35216
rect 108948 33736 109000 33788
rect 155224 33736 155276 33788
rect 280896 33736 280948 33788
rect 325700 33736 325752 33788
rect 3516 33056 3568 33108
rect 58624 33056 58676 33108
rect 70216 32376 70268 32428
rect 133144 32376 133196 32428
rect 46848 31016 46900 31068
rect 160836 31016 160888 31068
rect 197360 31016 197412 31068
rect 342260 31016 342312 31068
rect 43996 29588 44048 29640
rect 166264 29588 166316 29640
rect 209688 29588 209740 29640
rect 278780 29588 278832 29640
rect 121368 28228 121420 28280
rect 175924 28228 175976 28280
rect 192576 28228 192628 28280
rect 328460 28228 328512 28280
rect 61936 26868 61988 26920
rect 160744 26868 160796 26920
rect 229836 26868 229888 26920
rect 260840 26868 260892 26920
rect 100668 25508 100720 25560
rect 162124 25508 162176 25560
rect 204168 25508 204220 25560
rect 324412 25508 324464 25560
rect 84016 24080 84068 24132
rect 152464 24080 152516 24132
rect 206284 24080 206336 24132
rect 247040 24080 247092 24132
rect 250536 24080 250588 24132
rect 331220 24080 331272 24132
rect 102048 22720 102100 22772
rect 141424 22720 141476 22772
rect 214564 22720 214616 22772
rect 347044 22720 347096 22772
rect 86776 21360 86828 21412
rect 137284 21360 137336 21412
rect 191748 21360 191800 21412
rect 264980 21360 265032 21412
rect 3424 20612 3476 20664
rect 93124 20612 93176 20664
rect 93768 19932 93820 19984
rect 169024 19932 169076 19984
rect 220084 19932 220136 19984
rect 284392 19932 284444 19984
rect 95056 18572 95108 18624
rect 130384 18572 130436 18624
rect 253296 18572 253348 18624
rect 344284 18572 344336 18624
rect 99288 17280 99340 17332
rect 215944 17280 215996 17332
rect 240784 17280 240836 17332
rect 256700 17280 256752 17332
rect 78588 17212 78640 17264
rect 126244 17212 126296 17264
rect 202788 17212 202840 17264
rect 321560 17212 321612 17264
rect 68928 15852 68980 15904
rect 174544 15852 174596 15904
rect 184848 15852 184900 15904
rect 280712 15852 280764 15904
rect 226984 14424 227036 14476
rect 303160 14424 303212 14476
rect 64788 13064 64840 13116
rect 177304 13064 177356 13116
rect 181536 13064 181588 13116
rect 281540 13064 281592 13116
rect 251180 11772 251232 11824
rect 252376 11772 252428 11824
rect 90916 11704 90968 11756
rect 153844 11704 153896 11756
rect 195244 11704 195296 11756
rect 312176 11704 312228 11756
rect 332692 11704 332744 11756
rect 333888 11704 333940 11756
rect 97908 10344 97960 10396
rect 148324 10344 148376 10396
rect 2688 10276 2740 10328
rect 101404 10276 101456 10328
rect 222844 10276 222896 10328
rect 334716 10276 334768 10328
rect 271788 9596 271840 9648
rect 276020 9596 276072 9648
rect 255964 8984 256016 9036
rect 302424 8984 302476 9036
rect 82084 8916 82136 8968
rect 170404 8916 170456 8968
rect 196624 8916 196676 8968
rect 258264 8916 258316 8968
rect 100300 7556 100352 7608
rect 159364 7556 159416 7608
rect 3424 6604 3476 6656
rect 7564 6604 7616 6656
rect 251180 6196 251232 6248
rect 263600 6196 263652 6248
rect 224868 6128 224920 6180
rect 254676 6128 254728 6180
rect 256056 6128 256108 6180
rect 292488 6128 292540 6180
rect 300124 5584 300176 5636
rect 306748 5584 306800 5636
rect 305736 5516 305788 5568
rect 309048 5516 309100 5568
rect 349804 5516 349856 5568
rect 351644 5516 351696 5568
rect 96252 4836 96304 4888
rect 173164 4836 173216 4888
rect 228364 4836 228416 4888
rect 239312 4836 239364 4888
rect 572 4768 624 4820
rect 97264 4768 97316 4820
rect 238024 4768 238076 4820
rect 270040 4768 270092 4820
rect 323584 4768 323636 4820
rect 330392 4768 330444 4820
rect 331864 4496 331916 4548
rect 337476 4496 337528 4548
rect 291844 4428 291896 4480
rect 297272 4428 297324 4480
rect 134524 4156 134576 4208
rect 136456 4156 136508 4208
rect 307024 4156 307076 4208
rect 315028 4156 315080 4208
rect 342996 4088 343048 4140
rect 346952 4088 347004 4140
rect 233884 4020 233936 4072
rect 240508 4020 240560 4072
rect 8760 3544 8812 3596
rect 22744 3544 22796 3596
rect 66720 3544 66772 3596
rect 76564 3544 76616 3596
rect 85672 3544 85724 3596
rect 86776 3544 86828 3596
rect 1676 3476 1728 3528
rect 2688 3476 2740 3528
rect 2872 3476 2924 3528
rect 3976 3476 4028 3528
rect 9956 3476 10008 3528
rect 10968 3476 11020 3528
rect 11152 3476 11204 3528
rect 12348 3476 12400 3528
rect 15936 3476 15988 3528
rect 16488 3476 16540 3528
rect 17040 3476 17092 3528
rect 17868 3476 17920 3528
rect 18236 3476 18288 3528
rect 19248 3476 19300 3528
rect 24216 3476 24268 3528
rect 24768 3476 24820 3528
rect 26516 3476 26568 3528
rect 27528 3476 27580 3528
rect 32404 3476 32456 3528
rect 33048 3476 33100 3528
rect 33600 3476 33652 3528
rect 34428 3476 34480 3528
rect 34796 3476 34848 3528
rect 35808 3476 35860 3528
rect 35992 3476 36044 3528
rect 37096 3476 37148 3528
rect 40684 3476 40736 3528
rect 41144 3476 41196 3528
rect 41880 3476 41932 3528
rect 42708 3476 42760 3528
rect 43076 3476 43128 3528
rect 43996 3476 44048 3528
rect 48964 3476 49016 3528
rect 49608 3476 49660 3528
rect 50160 3476 50212 3528
rect 50712 3476 50764 3528
rect 52552 3476 52604 3528
rect 53656 3476 53708 3528
rect 57244 3476 57296 3528
rect 57888 3476 57940 3528
rect 58440 3476 58492 3528
rect 59268 3476 59320 3528
rect 59636 3476 59688 3528
rect 60648 3476 60700 3528
rect 60832 3476 60884 3528
rect 61936 3476 61988 3528
rect 64328 3476 64380 3528
rect 64788 3476 64840 3528
rect 65524 3476 65576 3528
rect 66168 3476 66220 3528
rect 67916 3476 67968 3528
rect 68928 3476 68980 3528
rect 69112 3476 69164 3528
rect 70216 3476 70268 3528
rect 72608 3476 72660 3528
rect 73068 3476 73120 3528
rect 75000 3476 75052 3528
rect 75828 3476 75880 3528
rect 76196 3476 76248 3528
rect 77208 3476 77260 3528
rect 80888 3476 80940 3528
rect 81348 3476 81400 3528
rect 89168 3476 89220 3528
rect 89628 3476 89680 3528
rect 90364 3476 90416 3528
rect 90916 3476 90968 3528
rect 91008 3476 91060 3528
rect 91560 3476 91612 3528
rect 92756 3476 92808 3528
rect 93768 3476 93820 3528
rect 93952 3476 94004 3528
rect 95056 3476 95108 3528
rect 97448 3476 97500 3528
rect 97908 3476 97960 3528
rect 98644 3476 98696 3528
rect 99288 3476 99340 3528
rect 99840 3476 99892 3528
rect 100668 3476 100720 3528
rect 101036 3476 101088 3528
rect 102048 3476 102100 3528
rect 102232 3476 102284 3528
rect 106832 3476 106884 3528
rect 106924 3476 106976 3528
rect 107568 3476 107620 3528
rect 108120 3476 108172 3528
rect 108948 3476 109000 3528
rect 109316 3476 109368 3528
rect 110328 3476 110380 3528
rect 114008 3476 114060 3528
rect 114468 3476 114520 3528
rect 115204 3476 115256 3528
rect 115848 3476 115900 3528
rect 116400 3476 116452 3528
rect 117228 3476 117280 3528
rect 117596 3476 117648 3528
rect 118608 3476 118660 3528
rect 122288 3476 122340 3528
rect 122748 3476 122800 3528
rect 123484 3476 123536 3528
rect 124128 3476 124180 3528
rect 124680 3476 124732 3528
rect 125508 3476 125560 3528
rect 143540 3476 143592 3528
rect 144828 3476 144880 3528
rect 147128 3476 147180 3528
rect 147588 3476 147640 3528
rect 249064 3476 249116 3528
rect 255872 3476 255924 3528
rect 260104 3476 260156 3528
rect 267740 3476 267792 3528
rect 280804 3476 280856 3528
rect 287796 3476 287848 3528
rect 299480 3476 299532 3528
rect 300768 3476 300820 3528
rect 302424 3476 302476 3528
rect 305552 3476 305604 3528
rect 324320 3476 324372 3528
rect 325608 3476 325660 3528
rect 340144 3476 340196 3528
rect 342168 3476 342220 3528
rect 1308 3408 1360 3460
rect 13544 3408 13596 3460
rect 32312 3408 32364 3460
rect 51356 3408 51408 3460
rect 66904 3408 66956 3460
rect 83280 3408 83332 3460
rect 84016 3408 84068 3460
rect 12348 3340 12400 3392
rect 27712 3340 27764 3392
rect 33784 3340 33836 3392
rect 77392 3340 77444 3392
rect 98552 3408 98604 3460
rect 105728 3408 105780 3460
rect 115112 3408 115164 3460
rect 213184 3408 213236 3460
rect 242900 3408 242952 3460
rect 246304 3408 246356 3460
rect 253480 3408 253532 3460
rect 267004 3408 267056 3460
rect 273628 3408 273680 3460
rect 320824 3408 320876 3460
rect 332692 3408 332744 3460
rect 334716 3408 334768 3460
rect 339868 3408 339920 3460
rect 344284 3408 344336 3460
rect 350448 3408 350500 3460
rect 574744 3408 574796 3460
rect 582196 3408 582248 3460
rect 253204 3340 253256 3392
rect 264152 3340 264204 3392
rect 309876 3340 309928 3392
rect 311440 3340 311492 3392
rect 289084 3272 289136 3324
rect 292580 3272 292632 3324
rect 340236 3272 340288 3324
rect 344560 3272 344612 3324
rect 317328 3204 317380 3256
rect 321652 3204 321704 3256
rect 581000 3204 581052 3256
rect 582472 3204 582524 3256
rect 25320 3136 25372 3188
rect 26148 3136 26200 3188
rect 118792 3068 118844 3120
rect 119804 3068 119856 3120
rect 299664 3068 299716 3120
rect 302240 3068 302292 3120
rect 347044 3068 347096 3120
rect 349252 3068 349304 3120
rect 55128 3000 55180 3052
rect 56048 3000 56100 3052
rect 258724 3000 258776 3052
rect 260656 3000 260708 3052
rect 304264 3000 304316 3052
rect 307944 3000 307996 3052
rect 282184 2932 282236 2984
rect 283104 2932 283156 2984
rect 292488 2932 292540 2984
rect 294880 2932 294932 2984
rect 270040 2796 270092 2848
rect 272432 2796 272484 2848
rect 140044 2728 140096 2780
rect 142988 2728 143040 2780
rect 7656 2048 7708 2100
rect 17224 2048 17276 2100
rect 19432 2048 19484 2100
rect 178684 2048 178736 2100
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 104912 703582 105308 703610
rect 8128 702710 8156 703520
rect 24320 702914 24348 703520
rect 24308 702908 24360 702914
rect 24308 702850 24360 702856
rect 40512 702778 40540 703520
rect 72988 703050 73016 703520
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 70308 702840 70360 702846
rect 70308 702782 70360 702788
rect 40500 702772 40552 702778
rect 40500 702714 40552 702720
rect 8116 702704 8168 702710
rect 8116 702646 8168 702652
rect 66168 702568 66220 702574
rect 66168 702510 66220 702516
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683194 3464 684247
rect 3424 683188 3476 683194
rect 3424 683130 3476 683136
rect 39304 683188 39356 683194
rect 39304 683130 39356 683136
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 14464 670744 14516 670750
rect 14464 670686 14516 670692
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 656946 3464 658135
rect 3424 656940 3476 656946
rect 3424 656882 3476 656888
rect 3422 632088 3478 632097
rect 3422 632023 3478 632032
rect 2778 606112 2834 606121
rect 2778 606047 2834 606056
rect 2792 605946 2820 606047
rect 2780 605940 2832 605946
rect 2780 605882 2832 605888
rect 3436 576842 3464 632023
rect 3514 619168 3570 619177
rect 3514 619103 3570 619112
rect 3528 618322 3556 619103
rect 3516 618316 3568 618322
rect 3516 618258 3568 618264
rect 11704 618316 11756 618322
rect 11704 618258 11756 618264
rect 4804 605940 4856 605946
rect 4804 605882 4856 605888
rect 4816 587178 4844 605882
rect 4804 587172 4856 587178
rect 4804 587114 4856 587120
rect 8114 581088 8170 581097
rect 8114 581023 8170 581032
rect 8128 580242 8156 581023
rect 3516 580236 3568 580242
rect 3516 580178 3568 580184
rect 8116 580236 8168 580242
rect 8116 580178 8168 580184
rect 3528 580009 3556 580178
rect 3514 580000 3570 580009
rect 3514 579935 3570 579944
rect 3424 576836 3476 576842
rect 3424 576778 3476 576784
rect 3422 566944 3478 566953
rect 3422 566879 3478 566888
rect 3330 553888 3386 553897
rect 3330 553823 3386 553832
rect 3344 553450 3372 553823
rect 3332 553444 3384 553450
rect 3332 553386 3384 553392
rect 3436 536790 3464 566879
rect 11716 540258 11744 618258
rect 14476 541113 14504 670686
rect 29644 553444 29696 553450
rect 29644 553386 29696 553392
rect 14462 541104 14518 541113
rect 14462 541039 14518 541048
rect 11704 540252 11756 540258
rect 11704 540194 11756 540200
rect 4804 538280 4856 538286
rect 4804 538222 4856 538228
rect 3424 536784 3476 536790
rect 3424 536726 3476 536732
rect 3424 529236 3476 529242
rect 3424 529178 3476 529184
rect 3436 501809 3464 529178
rect 3514 527912 3570 527921
rect 3514 527847 3516 527856
rect 3568 527847 3570 527856
rect 3516 527818 3568 527824
rect 3514 514856 3570 514865
rect 3514 514791 3516 514800
rect 3568 514791 3570 514800
rect 3516 514762 3568 514768
rect 3422 501800 3478 501809
rect 3422 501735 3478 501744
rect 4816 476134 4844 538222
rect 29656 538218 29684 553386
rect 39316 543726 39344 683130
rect 57888 582616 57940 582622
rect 57888 582558 57940 582564
rect 50988 582480 51040 582486
rect 50988 582422 51040 582428
rect 41328 571396 41380 571402
rect 41328 571338 41380 571344
rect 39304 543720 39356 543726
rect 39304 543662 39356 543668
rect 29644 538212 29696 538218
rect 29644 538154 29696 538160
rect 7564 514820 7616 514826
rect 7564 514762 7616 514768
rect 2780 476128 2832 476134
rect 2780 476070 2832 476076
rect 3424 476128 3476 476134
rect 3424 476070 3476 476076
rect 4804 476128 4856 476134
rect 4804 476070 4856 476076
rect 2792 475697 2820 476070
rect 2778 475688 2834 475697
rect 2778 475623 2834 475632
rect 3146 449576 3202 449585
rect 3146 449511 3202 449520
rect 3160 448594 3188 449511
rect 3148 448588 3200 448594
rect 3148 448530 3200 448536
rect 2964 411256 3016 411262
rect 2964 411198 3016 411204
rect 2976 410553 3004 411198
rect 2962 410544 3018 410553
rect 2962 410479 3018 410488
rect 3436 387802 3464 476070
rect 3514 462632 3570 462641
rect 3514 462567 3570 462576
rect 3528 462398 3556 462567
rect 3516 462392 3568 462398
rect 3516 462334 3568 462340
rect 7576 441590 7604 514762
rect 32404 462392 32456 462398
rect 32404 462334 32456 462340
rect 11704 448588 11756 448594
rect 11704 448530 11756 448536
rect 7564 441584 7616 441590
rect 7564 441526 7616 441532
rect 3516 423632 3568 423638
rect 3514 423600 3516 423609
rect 3568 423600 3570 423609
rect 3514 423535 3570 423544
rect 7564 397520 7616 397526
rect 3514 397488 3570 397497
rect 7564 397462 7616 397468
rect 3514 397423 3570 397432
rect 3424 387796 3476 387802
rect 3424 387738 3476 387744
rect 3528 386345 3556 397423
rect 3514 386336 3570 386345
rect 3514 386271 3570 386280
rect 3424 380928 3476 380934
rect 3424 380870 3476 380876
rect 3436 371385 3464 380870
rect 3422 371376 3478 371385
rect 3422 371311 3478 371320
rect 7576 358698 7604 397462
rect 11716 389201 11744 448530
rect 17224 436144 17276 436150
rect 17224 436086 17276 436092
rect 11702 389192 11758 389201
rect 11702 389127 11758 389136
rect 3240 358692 3292 358698
rect 3240 358634 3292 358640
rect 7564 358692 7616 358698
rect 7564 358634 7616 358640
rect 3252 358465 3280 358634
rect 3238 358456 3294 358465
rect 3238 358391 3294 358400
rect 3422 345400 3478 345409
rect 3422 345335 3424 345344
rect 3476 345335 3478 345344
rect 7564 345364 7616 345370
rect 3424 345306 3476 345312
rect 7564 345306 7616 345312
rect 4068 319456 4120 319462
rect 4068 319398 4120 319404
rect 4080 319297 4108 319398
rect 4066 319288 4122 319297
rect 4066 319223 4122 319232
rect 1306 309224 1362 309233
rect 1306 309159 1362 309168
rect 572 4820 624 4826
rect 572 4762 624 4768
rect 584 480 612 4762
rect 1320 3466 1348 309159
rect 3238 306232 3294 306241
rect 3238 306167 3294 306176
rect 3252 305046 3280 306167
rect 3240 305040 3292 305046
rect 3240 304982 3292 304988
rect 3422 293176 3478 293185
rect 3422 293111 3478 293120
rect 3148 255264 3200 255270
rect 3148 255206 3200 255212
rect 3160 254153 3188 255206
rect 3146 254144 3202 254153
rect 3146 254079 3202 254088
rect 3436 227730 3464 293111
rect 3514 283248 3570 283257
rect 3514 283183 3570 283192
rect 3528 267209 3556 283183
rect 4080 279478 4108 319223
rect 7576 288386 7604 345306
rect 12348 332648 12400 332654
rect 12348 332590 12400 332596
rect 7564 288380 7616 288386
rect 7564 288322 7616 288328
rect 4068 279472 4120 279478
rect 4068 279414 4120 279420
rect 3514 267200 3570 267209
rect 3514 267135 3570 267144
rect 3516 241460 3568 241466
rect 3516 241402 3568 241408
rect 3528 241097 3556 241402
rect 3514 241088 3570 241097
rect 3514 241023 3570 241032
rect 3516 235272 3568 235278
rect 3516 235214 3568 235220
rect 3424 227724 3476 227730
rect 3424 227666 3476 227672
rect 3528 219434 3556 235214
rect 6826 232520 6882 232529
rect 6826 232455 6882 232464
rect 4066 220144 4122 220153
rect 4066 220079 4122 220088
rect 3436 219406 3556 219434
rect 3436 214985 3464 219406
rect 3422 214976 3478 214985
rect 3422 214911 3478 214920
rect 3436 204270 3464 214911
rect 3424 204264 3476 204270
rect 3424 204206 3476 204212
rect 3240 202156 3292 202162
rect 3240 202098 3292 202104
rect 3252 201929 3280 202098
rect 3238 201920 3294 201929
rect 3238 201855 3294 201864
rect 3884 192500 3936 192506
rect 3884 192442 3936 192448
rect 3896 190454 3924 192442
rect 3896 190426 4016 190454
rect 3424 189032 3476 189038
rect 3424 188974 3476 188980
rect 3436 188873 3464 188974
rect 3422 188864 3478 188873
rect 3422 188799 3478 188808
rect 3424 162920 3476 162926
rect 3422 162888 3424 162897
rect 3476 162888 3478 162897
rect 3422 162823 3478 162832
rect 3330 149832 3386 149841
rect 3330 149767 3386 149776
rect 3344 145586 3372 149767
rect 3332 145580 3384 145586
rect 3332 145522 3384 145528
rect 3240 137964 3292 137970
rect 3240 137906 3292 137912
rect 3252 136785 3280 137906
rect 3238 136776 3294 136785
rect 3238 136711 3294 136720
rect 3424 135924 3476 135930
rect 3424 135866 3476 135872
rect 3436 110673 3464 135866
rect 3422 110664 3478 110673
rect 3422 110599 3478 110608
rect 3424 97980 3476 97986
rect 3424 97922 3476 97928
rect 3436 97617 3464 97922
rect 3422 97608 3478 97617
rect 3422 97543 3478 97552
rect 3148 85536 3200 85542
rect 3148 85478 3200 85484
rect 3160 84697 3188 85478
rect 3146 84688 3202 84697
rect 3146 84623 3202 84632
rect 3422 83464 3478 83473
rect 3422 83399 3478 83408
rect 3436 71641 3464 83399
rect 3422 71632 3478 71641
rect 3422 71567 3478 71576
rect 2964 59356 3016 59362
rect 2964 59298 3016 59304
rect 2976 58585 3004 59298
rect 2962 58576 3018 58585
rect 2962 58511 3018 58520
rect 3424 45552 3476 45558
rect 3422 45520 3424 45529
rect 3476 45520 3478 45529
rect 3422 45455 3478 45464
rect 3516 33108 3568 33114
rect 3516 33050 3568 33056
rect 3528 32473 3556 33050
rect 3514 32464 3570 32473
rect 3514 32399 3570 32408
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 2688 10328 2740 10334
rect 2688 10270 2740 10276
rect 2700 3534 2728 10270
rect 3424 6656 3476 6662
rect 3424 6598 3476 6604
rect 3436 6497 3464 6598
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 3988 3534 4016 190426
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 2688 3528 2740 3534
rect 2688 3470 2740 3476
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 3976 3528 4028 3534
rect 3976 3470 4028 3476
rect 1308 3460 1360 3466
rect 1308 3402 1360 3408
rect 1688 480 1716 3470
rect 2884 480 2912 3470
rect 4080 480 4108 220079
rect 5448 186992 5500 186998
rect 5448 186934 5500 186940
rect 5460 6914 5488 186934
rect 6840 6914 6868 232455
rect 7564 204264 7616 204270
rect 7564 204206 7616 204212
rect 7576 113830 7604 204206
rect 10966 146976 11022 146985
rect 10966 146911 11022 146920
rect 7564 113824 7616 113830
rect 7564 113766 7616 113772
rect 7564 106344 7616 106350
rect 7564 106286 7616 106292
rect 5276 6886 5488 6914
rect 6472 6886 6868 6914
rect 5276 480 5304 6886
rect 6472 480 6500 6886
rect 7576 6662 7604 106286
rect 7564 6656 7616 6662
rect 7564 6598 7616 6604
rect 8760 3596 8812 3602
rect 8760 3538 8812 3544
rect 7656 2100 7708 2106
rect 7656 2042 7708 2048
rect 7668 480 7696 2042
rect 8772 480 8800 3538
rect 10980 3534 11008 146911
rect 12360 3534 12388 332590
rect 17236 319462 17264 436086
rect 32416 388385 32444 462334
rect 39304 451308 39356 451314
rect 39304 451250 39356 451256
rect 37096 445868 37148 445874
rect 37096 445810 37148 445816
rect 33784 443012 33836 443018
rect 33784 442954 33836 442960
rect 33796 411262 33824 442954
rect 33784 411256 33836 411262
rect 33784 411198 33836 411204
rect 32402 388376 32458 388385
rect 32402 388311 32458 388320
rect 35808 334008 35860 334014
rect 35808 333950 35860 333956
rect 22006 324456 22062 324465
rect 22006 324391 22062 324400
rect 17224 319456 17276 319462
rect 17224 319398 17276 319404
rect 17866 307864 17922 307873
rect 17866 307799 17922 307808
rect 16486 297392 16542 297401
rect 16486 297327 16542 297336
rect 14464 280220 14516 280226
rect 14464 280162 14516 280168
rect 14476 255270 14504 280162
rect 14556 260908 14608 260914
rect 14556 260850 14608 260856
rect 14464 255264 14516 255270
rect 14464 255206 14516 255212
rect 14568 241466 14596 260850
rect 14556 241460 14608 241466
rect 14556 241402 14608 241408
rect 15106 236600 15162 236609
rect 15106 236535 15162 236544
rect 15120 6914 15148 236535
rect 14752 6886 15148 6914
rect 9956 3528 10008 3534
rect 9956 3470 10008 3476
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 11152 3528 11204 3534
rect 11152 3470 11204 3476
rect 12348 3528 12400 3534
rect 12348 3470 12400 3476
rect 9968 480 9996 3470
rect 11164 480 11192 3470
rect 13544 3460 13596 3466
rect 13544 3402 13596 3408
rect 12348 3392 12400 3398
rect 12348 3334 12400 3340
rect 12360 480 12388 3334
rect 13556 480 13584 3402
rect 14752 480 14780 6886
rect 16500 3534 16528 297327
rect 17224 185632 17276 185638
rect 17224 185574 17276 185580
rect 15936 3528 15988 3534
rect 15936 3470 15988 3476
rect 16488 3528 16540 3534
rect 16488 3470 16540 3476
rect 17040 3528 17092 3534
rect 17040 3470 17092 3476
rect 15948 480 15976 3470
rect 17052 480 17080 3470
rect 17236 2106 17264 185574
rect 17880 3534 17908 307799
rect 18604 305040 18656 305046
rect 18604 304982 18656 304988
rect 18616 253230 18644 304982
rect 18604 253224 18656 253230
rect 18604 253166 18656 253172
rect 18604 230580 18656 230586
rect 18604 230522 18656 230528
rect 18616 189038 18644 230522
rect 19246 221504 19302 221513
rect 19246 221439 19302 221448
rect 18604 189032 18656 189038
rect 18604 188974 18656 188980
rect 19260 3534 19288 221439
rect 20628 196648 20680 196654
rect 20628 196590 20680 196596
rect 17868 3528 17920 3534
rect 17868 3470 17920 3476
rect 18236 3528 18288 3534
rect 18236 3470 18288 3476
rect 19248 3528 19300 3534
rect 19248 3470 19300 3476
rect 17224 2100 17276 2106
rect 17224 2042 17276 2048
rect 18248 480 18276 3470
rect 19432 2100 19484 2106
rect 19432 2042 19484 2048
rect 19444 480 19472 2042
rect 20640 480 20668 196590
rect 22020 6914 22048 324391
rect 33782 314800 33838 314809
rect 33782 314735 33838 314744
rect 22742 313304 22798 313313
rect 22742 313239 22798 313248
rect 21836 6886 22048 6914
rect 21836 480 21864 6886
rect 22756 3602 22784 313239
rect 30286 311944 30342 311953
rect 30286 311879 30342 311888
rect 26146 302560 26202 302569
rect 26146 302495 26202 302504
rect 24766 233880 24822 233889
rect 24766 233815 24822 233824
rect 23386 203552 23442 203561
rect 23386 203487 23442 203496
rect 23400 6914 23428 203487
rect 23032 6886 23428 6914
rect 22744 3596 22796 3602
rect 22744 3538 22796 3544
rect 23032 480 23060 6886
rect 24780 3534 24808 233815
rect 24216 3528 24268 3534
rect 24216 3470 24268 3476
rect 24768 3528 24820 3534
rect 24768 3470 24820 3476
rect 24228 480 24256 3470
rect 26160 3194 26188 302495
rect 27528 188352 27580 188358
rect 27528 188294 27580 188300
rect 27540 3534 27568 188294
rect 28908 184204 28960 184210
rect 28908 184146 28960 184152
rect 26516 3528 26568 3534
rect 26516 3470 26568 3476
rect 27528 3528 27580 3534
rect 27528 3470 27580 3476
rect 25320 3188 25372 3194
rect 25320 3130 25372 3136
rect 26148 3188 26200 3194
rect 26148 3130 26200 3136
rect 25332 480 25360 3130
rect 26528 480 26556 3470
rect 27712 3392 27764 3398
rect 27712 3334 27764 3340
rect 27724 480 27752 3334
rect 28920 480 28948 184146
rect 30300 6914 30328 311879
rect 32402 306776 32458 306785
rect 32402 306711 32458 306720
rect 31666 200696 31722 200705
rect 31666 200631 31722 200640
rect 31680 6914 31708 200631
rect 32416 6914 32444 306711
rect 33046 152416 33102 152425
rect 33046 152351 33102 152360
rect 30116 6886 30328 6914
rect 31312 6886 31708 6914
rect 32324 6886 32444 6914
rect 30116 480 30144 6886
rect 31312 480 31340 6886
rect 32324 3466 32352 6886
rect 33060 3534 33088 152351
rect 32404 3528 32456 3534
rect 32404 3470 32456 3476
rect 33048 3528 33100 3534
rect 33048 3470 33100 3476
rect 33600 3528 33652 3534
rect 33600 3470 33652 3476
rect 32312 3460 32364 3466
rect 32312 3402 32364 3408
rect 32416 480 32444 3470
rect 33612 480 33640 3470
rect 33796 3398 33824 314735
rect 34426 202192 34482 202201
rect 34426 202127 34482 202136
rect 34440 3534 34468 202127
rect 35820 3534 35848 333950
rect 37108 288386 37136 445810
rect 39316 423638 39344 451250
rect 41340 449206 41368 571338
rect 48044 560312 48096 560318
rect 48044 560254 48096 560260
rect 44088 557592 44140 557598
rect 44088 557534 44140 557540
rect 44100 453257 44128 557534
rect 44086 453248 44142 453257
rect 44086 453183 44142 453192
rect 41328 449200 41380 449206
rect 41328 449142 41380 449148
rect 48056 438870 48084 560254
rect 48228 558952 48280 558958
rect 48228 558894 48280 558900
rect 48136 442264 48188 442270
rect 48136 442206 48188 442212
rect 48044 438864 48096 438870
rect 48044 438806 48096 438812
rect 45466 434888 45522 434897
rect 45466 434823 45522 434832
rect 39304 423632 39356 423638
rect 39304 423574 39356 423580
rect 39948 415472 40000 415478
rect 39948 415414 40000 415420
rect 37188 327140 37240 327146
rect 37188 327082 37240 327088
rect 37096 288380 37148 288386
rect 37096 288322 37148 288328
rect 37108 287706 37136 288322
rect 37096 287700 37148 287706
rect 37096 287642 37148 287648
rect 37094 214568 37150 214577
rect 37094 214503 37150 214512
rect 37108 3534 37136 214503
rect 34428 3528 34480 3534
rect 34428 3470 34480 3476
rect 34796 3528 34848 3534
rect 34796 3470 34848 3476
rect 35808 3528 35860 3534
rect 35808 3470 35860 3476
rect 35992 3528 36044 3534
rect 35992 3470 36044 3476
rect 37096 3528 37148 3534
rect 37096 3470 37148 3476
rect 33784 3392 33836 3398
rect 33784 3334 33836 3340
rect 34808 480 34836 3470
rect 36004 480 36032 3470
rect 37200 480 37228 327082
rect 39960 298217 39988 415414
rect 41328 411936 41380 411942
rect 41328 411878 41380 411884
rect 41142 310584 41198 310593
rect 41142 310519 41198 310528
rect 39946 298208 40002 298217
rect 39946 298143 40002 298152
rect 39856 290488 39908 290494
rect 39856 290430 39908 290436
rect 39304 262880 39356 262886
rect 39304 262822 39356 262828
rect 39316 235278 39344 262822
rect 39304 235272 39356 235278
rect 39304 235214 39356 235220
rect 38566 224224 38622 224233
rect 38566 224159 38622 224168
rect 38580 6914 38608 224159
rect 39868 141438 39896 290430
rect 39960 264246 39988 298143
rect 39948 264240 40000 264246
rect 39948 264182 40000 264188
rect 39946 235240 40002 235249
rect 39946 235175 40002 235184
rect 39856 141432 39908 141438
rect 39856 141374 39908 141380
rect 39960 6914 39988 235175
rect 38396 6886 38608 6914
rect 39592 6886 39988 6914
rect 38396 480 38424 6886
rect 39592 480 39620 6886
rect 41156 3534 41184 310519
rect 41340 309806 41368 411878
rect 44088 409148 44140 409154
rect 44088 409090 44140 409096
rect 41328 309800 41380 309806
rect 41328 309742 41380 309748
rect 41340 296714 41368 309742
rect 41248 296686 41368 296714
rect 41248 260137 41276 296686
rect 43996 271924 44048 271930
rect 43996 271866 44048 271872
rect 41234 260128 41290 260137
rect 41234 260063 41290 260072
rect 41236 249824 41288 249830
rect 41236 249766 41288 249772
rect 41248 101454 41276 249766
rect 42706 197976 42762 197985
rect 42706 197911 42762 197920
rect 41236 101448 41288 101454
rect 41236 101390 41288 101396
rect 42720 3534 42748 197911
rect 44008 155242 44036 271866
rect 44100 255921 44128 409090
rect 45480 285598 45508 434823
rect 46848 427848 46900 427854
rect 46848 427790 46900 427796
rect 45468 285592 45520 285598
rect 45468 285534 45520 285540
rect 45376 279472 45428 279478
rect 45376 279414 45428 279420
rect 44086 255912 44142 255921
rect 44086 255847 44142 255856
rect 44088 193860 44140 193866
rect 44088 193802 44140 193808
rect 43996 155236 44048 155242
rect 43996 155178 44048 155184
rect 44008 121446 44036 155178
rect 43996 121440 44048 121446
rect 43996 121382 44048 121388
rect 43996 29640 44048 29646
rect 43996 29582 44048 29588
rect 44008 3534 44036 29582
rect 40684 3528 40736 3534
rect 40684 3470 40736 3476
rect 41144 3528 41196 3534
rect 41144 3470 41196 3476
rect 41880 3528 41932 3534
rect 41880 3470 41932 3476
rect 42708 3528 42760 3534
rect 42708 3470 42760 3476
rect 43076 3528 43128 3534
rect 43076 3470 43128 3476
rect 43996 3528 44048 3534
rect 43996 3470 44048 3476
rect 44100 3482 44128 193802
rect 45388 158030 45416 279414
rect 46860 271182 46888 427790
rect 48044 421592 48096 421598
rect 48044 421534 48096 421540
rect 46848 271176 46900 271182
rect 46848 271118 46900 271124
rect 48056 265674 48084 421534
rect 48148 285530 48176 442206
rect 48240 399537 48268 558894
rect 50804 534744 50856 534750
rect 50804 534686 50856 534692
rect 49608 413296 49660 413302
rect 49608 413238 49660 413244
rect 48226 399528 48282 399537
rect 48226 399463 48282 399472
rect 48136 285524 48188 285530
rect 48136 285466 48188 285472
rect 48044 265668 48096 265674
rect 48044 265610 48096 265616
rect 46846 254008 46902 254017
rect 46846 253943 46902 253952
rect 45466 204912 45522 204921
rect 45466 204847 45522 204856
rect 45376 158024 45428 158030
rect 45376 157966 45428 157972
rect 40696 480 40724 3470
rect 41892 480 41920 3470
rect 43088 480 43116 3470
rect 44100 3454 44312 3482
rect 44284 480 44312 3454
rect 45480 480 45508 204847
rect 46204 142180 46256 142186
rect 46204 142122 46256 142128
rect 46216 97986 46244 142122
rect 46860 105602 46888 253943
rect 48148 217326 48176 285466
rect 49620 258738 49648 413238
rect 50816 412622 50844 534686
rect 51000 445738 51028 582422
rect 53564 579692 53616 579698
rect 53564 579634 53616 579640
rect 52368 563100 52420 563106
rect 52368 563042 52420 563048
rect 50988 445732 51040 445738
rect 50988 445674 51040 445680
rect 52380 442270 52408 563042
rect 52368 442264 52420 442270
rect 52368 442206 52420 442212
rect 53576 433401 53604 579634
rect 56508 564460 56560 564466
rect 56508 564402 56560 564408
rect 55128 549296 55180 549302
rect 55128 549238 55180 549244
rect 55036 533384 55088 533390
rect 55036 533326 55088 533332
rect 53656 518220 53708 518226
rect 53656 518162 53708 518168
rect 53562 433392 53618 433401
rect 53562 433327 53618 433336
rect 50896 426488 50948 426494
rect 50896 426430 50948 426436
rect 50804 412616 50856 412622
rect 50804 412558 50856 412564
rect 50816 411942 50844 412558
rect 50804 411936 50856 411942
rect 50804 411878 50856 411884
rect 50712 379568 50764 379574
rect 50712 379510 50764 379516
rect 49608 258732 49660 258738
rect 49608 258674 49660 258680
rect 50724 258058 50752 379510
rect 50908 272542 50936 426430
rect 52368 423632 52420 423638
rect 52368 423574 52420 423580
rect 50988 410576 51040 410582
rect 50988 410518 51040 410524
rect 51000 380866 51028 410518
rect 52276 407176 52328 407182
rect 52276 407118 52328 407124
rect 50988 380860 51040 380866
rect 50988 380802 51040 380808
rect 51000 379574 51028 380802
rect 50988 379568 51040 379574
rect 50988 379510 51040 379516
rect 52288 379506 52316 407118
rect 52276 379500 52328 379506
rect 52276 379442 52328 379448
rect 50988 285796 51040 285802
rect 50988 285738 51040 285744
rect 50896 272536 50948 272542
rect 50896 272478 50948 272484
rect 50802 261488 50858 261497
rect 50802 261423 50858 261432
rect 50712 258052 50764 258058
rect 50712 257994 50764 258000
rect 49606 229800 49662 229809
rect 49606 229735 49662 229744
rect 48226 225584 48282 225593
rect 48226 225519 48282 225528
rect 48136 217320 48188 217326
rect 48136 217262 48188 217268
rect 46848 105596 46900 105602
rect 46848 105538 46900 105544
rect 46204 97980 46256 97986
rect 46204 97922 46256 97928
rect 46848 31068 46900 31074
rect 46848 31010 46900 31016
rect 46860 6914 46888 31010
rect 48240 6914 48268 225519
rect 46676 6886 46888 6914
rect 47872 6886 48268 6914
rect 46676 480 46704 6886
rect 47872 480 47900 6886
rect 49620 3534 49648 229735
rect 50710 151056 50766 151065
rect 50710 150991 50766 151000
rect 50724 3534 50752 150991
rect 50816 112470 50844 261423
rect 50896 240780 50948 240786
rect 50896 240722 50948 240728
rect 50804 112464 50856 112470
rect 50804 112406 50856 112412
rect 50908 90409 50936 240722
rect 51000 132462 51028 285738
rect 51724 285592 51776 285598
rect 51724 285534 51776 285540
rect 51736 138718 51764 285534
rect 52288 258074 52316 379442
rect 52380 267034 52408 423574
rect 53668 409834 53696 518162
rect 53748 436212 53800 436218
rect 53748 436154 53800 436160
rect 52460 409828 52512 409834
rect 52460 409770 52512 409776
rect 53656 409828 53708 409834
rect 53656 409770 53708 409776
rect 52472 409154 52500 409770
rect 52460 409148 52512 409154
rect 52460 409090 52512 409096
rect 53656 400240 53708 400246
rect 53656 400182 53708 400188
rect 53668 291854 53696 400182
rect 53656 291848 53708 291854
rect 53656 291790 53708 291796
rect 53564 278724 53616 278730
rect 53564 278666 53616 278672
rect 53576 278050 53604 278666
rect 53564 278044 53616 278050
rect 53564 277986 53616 277992
rect 52368 267028 52420 267034
rect 52368 266970 52420 266976
rect 52288 258046 52408 258074
rect 52380 255241 52408 258046
rect 52366 255232 52422 255241
rect 52366 255167 52422 255176
rect 52380 254017 52408 255167
rect 53472 254584 53524 254590
rect 53472 254526 53524 254532
rect 52366 254008 52422 254017
rect 52366 253943 52422 253952
rect 52368 238808 52420 238814
rect 52368 238750 52420 238756
rect 52380 209681 52408 238750
rect 53484 237425 53512 254526
rect 53470 237416 53526 237425
rect 53470 237351 53526 237360
rect 53576 224262 53604 277986
rect 53668 251190 53696 291790
rect 53760 278730 53788 436154
rect 55048 435402 55076 533326
rect 55036 435396 55088 435402
rect 55036 435338 55088 435344
rect 55048 431954 55076 435338
rect 54956 431926 55076 431954
rect 54956 423638 54984 431926
rect 55036 423700 55088 423706
rect 55036 423642 55088 423648
rect 54944 423632 54996 423638
rect 54944 423574 54996 423580
rect 54944 403028 54996 403034
rect 54944 402970 54996 402976
rect 53748 278724 53800 278730
rect 53748 278666 53800 278672
rect 53748 273964 53800 273970
rect 53748 273906 53800 273912
rect 53656 251184 53708 251190
rect 53656 251126 53708 251132
rect 53654 237416 53710 237425
rect 53654 237351 53710 237360
rect 53564 224256 53616 224262
rect 53564 224198 53616 224204
rect 53564 210452 53616 210458
rect 53564 210394 53616 210400
rect 52366 209672 52422 209681
rect 52366 209607 52422 209616
rect 51816 162920 51868 162926
rect 51816 162862 51868 162868
rect 51828 144906 51856 162862
rect 51816 144900 51868 144906
rect 51816 144842 51868 144848
rect 51724 138712 51776 138718
rect 51724 138654 51776 138660
rect 50988 132456 51040 132462
rect 50988 132398 51040 132404
rect 52380 92478 52408 209607
rect 53470 158808 53526 158817
rect 53470 158743 53526 158752
rect 53484 124914 53512 158743
rect 53472 124908 53524 124914
rect 53472 124850 53524 124856
rect 52368 92472 52420 92478
rect 52368 92414 52420 92420
rect 50894 90400 50950 90409
rect 50894 90335 50950 90344
rect 53576 89690 53604 210394
rect 53668 104854 53696 237351
rect 53760 158817 53788 273906
rect 54852 268388 54904 268394
rect 54852 268330 54904 268336
rect 53746 158808 53802 158817
rect 53746 158743 53802 158752
rect 54864 152522 54892 268330
rect 54956 251870 54984 402970
rect 55048 268394 55076 423642
rect 55140 391513 55168 549238
rect 56416 392012 56468 392018
rect 56416 391954 56468 391960
rect 55126 391504 55182 391513
rect 55126 391439 55182 391448
rect 56428 358057 56456 391954
rect 56520 389842 56548 564402
rect 57796 553444 57848 553450
rect 57796 553386 57848 553392
rect 57704 465044 57756 465050
rect 57704 464986 57756 464992
rect 57716 463758 57744 464986
rect 57704 463752 57756 463758
rect 57704 463694 57756 463700
rect 57716 422249 57744 463694
rect 57702 422240 57758 422249
rect 57702 422175 57758 422184
rect 57716 421598 57744 422175
rect 57704 421592 57756 421598
rect 57704 421534 57756 421540
rect 57808 415478 57836 553386
rect 57900 465050 57928 582558
rect 59268 581052 59320 581058
rect 59268 580994 59320 581000
rect 59176 539640 59228 539646
rect 59176 539582 59228 539588
rect 57888 465044 57940 465050
rect 57888 464986 57940 464992
rect 57888 425740 57940 425746
rect 57888 425682 57940 425688
rect 57796 415472 57848 415478
rect 57796 415414 57848 415420
rect 56508 389836 56560 389842
rect 56508 389778 56560 389784
rect 57704 387864 57756 387870
rect 57704 387806 57756 387812
rect 56414 358048 56470 358057
rect 56414 357983 56470 357992
rect 55126 289232 55182 289241
rect 55126 289167 55182 289176
rect 55036 268388 55088 268394
rect 55036 268330 55088 268336
rect 54944 251864 54996 251870
rect 54944 251806 54996 251812
rect 54956 248414 54984 251806
rect 55140 249082 55168 289167
rect 56324 288516 56376 288522
rect 56324 288458 56376 288464
rect 55128 249076 55180 249082
rect 55128 249018 55180 249024
rect 55864 249076 55916 249082
rect 55864 249018 55916 249024
rect 54956 248386 55076 248414
rect 54944 165640 54996 165646
rect 54944 165582 54996 165588
rect 54852 152516 54904 152522
rect 54852 152458 54904 152464
rect 53746 148336 53802 148345
rect 53746 148271 53802 148280
rect 53656 104848 53708 104854
rect 53656 104790 53708 104796
rect 53564 89684 53616 89690
rect 53564 89626 53616 89632
rect 53656 47592 53708 47598
rect 53656 47534 53708 47540
rect 53668 3534 53696 47534
rect 48964 3528 49016 3534
rect 48964 3470 49016 3476
rect 49608 3528 49660 3534
rect 49608 3470 49660 3476
rect 50160 3528 50212 3534
rect 50160 3470 50212 3476
rect 50712 3528 50764 3534
rect 50712 3470 50764 3476
rect 52552 3528 52604 3534
rect 52552 3470 52604 3476
rect 53656 3528 53708 3534
rect 53656 3470 53708 3476
rect 48976 480 49004 3470
rect 50172 480 50200 3470
rect 51356 3460 51408 3466
rect 51356 3402 51408 3408
rect 51368 480 51396 3402
rect 52564 480 52592 3470
rect 53760 480 53788 148271
rect 54864 118658 54892 152458
rect 54956 126954 54984 165582
rect 54944 126948 54996 126954
rect 54944 126890 54996 126896
rect 54852 118652 54904 118658
rect 54852 118594 54904 118600
rect 55048 102814 55076 248386
rect 55126 189680 55182 189689
rect 55126 189615 55182 189624
rect 55036 102808 55088 102814
rect 55036 102750 55088 102756
rect 55036 37936 55088 37942
rect 55036 37878 55088 37884
rect 55048 6914 55076 37878
rect 54956 6886 55076 6914
rect 54956 480 54984 6886
rect 55140 3058 55168 189615
rect 55876 99482 55904 249018
rect 56336 236706 56364 288458
rect 56428 244254 56456 357983
rect 57244 265668 57296 265674
rect 57244 265610 57296 265616
rect 57256 264994 57284 265610
rect 57244 264988 57296 264994
rect 57244 264930 57296 264936
rect 56508 260160 56560 260166
rect 56508 260102 56560 260108
rect 56416 244248 56468 244254
rect 56416 244190 56468 244196
rect 56324 236700 56376 236706
rect 56324 236642 56376 236648
rect 56414 151192 56470 151201
rect 56414 151127 56470 151136
rect 56428 118590 56456 151127
rect 56416 118584 56468 118590
rect 56416 118526 56468 118532
rect 56520 111790 56548 260102
rect 57716 242185 57744 387806
rect 57796 282192 57848 282198
rect 57796 282134 57848 282140
rect 57702 242176 57758 242185
rect 57702 242111 57758 242120
rect 57704 156052 57756 156058
rect 57704 155994 57756 156000
rect 57242 136776 57298 136785
rect 57242 136711 57298 136720
rect 56508 111784 56560 111790
rect 56508 111726 56560 111732
rect 55864 99476 55916 99482
rect 55864 99418 55916 99424
rect 57256 59362 57284 136711
rect 57716 122806 57744 155994
rect 57808 131102 57836 282134
rect 57900 269074 57928 425682
rect 59084 393372 59136 393378
rect 59084 393314 59136 393320
rect 58900 376032 58952 376038
rect 58900 375974 58952 375980
rect 57888 269068 57940 269074
rect 57888 269010 57940 269016
rect 57888 264988 57940 264994
rect 57888 264930 57940 264936
rect 57900 153882 57928 264930
rect 58912 241466 58940 375974
rect 59096 367062 59124 393314
rect 59188 389337 59216 539582
rect 59280 413302 59308 580994
rect 64788 579760 64840 579766
rect 64788 579702 64840 579708
rect 63408 572756 63460 572762
rect 63408 572698 63460 572704
rect 61936 570036 61988 570042
rect 61936 569978 61988 569984
rect 60554 537432 60610 537441
rect 60554 537367 60610 537376
rect 59268 413296 59320 413302
rect 59268 413238 59320 413244
rect 60568 393446 60596 537367
rect 61948 448594 61976 569978
rect 62028 565888 62080 565894
rect 62028 565830 62080 565836
rect 61936 448588 61988 448594
rect 61936 448530 61988 448536
rect 61750 439512 61806 439521
rect 61750 439447 61806 439456
rect 60646 425096 60702 425105
rect 60646 425031 60702 425040
rect 60556 393440 60608 393446
rect 60556 393382 60608 393388
rect 59174 389328 59230 389337
rect 59174 389263 59230 389272
rect 59084 367056 59136 367062
rect 59084 366998 59136 367004
rect 59096 354674 59124 366998
rect 59004 354646 59124 354674
rect 59004 245614 59032 354646
rect 60556 304292 60608 304298
rect 60556 304234 60608 304240
rect 60568 279478 60596 304234
rect 60556 279472 60608 279478
rect 60556 279414 60608 279420
rect 60464 272536 60516 272542
rect 60464 272478 60516 272484
rect 60476 270745 60504 272478
rect 60556 271176 60608 271182
rect 60556 271118 60608 271124
rect 60462 270736 60518 270745
rect 60462 270671 60518 270680
rect 59176 270496 59228 270502
rect 59176 270438 59228 270444
rect 59084 263628 59136 263634
rect 59084 263570 59136 263576
rect 58992 245608 59044 245614
rect 58992 245550 59044 245556
rect 58532 241460 58584 241466
rect 58532 241402 58584 241408
rect 58900 241460 58952 241466
rect 58900 241402 58952 241408
rect 58544 240786 58572 241402
rect 58532 240780 58584 240786
rect 58532 240722 58584 240728
rect 57888 153876 57940 153882
rect 57888 153818 57940 153824
rect 57796 131096 57848 131102
rect 57796 131038 57848 131044
rect 57704 122800 57756 122806
rect 57704 122742 57756 122748
rect 57900 115938 57928 153818
rect 59096 139466 59124 263570
rect 59084 139460 59136 139466
rect 59084 139402 59136 139408
rect 58622 135416 58678 135425
rect 58622 135351 58678 135360
rect 57888 115932 57940 115938
rect 57888 115874 57940 115880
rect 57244 59356 57296 59362
rect 57244 59298 57296 59304
rect 57888 58676 57940 58682
rect 57888 58618 57940 58624
rect 57900 3534 57928 58618
rect 58636 33114 58664 135351
rect 59096 114510 59124 139402
rect 59188 138145 59216 270438
rect 59266 258224 59322 258233
rect 59266 258159 59322 258168
rect 59280 254590 59308 258159
rect 59268 254584 59320 254590
rect 59268 254526 59320 254532
rect 59268 242956 59320 242962
rect 59268 242898 59320 242904
rect 59280 191146 59308 242898
rect 59268 191140 59320 191146
rect 59268 191082 59320 191088
rect 59174 138136 59230 138145
rect 59174 138071 59230 138080
rect 59188 120018 59216 138071
rect 59176 120012 59228 120018
rect 59176 119954 59228 119960
rect 59084 114504 59136 114510
rect 59084 114446 59136 114452
rect 59280 95198 59308 191082
rect 60476 146946 60504 270671
rect 60568 270570 60596 271118
rect 60556 270564 60608 270570
rect 60556 270506 60608 270512
rect 60464 146940 60516 146946
rect 60464 146882 60516 146888
rect 60476 120086 60504 146882
rect 60568 142254 60596 270506
rect 60660 270502 60688 425031
rect 61658 311128 61714 311137
rect 61658 311063 61714 311072
rect 61672 277370 61700 311063
rect 61764 290494 61792 439447
rect 61842 436112 61898 436121
rect 61842 436047 61898 436056
rect 61856 311137 61884 436047
rect 61948 429146 61976 448530
rect 61936 429140 61988 429146
rect 61936 429082 61988 429088
rect 62040 410582 62068 565830
rect 63316 545148 63368 545154
rect 63316 545090 63368 545096
rect 63328 496126 63356 545090
rect 63316 496120 63368 496126
rect 63316 496062 63368 496068
rect 63316 440292 63368 440298
rect 63316 440234 63368 440240
rect 62762 438152 62818 438161
rect 62762 438087 62818 438096
rect 62028 410576 62080 410582
rect 62028 410518 62080 410524
rect 62028 404388 62080 404394
rect 62028 404330 62080 404336
rect 61842 311128 61898 311137
rect 61842 311063 61898 311072
rect 61752 290488 61804 290494
rect 61752 290430 61804 290436
rect 61844 290148 61896 290154
rect 61844 290090 61896 290096
rect 61856 285705 61884 290090
rect 61842 285696 61898 285705
rect 61842 285631 61898 285640
rect 61752 280288 61804 280294
rect 61752 280230 61804 280236
rect 61660 277364 61712 277370
rect 61660 277306 61712 277312
rect 60648 270496 60700 270502
rect 60648 270438 60700 270444
rect 60660 269249 60688 270438
rect 60646 269240 60702 269249
rect 60646 269175 60702 269184
rect 60648 269068 60700 269074
rect 60648 269010 60700 269016
rect 60660 268462 60688 269010
rect 60648 268456 60700 268462
rect 60648 268398 60700 268404
rect 60660 218754 60688 268398
rect 61764 242214 61792 280230
rect 61752 242208 61804 242214
rect 61752 242150 61804 242156
rect 61856 236774 61884 285631
rect 61934 265160 61990 265169
rect 61934 265095 61990 265104
rect 61844 236768 61896 236774
rect 61844 236710 61896 236716
rect 60648 218748 60700 218754
rect 60648 218690 60700 218696
rect 60646 167648 60702 167657
rect 60646 167583 60702 167592
rect 60556 142248 60608 142254
rect 60556 142190 60608 142196
rect 60568 121378 60596 142190
rect 60556 121372 60608 121378
rect 60556 121314 60608 121320
rect 60464 120080 60516 120086
rect 60464 120022 60516 120028
rect 59268 95192 59320 95198
rect 59268 95134 59320 95140
rect 59268 46232 59320 46238
rect 59268 46174 59320 46180
rect 58624 33108 58676 33114
rect 58624 33050 58676 33056
rect 59280 3534 59308 46174
rect 60660 3534 60688 167583
rect 61842 162888 61898 162897
rect 61842 162823 61898 162832
rect 61660 128716 61712 128722
rect 61660 128658 61712 128664
rect 61672 35222 61700 128658
rect 61856 126886 61884 162823
rect 61948 147762 61976 265095
rect 62040 252770 62068 404330
rect 62776 290154 62804 438087
rect 63132 419552 63184 419558
rect 63132 419494 63184 419500
rect 62764 290148 62816 290154
rect 62764 290090 62816 290096
rect 63144 265169 63172 419494
rect 63328 419490 63356 440234
rect 63316 419484 63368 419490
rect 63316 419426 63368 419432
rect 63420 405793 63448 572698
rect 64696 547936 64748 547942
rect 64696 547878 64748 547884
rect 64604 526448 64656 526454
rect 64604 526390 64656 526396
rect 63406 405784 63462 405793
rect 63406 405719 63462 405728
rect 64616 395486 64644 526390
rect 64708 520946 64736 547878
rect 64696 520940 64748 520946
rect 64696 520882 64748 520888
rect 64800 490618 64828 579702
rect 65982 567624 66038 567633
rect 65982 567559 66038 567568
rect 65890 550896 65946 550905
rect 65890 550831 65946 550840
rect 65798 544096 65854 544105
rect 65798 544031 65854 544040
rect 64788 490612 64840 490618
rect 64788 490554 64840 490560
rect 65812 438161 65840 544031
rect 65904 532030 65932 550831
rect 65892 532024 65944 532030
rect 65892 531966 65944 531972
rect 65996 522345 66024 567559
rect 66180 566817 66208 702510
rect 68928 625864 68980 625870
rect 68928 625806 68980 625812
rect 68940 588402 68968 625806
rect 67732 588396 67784 588402
rect 67732 588338 67784 588344
rect 68928 588396 68980 588402
rect 68928 588338 68980 588344
rect 66534 580000 66590 580009
rect 66534 579935 66590 579944
rect 66548 579766 66576 579935
rect 66536 579760 66588 579766
rect 66536 579702 66588 579708
rect 67546 578640 67602 578649
rect 67546 578575 67602 578584
rect 67454 577280 67510 577289
rect 67454 577215 67510 577224
rect 66534 573200 66590 573209
rect 66534 573135 66590 573144
rect 66548 572762 66576 573135
rect 66536 572756 66588 572762
rect 66536 572698 66588 572704
rect 66534 571840 66590 571849
rect 66534 571775 66590 571784
rect 66548 571402 66576 571775
rect 66536 571396 66588 571402
rect 66536 571338 66588 571344
rect 66902 570208 66958 570217
rect 66902 570143 66958 570152
rect 66916 570042 66944 570143
rect 66904 570036 66956 570042
rect 66904 569978 66956 569984
rect 67362 568848 67418 568857
rect 67362 568783 67418 568792
rect 66166 566808 66222 566817
rect 66166 566743 66222 566752
rect 66180 565894 66208 566743
rect 66168 565888 66220 565894
rect 66168 565830 66220 565836
rect 66534 564768 66590 564777
rect 66534 564703 66590 564712
rect 66548 564466 66576 564703
rect 66536 564460 66588 564466
rect 66536 564402 66588 564408
rect 66534 563408 66590 563417
rect 66534 563343 66590 563352
rect 66548 563106 66576 563343
rect 66536 563100 66588 563106
rect 66536 563042 66588 563048
rect 66718 560688 66774 560697
rect 66718 560623 66774 560632
rect 66732 560318 66760 560623
rect 66720 560312 66772 560318
rect 66720 560254 66772 560260
rect 66718 559328 66774 559337
rect 66718 559263 66774 559272
rect 66732 558958 66760 559263
rect 66720 558952 66772 558958
rect 66720 558894 66772 558900
rect 66718 557968 66774 557977
rect 66718 557903 66774 557912
rect 66732 557598 66760 557903
rect 66720 557592 66772 557598
rect 66720 557534 66772 557540
rect 66074 555248 66130 555257
rect 66074 555183 66130 555192
rect 65982 522336 66038 522345
rect 65982 522271 66038 522280
rect 66088 501634 66116 555183
rect 66534 553752 66590 553761
rect 66534 553687 66590 553696
rect 66548 553450 66576 553687
rect 66536 553444 66588 553450
rect 66536 553386 66588 553392
rect 66534 549672 66590 549681
rect 66534 549607 66590 549616
rect 66548 549302 66576 549607
rect 66536 549296 66588 549302
rect 66536 549238 66588 549244
rect 66810 548176 66866 548185
rect 66810 548111 66866 548120
rect 66824 547942 66852 548111
rect 66812 547936 66864 547942
rect 66812 547878 66864 547884
rect 66718 545456 66774 545465
rect 66718 545391 66774 545400
rect 66732 545154 66760 545391
rect 66720 545148 66772 545154
rect 66720 545090 66772 545096
rect 67272 543720 67324 543726
rect 67272 543662 67324 543668
rect 67284 543425 67312 543662
rect 67270 543416 67326 543425
rect 67270 543351 67326 543360
rect 66442 540152 66498 540161
rect 66442 540087 66498 540096
rect 66456 539646 66484 540087
rect 66444 539640 66496 539646
rect 66444 539582 66496 539588
rect 67376 525094 67404 568783
rect 67364 525088 67416 525094
rect 67364 525030 67416 525036
rect 66076 501628 66128 501634
rect 66076 501570 66128 501576
rect 65982 475416 66038 475425
rect 65982 475351 66038 475360
rect 65798 438152 65854 438161
rect 65798 438087 65854 438096
rect 64696 434784 64748 434790
rect 64696 434726 64748 434732
rect 64604 395480 64656 395486
rect 64604 395422 64656 395428
rect 63408 307080 63460 307086
rect 63408 307022 63460 307028
rect 63224 267028 63276 267034
rect 63224 266970 63276 266976
rect 63130 265160 63186 265169
rect 63130 265095 63186 265104
rect 62118 252784 62174 252793
rect 62040 252742 62118 252770
rect 62118 252719 62174 252728
rect 62026 240272 62082 240281
rect 62026 240207 62082 240216
rect 61936 147756 61988 147762
rect 61936 147698 61988 147704
rect 61844 126880 61896 126886
rect 61844 126822 61896 126828
rect 61948 115462 61976 147698
rect 61936 115456 61988 115462
rect 61936 115398 61988 115404
rect 61752 102808 61804 102814
rect 61752 102750 61804 102756
rect 61764 81161 61792 102750
rect 61844 100768 61896 100774
rect 61844 100710 61896 100716
rect 61750 81152 61806 81161
rect 61750 81087 61806 81096
rect 61856 67590 61884 100710
rect 62040 92546 62068 240207
rect 63236 222902 63264 266970
rect 63316 266416 63368 266422
rect 63316 266358 63368 266364
rect 63224 222896 63276 222902
rect 63224 222838 63276 222844
rect 63222 161664 63278 161673
rect 63222 161599 63278 161608
rect 63132 145036 63184 145042
rect 63132 144978 63184 144984
rect 63144 117298 63172 144978
rect 63236 125390 63264 161599
rect 63328 145042 63356 266358
rect 63420 256902 63448 307022
rect 64602 291816 64658 291825
rect 64602 291751 64658 291760
rect 63408 256896 63460 256902
rect 63408 256838 63460 256844
rect 63406 252784 63462 252793
rect 63406 252719 63462 252728
rect 63316 145036 63368 145042
rect 63316 144978 63368 144984
rect 63316 141568 63368 141574
rect 63316 141510 63368 141516
rect 63224 125384 63276 125390
rect 63224 125326 63276 125332
rect 63132 117292 63184 117298
rect 63132 117234 63184 117240
rect 63224 113824 63276 113830
rect 63224 113766 63276 113772
rect 62028 92540 62080 92546
rect 62028 92482 62080 92488
rect 63236 88330 63264 113766
rect 63328 90982 63356 141510
rect 63420 103494 63448 252719
rect 64616 238746 64644 291751
rect 64708 283014 64736 434726
rect 65798 433392 65854 433401
rect 64788 433356 64840 433362
rect 65798 433327 65854 433336
rect 64788 433298 64840 433304
rect 64800 422278 64828 433298
rect 64788 422272 64840 422278
rect 64788 422214 64840 422220
rect 64788 414044 64840 414050
rect 64788 413986 64840 413992
rect 64696 283008 64748 283014
rect 64696 282950 64748 282956
rect 64604 238740 64656 238746
rect 64604 238682 64656 238688
rect 63500 158024 63552 158030
rect 63500 157966 63552 157972
rect 63512 157418 63540 157966
rect 63500 157412 63552 157418
rect 63500 157354 63552 157360
rect 64604 157412 64656 157418
rect 64604 157354 64656 157360
rect 64512 138032 64564 138038
rect 64512 137974 64564 137980
rect 64524 110430 64552 137974
rect 64616 128314 64644 157354
rect 64708 139641 64736 282950
rect 64800 261497 64828 413986
rect 65812 288425 65840 433327
rect 65904 393446 65932 393477
rect 65892 393440 65944 393446
rect 65890 393408 65892 393417
rect 65944 393408 65946 393417
rect 65890 393343 65946 393352
rect 65904 373969 65932 393343
rect 65996 389162 66024 475351
rect 67272 449948 67324 449954
rect 67272 449890 67324 449896
rect 66168 445800 66220 445806
rect 66168 445742 66220 445748
rect 66074 443048 66130 443057
rect 66074 442983 66130 442992
rect 66088 425746 66116 442983
rect 66180 431474 66208 445742
rect 67180 439544 67232 439550
rect 67180 439486 67232 439492
rect 66258 431488 66314 431497
rect 66180 431446 66258 431474
rect 66076 425740 66128 425746
rect 66076 425682 66128 425688
rect 65984 389156 66036 389162
rect 65984 389098 66036 389104
rect 66076 387864 66128 387870
rect 66076 387806 66128 387812
rect 66088 387433 66116 387806
rect 66074 387424 66130 387433
rect 66074 387359 66130 387368
rect 65984 381540 66036 381546
rect 65984 381482 66036 381488
rect 65890 373960 65946 373969
rect 65890 373895 65946 373904
rect 65798 288416 65854 288425
rect 65798 288351 65854 288360
rect 65892 282260 65944 282266
rect 65892 282202 65944 282208
rect 65904 273970 65932 282202
rect 65892 273964 65944 273970
rect 65892 273906 65944 273912
rect 64786 261488 64842 261497
rect 64786 261423 64842 261432
rect 65890 259584 65946 259593
rect 65890 259519 65946 259528
rect 64788 258732 64840 258738
rect 64788 258674 64840 258680
rect 64800 235385 64828 258674
rect 64786 235376 64842 235385
rect 64786 235311 64842 235320
rect 65904 229094 65932 259519
rect 65996 239873 66024 381482
rect 66074 288416 66130 288425
rect 66074 288351 66130 288360
rect 66088 287337 66116 288351
rect 66074 287328 66130 287337
rect 66074 287263 66130 287272
rect 66088 277394 66116 287263
rect 66180 282266 66208 431446
rect 66258 431423 66314 431432
rect 67192 430409 67220 439486
rect 67178 430400 67234 430409
rect 67178 430335 67234 430344
rect 66812 429140 66864 429146
rect 66812 429082 66864 429088
rect 66258 428224 66314 428233
rect 66258 428159 66314 428168
rect 66272 427854 66300 428159
rect 66260 427848 66312 427854
rect 66260 427790 66312 427796
rect 66824 426306 66852 429082
rect 66902 427408 66958 427417
rect 66902 427343 66958 427352
rect 66916 426494 66944 427343
rect 66904 426488 66956 426494
rect 66904 426430 66956 426436
rect 66824 426278 66944 426306
rect 66628 425740 66680 425746
rect 66628 425682 66680 425688
rect 66640 425241 66668 425682
rect 66626 425232 66682 425241
rect 66626 425167 66682 425176
rect 66810 424144 66866 424153
rect 66810 424079 66866 424088
rect 66824 423706 66852 424079
rect 66812 423700 66864 423706
rect 66812 423642 66864 423648
rect 66628 423632 66680 423638
rect 66628 423574 66680 423580
rect 66640 423337 66668 423574
rect 66626 423328 66682 423337
rect 66626 423263 66682 423272
rect 66916 422294 66944 426278
rect 66812 422272 66864 422278
rect 66810 422240 66812 422249
rect 66916 422266 67036 422294
rect 66864 422240 66866 422249
rect 66810 422175 66866 422184
rect 66902 420064 66958 420073
rect 66902 419999 66958 420008
rect 66916 419558 66944 419999
rect 66904 419552 66956 419558
rect 66904 419494 66956 419500
rect 66812 419484 66864 419490
rect 66812 419426 66864 419432
rect 66824 418985 66852 419426
rect 66810 418976 66866 418985
rect 66810 418911 66866 418920
rect 67008 417081 67036 422266
rect 66994 417072 67050 417081
rect 66994 417007 67050 417016
rect 66902 415984 66958 415993
rect 66902 415919 66958 415928
rect 66916 415478 66944 415919
rect 66904 415472 66956 415478
rect 66904 415414 66956 415420
rect 66718 414896 66774 414905
rect 66718 414831 66774 414840
rect 66732 414050 66760 414831
rect 67284 414089 67312 449890
rect 67468 441658 67496 577215
rect 67456 441652 67508 441658
rect 67456 441594 67508 441600
rect 67468 431954 67496 441594
rect 67376 431926 67496 431954
rect 67270 414080 67326 414089
rect 66720 414044 66772 414050
rect 67270 414015 67326 414024
rect 66720 413986 66772 413992
rect 66260 413296 66312 413302
rect 66260 413238 66312 413244
rect 66272 413001 66300 413238
rect 66258 412992 66314 413001
rect 66258 412927 66314 412936
rect 66812 412616 66864 412622
rect 66812 412558 66864 412564
rect 66824 411913 66852 412558
rect 66810 411904 66866 411913
rect 66810 411839 66866 411848
rect 66902 410816 66958 410825
rect 66902 410751 66958 410760
rect 66916 410582 66944 410751
rect 66904 410576 66956 410582
rect 66904 410518 66956 410524
rect 66812 409828 66864 409834
rect 66812 409770 66864 409776
rect 66824 408921 66852 409770
rect 66810 408912 66866 408921
rect 66810 408847 66866 408856
rect 66810 407824 66866 407833
rect 66810 407759 66866 407768
rect 66824 407182 66852 407759
rect 66812 407176 66864 407182
rect 66812 407118 66864 407124
rect 67376 405657 67404 431926
rect 67454 418160 67510 418169
rect 67454 418095 67510 418104
rect 67362 405648 67418 405657
rect 67362 405583 67418 405592
rect 66902 404560 66958 404569
rect 66902 404495 66958 404504
rect 66916 404394 66944 404495
rect 66904 404388 66956 404394
rect 66904 404330 66956 404336
rect 66810 403744 66866 403753
rect 66810 403679 66866 403688
rect 66824 403034 66852 403679
rect 66812 403028 66864 403034
rect 66812 402970 66864 402976
rect 67270 401704 67326 401713
rect 67270 401639 67326 401648
rect 66718 401568 66774 401577
rect 66718 401503 66774 401512
rect 66732 400246 66760 401503
rect 66720 400240 66772 400246
rect 66720 400182 66772 400188
rect 67180 395480 67232 395486
rect 67180 395422 67232 395428
rect 67192 395321 67220 395422
rect 67178 395312 67234 395321
rect 67178 395247 67234 395256
rect 66810 394496 66866 394505
rect 66810 394431 66866 394440
rect 66824 393378 66852 394431
rect 66812 393372 66864 393378
rect 66812 393314 66864 393320
rect 66258 392320 66314 392329
rect 66258 392255 66314 392264
rect 66272 392018 66300 392255
rect 66260 392012 66312 392018
rect 66260 391954 66312 391960
rect 67192 372609 67220 395247
rect 67284 378146 67312 401639
rect 67362 400480 67418 400489
rect 67362 400415 67418 400424
rect 67376 390658 67404 400415
rect 67364 390652 67416 390658
rect 67364 390594 67416 390600
rect 67272 378140 67324 378146
rect 67272 378082 67324 378088
rect 67178 372600 67234 372609
rect 67178 372535 67234 372544
rect 67468 314702 67496 418095
rect 67560 402665 67588 578575
rect 67640 576836 67692 576842
rect 67640 576778 67692 576784
rect 67652 575929 67680 576778
rect 67638 575920 67694 575929
rect 67638 575855 67694 575864
rect 67652 474065 67680 575855
rect 67744 575385 67772 588338
rect 68940 587926 68968 588338
rect 68928 587920 68980 587926
rect 68928 587862 68980 587868
rect 70320 586514 70348 702782
rect 69768 586486 70348 586514
rect 69768 581074 69796 586486
rect 71792 585177 71820 702986
rect 86224 702908 86276 702914
rect 86224 702850 86276 702856
rect 84108 702636 84160 702642
rect 84108 702578 84160 702584
rect 77208 702500 77260 702506
rect 77208 702442 77260 702448
rect 74540 656940 74592 656946
rect 74540 656882 74592 656888
rect 74552 596174 74580 656882
rect 74552 596146 74672 596174
rect 72424 585200 72476 585206
rect 71778 585168 71834 585177
rect 72424 585142 72476 585148
rect 71778 585103 71834 585112
rect 69940 582480 69992 582486
rect 69940 582422 69992 582428
rect 69032 581046 69796 581074
rect 69952 581074 69980 582422
rect 72436 581074 72464 585142
rect 74264 583840 74316 583846
rect 74264 583782 74316 583788
rect 73526 582584 73582 582593
rect 73526 582519 73582 582528
rect 73540 581074 73568 582519
rect 74276 581074 74304 583782
rect 69952 581046 70288 581074
rect 72128 581046 72464 581074
rect 73232 581046 73568 581074
rect 74152 581046 74304 581074
rect 74644 581074 74672 596146
rect 77220 590442 77248 702442
rect 79968 700324 80020 700330
rect 79968 700266 80020 700272
rect 79980 592074 80008 700266
rect 79324 592068 79376 592074
rect 79324 592010 79376 592016
rect 79968 592068 80020 592074
rect 79968 592010 80020 592016
rect 76472 590436 76524 590442
rect 76472 590378 76524 590384
rect 77208 590436 77260 590442
rect 77208 590378 77260 590384
rect 76484 589354 76512 590378
rect 76472 589348 76524 589354
rect 76472 589290 76524 589296
rect 76288 581120 76340 581126
rect 75366 581088 75422 581097
rect 74644 581046 75366 581074
rect 69032 580718 69060 581046
rect 75992 581068 76288 581074
rect 75992 581062 76340 581068
rect 76484 581074 76512 589290
rect 79336 582690 79364 592010
rect 84120 587246 84148 702578
rect 81808 587240 81860 587246
rect 81808 587182 81860 587188
rect 84108 587240 84160 587246
rect 84108 587182 84160 587188
rect 78128 582684 78180 582690
rect 78128 582626 78180 582632
rect 79324 582684 79376 582690
rect 79324 582626 79376 582632
rect 78140 581074 78168 582626
rect 79048 582412 79100 582418
rect 79048 582354 79100 582360
rect 79060 581074 79088 582354
rect 80242 581224 80298 581233
rect 80242 581159 80298 581168
rect 75992 581046 76328 581062
rect 76484 581046 76912 581074
rect 77832 581046 78168 581074
rect 78752 581046 79088 581074
rect 80256 581074 80284 581159
rect 81820 581074 81848 587182
rect 85486 582720 85542 582729
rect 85486 582655 85542 582664
rect 82726 581088 82782 581097
rect 80256 581046 80592 581074
rect 81512 581046 81848 581074
rect 82432 581046 82726 581074
rect 75366 581023 75422 581032
rect 85500 581074 85528 582655
rect 86236 582554 86264 702850
rect 89180 700330 89208 703520
rect 104808 702976 104860 702982
rect 104808 702918 104860 702924
rect 90364 702908 90416 702914
rect 90364 702850 90416 702856
rect 89168 700324 89220 700330
rect 89168 700266 89220 700272
rect 90376 596174 90404 702850
rect 94688 702772 94740 702778
rect 94688 702714 94740 702720
rect 94700 596174 94728 702714
rect 96620 702704 96672 702710
rect 96620 702646 96672 702652
rect 90376 596146 90496 596174
rect 94700 596146 94912 596174
rect 87512 585268 87564 585274
rect 87512 585210 87564 585216
rect 86224 582548 86276 582554
rect 86224 582490 86276 582496
rect 86236 581346 86264 582490
rect 86868 582412 86920 582418
rect 86868 582354 86920 582360
rect 86236 581318 86310 581346
rect 83016 581058 83352 581074
rect 82726 581023 82782 581032
rect 83004 581052 83352 581058
rect 83056 581046 83352 581052
rect 85376 581046 85528 581074
rect 86282 581060 86310 581318
rect 83004 580994 83056 581000
rect 70858 580816 70914 580825
rect 79874 580816 79930 580825
rect 70914 580774 71208 580802
rect 79672 580774 79874 580802
rect 70858 580751 70914 580760
rect 79874 580751 79930 580760
rect 84198 580816 84254 580825
rect 84254 580774 84456 580802
rect 84198 580751 84254 580760
rect 86880 580718 86908 582354
rect 87524 581074 87552 585210
rect 88248 583772 88300 583778
rect 88248 583714 88300 583720
rect 88260 581074 88288 583714
rect 90468 582622 90496 596146
rect 92110 583808 92166 583817
rect 92110 583743 92166 583752
rect 90456 582616 90508 582622
rect 90456 582558 90508 582564
rect 90272 582412 90324 582418
rect 90272 582354 90324 582360
rect 90284 581074 90312 582354
rect 87216 581046 87552 581074
rect 88136 581046 88288 581074
rect 89976 581046 90312 581074
rect 90468 581074 90496 582558
rect 92124 581074 92152 583743
rect 90468 581046 90896 581074
rect 91816 581046 92152 581074
rect 93656 581058 93808 581074
rect 93656 581052 93820 581058
rect 93656 581046 93768 581052
rect 93768 580994 93820 581000
rect 88890 580816 88946 580825
rect 92570 580816 92626 580825
rect 88946 580774 89056 580802
rect 88890 580751 88946 580760
rect 92626 580774 92736 580802
rect 92570 580751 92626 580760
rect 69020 580712 69072 580718
rect 69020 580654 69072 580660
rect 86868 580712 86920 580718
rect 86868 580654 86920 580660
rect 94576 580514 94728 580530
rect 94576 580508 94740 580514
rect 94576 580502 94688 580508
rect 94688 580450 94740 580456
rect 67730 575376 67786 575385
rect 67730 575311 67786 575320
rect 94884 567194 94912 596146
rect 95976 582412 96028 582418
rect 95976 582354 96028 582360
rect 95884 580508 95936 580514
rect 95884 580450 95936 580456
rect 95238 574832 95294 574841
rect 95238 574767 95294 574776
rect 94700 567166 94912 567194
rect 94700 558657 94728 567166
rect 94686 558648 94742 558657
rect 94686 558583 94742 558592
rect 67730 556608 67786 556617
rect 67730 556543 67786 556552
rect 67744 536110 67772 556543
rect 67822 552256 67878 552265
rect 67822 552191 67878 552200
rect 94686 552256 94742 552265
rect 94686 552191 94742 552200
rect 67836 539102 67864 552191
rect 73160 539844 73212 539850
rect 73160 539786 73212 539792
rect 91008 539844 91060 539850
rect 91008 539786 91060 539792
rect 73172 539730 73200 539786
rect 73172 539716 73416 539730
rect 73172 539702 73430 539716
rect 68816 539158 68968 539186
rect 67824 539096 67876 539102
rect 67824 539038 67876 539044
rect 67732 536104 67784 536110
rect 67732 536046 67784 536052
rect 68940 535537 68968 539158
rect 69400 539158 69736 539186
rect 70656 539158 70716 539186
rect 69400 538214 69428 539158
rect 70688 538218 70716 539158
rect 70872 539158 71576 539186
rect 71792 539158 72496 539186
rect 69032 538186 69428 538214
rect 70676 538212 70728 538218
rect 69032 536790 69060 538186
rect 70676 538154 70728 538160
rect 69020 536784 69072 536790
rect 69020 536726 69072 536732
rect 68926 535528 68982 535537
rect 68926 535463 68982 535472
rect 67732 479528 67784 479534
rect 67732 479470 67784 479476
rect 67638 474056 67694 474065
rect 67638 473991 67694 474000
rect 67640 448384 67692 448390
rect 67640 448326 67692 448332
rect 67652 418169 67680 448326
rect 67638 418160 67694 418169
rect 67638 418095 67694 418104
rect 67546 402656 67602 402665
rect 67546 402591 67602 402600
rect 67560 401713 67588 402591
rect 67546 401704 67602 401713
rect 67546 401639 67602 401648
rect 67546 399664 67602 399673
rect 67546 399599 67602 399608
rect 67560 392057 67588 399599
rect 67744 397526 67772 479470
rect 68926 471880 68982 471889
rect 68926 471815 68982 471824
rect 68940 470665 68968 471815
rect 68926 470656 68982 470665
rect 68926 470591 68982 470600
rect 68940 456074 68968 470591
rect 68928 456068 68980 456074
rect 68928 456010 68980 456016
rect 69032 440337 69060 536726
rect 70688 530602 70716 538154
rect 70676 530596 70728 530602
rect 70676 530538 70728 530544
rect 70872 528554 70900 539158
rect 70504 528526 70900 528554
rect 69664 520940 69716 520946
rect 69664 520882 69716 520888
rect 69676 465225 69704 520882
rect 69662 465216 69718 465225
rect 69662 465151 69718 465160
rect 69112 443692 69164 443698
rect 69112 443634 69164 443640
rect 69018 440328 69074 440337
rect 69018 440263 69074 440272
rect 68926 437200 68982 437209
rect 68926 437135 68982 437144
rect 68558 436248 68614 436257
rect 68558 436183 68614 436192
rect 67822 433664 67878 433673
rect 67822 433599 67878 433608
rect 67836 429865 67864 433599
rect 68572 431954 68600 436183
rect 68940 436121 68968 437135
rect 68926 436112 68982 436121
rect 68926 436047 68982 436056
rect 68940 434194 68968 436047
rect 69124 434330 69152 443634
rect 69676 441614 69704 465151
rect 70504 443057 70532 528526
rect 71688 468580 71740 468586
rect 71688 468522 71740 468528
rect 70490 443048 70546 443057
rect 70490 442983 70546 442992
rect 71134 443048 71190 443057
rect 71134 442983 71190 442992
rect 69676 441586 69888 441614
rect 69860 436218 69888 441586
rect 70504 437510 70532 442983
rect 70492 437504 70544 437510
rect 70492 437446 70544 437452
rect 69848 436212 69900 436218
rect 69848 436154 69900 436160
rect 70860 436212 70912 436218
rect 70860 436154 70912 436160
rect 69860 434330 69888 436154
rect 69124 434302 69552 434330
rect 69860 434302 70288 434330
rect 68816 434166 68968 434194
rect 70872 434058 70900 436154
rect 70872 434030 71024 434058
rect 71148 433673 71176 442983
rect 71700 442921 71728 468522
rect 71792 460193 71820 539158
rect 71872 539096 71924 539102
rect 71872 539038 71924 539044
rect 73402 539050 73430 539702
rect 86224 539640 86276 539646
rect 76746 539608 76802 539617
rect 76802 539566 77096 539594
rect 86224 539582 86276 539588
rect 76746 539543 76802 539552
rect 73632 539158 74336 539186
rect 74552 539158 75256 539186
rect 75932 539158 76176 539186
rect 77312 539158 78016 539186
rect 78692 539158 78936 539186
rect 80040 539158 80100 539186
rect 71778 460184 71834 460193
rect 71778 460119 71834 460128
rect 71686 442912 71742 442921
rect 71686 442847 71742 442856
rect 71700 441614 71728 442847
rect 71608 441586 71728 441614
rect 71608 437209 71636 441586
rect 71594 437200 71650 437209
rect 71594 437135 71650 437144
rect 71688 436144 71740 436150
rect 71884 436121 71912 539038
rect 73402 539022 73476 539050
rect 73448 536790 73476 539022
rect 73436 536784 73488 536790
rect 73436 536726 73488 536732
rect 73632 528554 73660 539158
rect 73802 535528 73858 535537
rect 73802 535463 73858 535472
rect 73172 528526 73660 528554
rect 73172 472569 73200 528526
rect 73816 487830 73844 535463
rect 73804 487824 73856 487830
rect 73804 487766 73856 487772
rect 73158 472560 73214 472569
rect 73158 472495 73214 472504
rect 72424 456884 72476 456890
rect 72424 456826 72476 456832
rect 72436 436150 72464 456826
rect 74552 455394 74580 539158
rect 75828 537532 75880 537538
rect 75828 537474 75880 537480
rect 75840 460970 75868 537474
rect 75184 460964 75236 460970
rect 75184 460906 75236 460912
rect 75828 460964 75880 460970
rect 75828 460906 75880 460912
rect 74540 455388 74592 455394
rect 74540 455330 74592 455336
rect 73252 447840 73304 447846
rect 73252 447782 73304 447788
rect 73264 441614 73292 447782
rect 73264 441586 73384 441614
rect 72424 436144 72476 436150
rect 71688 436086 71740 436092
rect 71870 436112 71926 436121
rect 71700 434330 71728 436086
rect 72424 436086 72476 436092
rect 72516 436144 72568 436150
rect 72516 436086 72568 436092
rect 72698 436112 72754 436121
rect 71870 436047 71926 436056
rect 72528 434489 72556 436086
rect 72698 436047 72754 436056
rect 72606 435024 72662 435033
rect 72606 434959 72662 434968
rect 72514 434480 72570 434489
rect 72514 434415 72570 434424
rect 72620 434330 72648 434959
rect 71576 434302 71728 434330
rect 72312 434302 72648 434330
rect 72712 434330 72740 436047
rect 73356 434330 73384 441586
rect 73988 438932 74040 438938
rect 73988 438874 74040 438880
rect 74000 434790 74028 438874
rect 74724 438864 74776 438870
rect 74724 438806 74776 438812
rect 73988 434784 74040 434790
rect 73988 434726 74040 434732
rect 74000 434330 74028 434726
rect 72712 434302 73048 434330
rect 73356 434302 73784 434330
rect 74000 434302 74336 434330
rect 74736 433673 74764 438806
rect 75196 436218 75224 460906
rect 75368 455388 75420 455394
rect 75368 455330 75420 455336
rect 75380 454170 75408 455330
rect 75368 454164 75420 454170
rect 75368 454106 75420 454112
rect 75276 452668 75328 452674
rect 75276 452610 75328 452616
rect 75288 438938 75316 452610
rect 75380 448390 75408 454106
rect 75368 448384 75420 448390
rect 75368 448326 75420 448332
rect 75366 444952 75422 444961
rect 75366 444887 75422 444896
rect 75276 438932 75328 438938
rect 75276 438874 75328 438880
rect 75380 438870 75408 444887
rect 75932 439521 75960 539158
rect 76564 536784 76616 536790
rect 76564 536726 76616 536732
rect 76576 493338 76604 536726
rect 76564 493332 76616 493338
rect 76564 493274 76616 493280
rect 77312 486470 77340 539158
rect 77300 486464 77352 486470
rect 77300 486406 77352 486412
rect 77944 485104 77996 485110
rect 77944 485046 77996 485052
rect 77208 463004 77260 463010
rect 77208 462946 77260 462952
rect 77220 441614 77248 462946
rect 77956 445874 77984 485046
rect 78692 475454 78720 539158
rect 80072 536081 80100 539158
rect 80164 539158 80960 539186
rect 81880 539158 82216 539186
rect 82800 539158 82860 539186
rect 83720 539158 84056 539186
rect 80058 536072 80114 536081
rect 80058 536007 80114 536016
rect 80164 528554 80192 539158
rect 82188 536178 82216 539158
rect 82728 538892 82780 538898
rect 82728 538834 82780 538840
rect 82176 536172 82228 536178
rect 82176 536114 82228 536120
rect 80072 528526 80192 528554
rect 78680 475448 78732 475454
rect 78680 475390 78732 475396
rect 80072 461650 80100 528526
rect 82740 466546 82768 538834
rect 82832 469878 82860 539158
rect 84028 536217 84056 539158
rect 84212 539158 84640 539186
rect 85560 539158 85620 539186
rect 84014 536208 84070 536217
rect 84014 536143 84070 536152
rect 83464 536104 83516 536110
rect 83464 536046 83516 536052
rect 82820 469872 82872 469878
rect 82820 469814 82872 469820
rect 82728 466540 82780 466546
rect 82728 466482 82780 466488
rect 80060 461644 80112 461650
rect 80060 461586 80112 461592
rect 78680 456816 78732 456822
rect 78680 456758 78732 456764
rect 78034 455696 78090 455705
rect 78034 455631 78090 455640
rect 77300 445868 77352 445874
rect 77300 445810 77352 445816
rect 77944 445868 77996 445874
rect 77944 445810 77996 445816
rect 76944 441586 77248 441614
rect 75918 439512 75974 439521
rect 75918 439447 75974 439456
rect 75368 438864 75420 438870
rect 75368 438806 75420 438812
rect 75184 436212 75236 436218
rect 75184 436154 75236 436160
rect 75644 436212 75696 436218
rect 75644 436154 75696 436160
rect 75656 434625 75684 436154
rect 75642 434616 75698 434625
rect 75642 434551 75698 434560
rect 75656 434058 75684 434551
rect 75656 434030 75808 434058
rect 71134 433664 71190 433673
rect 71134 433599 71190 433608
rect 74722 433664 74778 433673
rect 76378 433664 76434 433673
rect 74778 433622 75072 433650
rect 74722 433599 74778 433608
rect 76944 433650 76972 441586
rect 77312 434602 77340 445810
rect 78048 436218 78076 455631
rect 78692 441614 78720 456758
rect 80060 456068 80112 456074
rect 80060 456010 80112 456016
rect 78692 441586 78904 441614
rect 78036 436212 78088 436218
rect 78036 436154 78088 436160
rect 77484 436144 77536 436150
rect 77484 436086 77536 436092
rect 77266 434574 77340 434602
rect 77266 434316 77294 434574
rect 77496 434330 77524 436086
rect 78876 434330 78904 441586
rect 80072 434602 80100 456010
rect 82740 441614 82768 466482
rect 82820 452736 82872 452742
rect 82820 452678 82872 452684
rect 82832 447846 82860 452678
rect 82820 447840 82872 447846
rect 82820 447782 82872 447788
rect 83476 447166 83504 536046
rect 84212 526454 84240 539158
rect 84200 526448 84252 526454
rect 84200 526390 84252 526396
rect 85592 468518 85620 539158
rect 85580 468512 85632 468518
rect 85580 468454 85632 468460
rect 86236 458250 86264 539582
rect 86480 539158 86724 539186
rect 86696 535566 86724 539158
rect 87156 539158 87400 539186
rect 88320 539158 88472 539186
rect 86684 535560 86736 535566
rect 86684 535502 86736 535508
rect 87156 534750 87184 539158
rect 87602 536072 87658 536081
rect 87602 536007 87658 536016
rect 87144 534744 87196 534750
rect 87144 534686 87196 534692
rect 87616 465730 87644 536007
rect 87696 535560 87748 535566
rect 87696 535502 87748 535508
rect 87708 481642 87736 535502
rect 88340 533452 88392 533458
rect 88340 533394 88392 533400
rect 87696 481636 87748 481642
rect 87696 481578 87748 481584
rect 88248 481636 88300 481642
rect 88248 481578 88300 481584
rect 88260 480962 88288 481578
rect 88248 480956 88300 480962
rect 88248 480898 88300 480904
rect 87604 465724 87656 465730
rect 87604 465666 87656 465672
rect 86868 464364 86920 464370
rect 86868 464306 86920 464312
rect 85488 458244 85540 458250
rect 85488 458186 85540 458192
rect 86224 458244 86276 458250
rect 86224 458186 86276 458192
rect 82912 447160 82964 447166
rect 82912 447102 82964 447108
rect 83464 447160 83516 447166
rect 83464 447102 83516 447108
rect 82464 441586 82768 441614
rect 82924 441614 82952 447102
rect 83464 444440 83516 444446
rect 83464 444382 83516 444388
rect 82924 441586 83136 441614
rect 81346 438288 81402 438297
rect 81346 438223 81402 438232
rect 80334 436248 80390 436257
rect 80334 436183 80390 436192
rect 80026 434574 80100 434602
rect 77496 434302 77832 434330
rect 78876 434302 79304 434330
rect 79874 433800 79930 433809
rect 80026 433786 80054 434574
rect 80348 434330 80376 436183
rect 81360 434897 81388 438223
rect 81346 434888 81402 434897
rect 81346 434823 81402 434832
rect 81360 434602 81388 434823
rect 81314 434574 81388 434602
rect 80348 434302 80592 434330
rect 81314 434316 81342 434574
rect 79930 433772 80054 433786
rect 79930 433758 80040 433772
rect 79874 433735 79930 433744
rect 76434 433622 76972 433650
rect 78218 433664 78274 433673
rect 76378 433599 76434 433608
rect 81898 433664 81954 433673
rect 78274 433622 78568 433650
rect 78218 433599 78274 433608
rect 82464 433650 82492 441586
rect 82910 439512 82966 439521
rect 82910 439447 82966 439456
rect 82924 438938 82952 439447
rect 82912 438932 82964 438938
rect 82912 438874 82964 438880
rect 82818 438152 82874 438161
rect 82818 438087 82874 438096
rect 82832 437442 82860 438087
rect 82820 437436 82872 437442
rect 82820 437378 82872 437384
rect 82924 434330 82952 438874
rect 82800 434302 82952 434330
rect 83108 434330 83136 441586
rect 83476 439550 83504 444382
rect 85500 441614 85528 458186
rect 85762 453248 85818 453257
rect 85762 453183 85818 453192
rect 85224 441586 85528 441614
rect 85776 441614 85804 453183
rect 85776 441586 85896 441614
rect 83464 439544 83516 439550
rect 83464 439486 83516 439492
rect 83924 437436 83976 437442
rect 83924 437378 83976 437384
rect 83108 434302 83536 434330
rect 83936 434058 83964 437378
rect 83936 434030 84088 434058
rect 81954 433622 82492 433650
rect 84658 433664 84714 433673
rect 81898 433599 81954 433608
rect 85224 433650 85252 441586
rect 85868 437474 85896 441586
rect 85868 437446 85988 437474
rect 85854 435296 85910 435305
rect 85854 435231 85910 435240
rect 85868 434330 85896 435231
rect 85560 434302 85896 434330
rect 85960 433673 85988 437446
rect 86880 435305 86908 464306
rect 88260 454714 88288 480898
rect 88352 472666 88380 533394
rect 88444 498846 88472 539158
rect 88904 539158 89240 539186
rect 90160 539158 90404 539186
rect 88904 533458 88932 539158
rect 90376 538218 90404 539158
rect 90364 538212 90416 538218
rect 90364 538154 90416 538160
rect 88892 533452 88944 533458
rect 88892 533394 88944 533400
rect 88432 498840 88484 498846
rect 88432 498782 88484 498788
rect 88340 472660 88392 472666
rect 88340 472602 88392 472608
rect 90376 463010 90404 538154
rect 91020 478922 91048 539786
rect 94318 539744 94374 539753
rect 94318 539679 94374 539688
rect 94332 539646 94360 539679
rect 94320 539640 94372 539646
rect 94320 539582 94372 539588
rect 91204 539158 91264 539186
rect 91848 539158 92184 539186
rect 93104 539158 93440 539186
rect 94024 539158 94544 539186
rect 91100 533452 91152 533458
rect 91100 533394 91152 533400
rect 90456 478916 90508 478922
rect 90456 478858 90508 478864
rect 91008 478916 91060 478922
rect 91008 478858 91060 478864
rect 90364 463004 90416 463010
rect 90364 462946 90416 462952
rect 88248 454708 88300 454714
rect 88248 454650 88300 454656
rect 87604 450016 87656 450022
rect 87604 449958 87656 449964
rect 87616 437442 87644 449958
rect 88432 442944 88484 442950
rect 88432 442886 88484 442892
rect 88444 442270 88472 442886
rect 88432 442264 88484 442270
rect 88432 442206 88484 442212
rect 88444 441614 88472 442206
rect 88444 441586 88656 441614
rect 88522 440328 88578 440337
rect 88522 440263 88578 440272
rect 87604 437436 87656 437442
rect 87604 437378 87656 437384
rect 87328 436484 87380 436490
rect 87328 436426 87380 436432
rect 86866 435296 86922 435305
rect 86866 435231 86922 435240
rect 86880 434897 86908 435231
rect 86866 434888 86922 434897
rect 86866 434823 86922 434832
rect 87340 434330 87368 436426
rect 88536 434330 88564 440263
rect 87032 434302 87368 434330
rect 88320 434302 88564 434330
rect 88628 434330 88656 441586
rect 90468 436490 90496 478858
rect 91112 468586 91140 533394
rect 91204 485110 91232 539158
rect 91848 533458 91876 539158
rect 93412 536081 93440 539158
rect 93950 538928 94006 538937
rect 93950 538863 94006 538872
rect 93964 538286 93992 538863
rect 93952 538280 94004 538286
rect 93952 538222 94004 538228
rect 93398 536072 93454 536081
rect 93398 536007 93454 536016
rect 91836 533452 91888 533458
rect 91836 533394 91888 533400
rect 94516 531282 94544 539158
rect 93768 531276 93820 531282
rect 93768 531218 93820 531224
rect 94504 531276 94556 531282
rect 94504 531218 94556 531224
rect 93780 529242 93808 531218
rect 93768 529236 93820 529242
rect 93768 529178 93820 529184
rect 92480 490612 92532 490618
rect 92480 490554 92532 490560
rect 91192 485104 91244 485110
rect 91192 485046 91244 485052
rect 91100 468580 91152 468586
rect 91100 468522 91152 468528
rect 92386 464400 92442 464409
rect 92386 464335 92442 464344
rect 92400 462466 92428 464335
rect 92388 462460 92440 462466
rect 92388 462402 92440 462408
rect 90456 436484 90508 436490
rect 90456 436426 90508 436432
rect 89718 436248 89774 436257
rect 89718 436183 89774 436192
rect 89732 434466 89760 436183
rect 92400 436150 92428 462402
rect 92388 436144 92440 436150
rect 92388 436086 92440 436092
rect 92492 434625 92520 490554
rect 93952 473884 94004 473890
rect 93952 473826 94004 473832
rect 92570 449984 92626 449993
rect 92570 449919 92626 449928
rect 92584 442950 92612 449919
rect 92572 442944 92624 442950
rect 92572 442886 92624 442892
rect 92478 434616 92534 434625
rect 92400 434574 92478 434602
rect 89732 434438 89806 434466
rect 88628 434302 89056 434330
rect 89778 434316 89806 434438
rect 92400 434194 92428 434574
rect 92478 434551 92534 434560
rect 93964 434330 93992 473826
rect 94516 438870 94544 531218
rect 94700 473890 94728 552191
rect 94778 543008 94834 543017
rect 94778 542943 94834 542952
rect 94688 473884 94740 473890
rect 94688 473826 94740 473832
rect 94700 473414 94728 473826
rect 94688 473408 94740 473414
rect 94688 473350 94740 473356
rect 94792 449954 94820 542943
rect 95252 464370 95280 574767
rect 95896 573374 95924 580450
rect 95988 574802 96016 582354
rect 95976 574796 96028 574802
rect 95976 574738 96028 574744
rect 95884 573368 95936 573374
rect 95884 573310 95936 573316
rect 95606 567216 95662 567225
rect 95606 567151 95662 567160
rect 95422 563680 95478 563689
rect 95422 563615 95478 563624
rect 95332 536172 95384 536178
rect 95332 536114 95384 536120
rect 95240 464364 95292 464370
rect 95240 464306 95292 464312
rect 95240 458312 95292 458318
rect 95240 458254 95292 458260
rect 94780 449948 94832 449954
rect 94780 449890 94832 449896
rect 95148 449948 95200 449954
rect 95148 449890 95200 449896
rect 95160 447846 95188 449890
rect 95148 447840 95200 447846
rect 95148 447782 95200 447788
rect 95146 446448 95202 446457
rect 95146 446383 95202 446392
rect 95160 445738 95188 446383
rect 95148 445732 95200 445738
rect 95148 445674 95200 445680
rect 94504 438864 94556 438870
rect 94504 438806 94556 438812
rect 94228 436144 94280 436150
rect 94228 436086 94280 436092
rect 93840 434302 93992 434330
rect 94240 434330 94268 436086
rect 95252 434602 95280 458254
rect 95344 443018 95372 536114
rect 95436 523705 95464 563615
rect 95514 558648 95570 558657
rect 95514 558583 95570 558592
rect 95528 538898 95556 558583
rect 95516 538892 95568 538898
rect 95516 538834 95568 538840
rect 95620 534721 95648 567151
rect 96632 552537 96660 702646
rect 96712 587172 96764 587178
rect 96712 587114 96764 587120
rect 96724 568721 96752 587114
rect 98644 583840 98696 583846
rect 98644 583782 98696 583788
rect 97170 578912 97226 578921
rect 97170 578847 97226 578856
rect 97184 578270 97212 578847
rect 97172 578264 97224 578270
rect 97172 578206 97224 578212
rect 97170 577552 97226 577561
rect 97170 577487 97226 577496
rect 97184 576910 97212 577487
rect 97172 576904 97224 576910
rect 97172 576846 97224 576852
rect 97906 576464 97962 576473
rect 97906 576399 97962 576408
rect 97920 576162 97948 576399
rect 97908 576156 97960 576162
rect 97908 576098 97960 576104
rect 97906 573472 97962 573481
rect 97962 573430 98040 573458
rect 97906 573407 97962 573416
rect 96802 572112 96858 572121
rect 96802 572047 96858 572056
rect 96816 571402 96844 572047
rect 97262 571432 97318 571441
rect 96804 571396 96856 571402
rect 97262 571367 97318 571376
rect 96804 571338 96856 571344
rect 96710 568712 96766 568721
rect 96710 568647 96766 568656
rect 97276 565865 97304 571367
rect 97906 570072 97962 570081
rect 97906 570007 97962 570016
rect 97920 569974 97948 570007
rect 97908 569968 97960 569974
rect 97908 569910 97960 569916
rect 97906 568712 97962 568721
rect 97906 568647 97908 568656
rect 97960 568647 97962 568656
rect 97908 568618 97960 568624
rect 96710 565856 96766 565865
rect 96710 565791 96766 565800
rect 97262 565856 97318 565865
rect 97262 565791 97318 565800
rect 96618 552528 96674 552537
rect 96618 552463 96674 552472
rect 96724 539850 96752 565791
rect 96802 562320 96858 562329
rect 96802 562255 96858 562264
rect 96816 561746 96844 562255
rect 96804 561740 96856 561746
rect 96804 561682 96856 561688
rect 96894 560960 96950 560969
rect 96894 560895 96950 560904
rect 96802 559600 96858 559609
rect 96802 559535 96858 559544
rect 96816 558958 96844 559535
rect 96804 558952 96856 558958
rect 96804 558894 96856 558900
rect 96802 556880 96858 556889
rect 96802 556815 96858 556824
rect 96712 539844 96764 539850
rect 96712 539786 96764 539792
rect 95606 534712 95662 534721
rect 95606 534647 95662 534656
rect 96816 533390 96844 556815
rect 96908 537538 96936 560895
rect 96986 555520 97042 555529
rect 96986 555455 97042 555464
rect 97000 554810 97028 555455
rect 96988 554804 97040 554810
rect 96988 554746 97040 554752
rect 96986 552800 97042 552809
rect 96986 552735 97042 552744
rect 97000 552090 97028 552735
rect 96988 552084 97040 552090
rect 96988 552026 97040 552032
rect 97906 550760 97962 550769
rect 97906 550695 97962 550704
rect 97920 550662 97948 550695
rect 97908 550656 97960 550662
rect 97908 550598 97960 550604
rect 96986 545728 97042 545737
rect 96986 545663 97042 545672
rect 96896 537532 96948 537538
rect 96896 537474 96948 537480
rect 96804 533384 96856 533390
rect 96804 533326 96856 533332
rect 95422 523696 95478 523705
rect 95422 523631 95478 523640
rect 97000 479534 97028 545663
rect 97078 544368 97134 544377
rect 97078 544303 97134 544312
rect 97092 543794 97120 544303
rect 97080 543788 97132 543794
rect 97080 543730 97132 543736
rect 97170 541648 97226 541657
rect 97170 541583 97226 541592
rect 97184 541006 97212 541583
rect 97172 541000 97224 541006
rect 97172 540942 97224 540948
rect 98012 518226 98040 573430
rect 98000 518220 98052 518226
rect 98000 518162 98052 518168
rect 96988 479528 97040 479534
rect 96988 479470 97040 479476
rect 98656 475386 98684 583782
rect 100208 582548 100260 582554
rect 100208 582490 100260 582496
rect 99380 487824 99432 487830
rect 99380 487766 99432 487772
rect 98736 475448 98788 475454
rect 98736 475390 98788 475396
rect 98644 475380 98696 475386
rect 98644 475322 98696 475328
rect 96618 456104 96674 456113
rect 96618 456039 96674 456048
rect 95332 443012 95384 443018
rect 95332 442954 95384 442960
rect 95344 440881 95372 442954
rect 95330 440872 95386 440881
rect 95330 440807 95386 440816
rect 96632 437474 96660 456039
rect 98644 449948 98696 449954
rect 98644 449890 98696 449896
rect 97356 438864 97408 438870
rect 97356 438806 97408 438812
rect 96632 437446 96752 437474
rect 95252 434574 95326 434602
rect 94240 434302 94576 434330
rect 95298 434316 95326 434574
rect 92400 434166 92552 434194
rect 96724 433809 96752 437446
rect 97368 437442 97396 438806
rect 98656 437442 98684 449890
rect 98748 437442 98776 475390
rect 97356 437436 97408 437442
rect 97356 437378 97408 437384
rect 98644 437436 98696 437442
rect 98644 437378 98696 437384
rect 98736 437436 98788 437442
rect 98736 437378 98788 437384
rect 97368 434602 97396 437378
rect 99392 436529 99420 487766
rect 99378 436520 99434 436529
rect 99378 436455 99434 436464
rect 99746 436520 99802 436529
rect 99746 436455 99802 436464
rect 97322 434574 97396 434602
rect 97322 434316 97350 434574
rect 99760 434330 99788 436455
rect 99760 434302 100096 434330
rect 100220 434042 100248 582490
rect 102784 580304 102836 580310
rect 102784 580246 102836 580252
rect 102796 487830 102824 580246
rect 104820 576162 104848 702918
rect 104912 625870 104940 703582
rect 105280 703474 105308 703582
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 136652 703582 137692 703610
rect 105464 703474 105492 703520
rect 105280 703446 105492 703474
rect 104900 625864 104952 625870
rect 104900 625806 104952 625812
rect 112444 592068 112496 592074
rect 112444 592010 112496 592016
rect 107014 582584 107070 582593
rect 107014 582519 107070 582528
rect 104808 576156 104860 576162
rect 104808 576098 104860 576104
rect 104164 574796 104216 574802
rect 104164 574738 104216 574744
rect 102876 493332 102928 493338
rect 102876 493274 102928 493280
rect 102140 487824 102192 487830
rect 102140 487766 102192 487772
rect 102784 487824 102836 487830
rect 102784 487766 102836 487772
rect 101218 436384 101274 436393
rect 101218 436319 101274 436328
rect 101232 434330 101260 436319
rect 102152 434330 102180 487766
rect 102888 466478 102916 493274
rect 104176 476134 104204 574738
rect 106924 571396 106976 571402
rect 106924 571338 106976 571344
rect 104440 568676 104492 568682
rect 104440 568618 104492 568624
rect 104348 543788 104400 543794
rect 104348 543730 104400 543736
rect 104254 536208 104310 536217
rect 104254 536143 104310 536152
rect 104164 476128 104216 476134
rect 104164 476070 104216 476076
rect 102416 466472 102468 466478
rect 102416 466414 102468 466420
rect 102876 466472 102928 466478
rect 102876 466414 102928 466420
rect 102428 441614 102456 466414
rect 102428 441586 102640 441614
rect 104176 441590 104204 476070
rect 104268 475250 104296 536143
rect 104360 521626 104388 543730
rect 104452 535537 104480 568618
rect 104438 535528 104494 535537
rect 104438 535463 104494 535472
rect 104348 521620 104400 521626
rect 104348 521562 104400 521568
rect 106936 478174 106964 571338
rect 107028 562970 107056 582519
rect 108304 581120 108356 581126
rect 108304 581062 108356 581068
rect 107016 562964 107068 562970
rect 107016 562906 107068 562912
rect 107016 532024 107068 532030
rect 107016 531966 107068 531972
rect 106924 478168 106976 478174
rect 106924 478110 106976 478116
rect 104256 475244 104308 475250
rect 104256 475186 104308 475192
rect 104808 475244 104860 475250
rect 104808 475186 104860 475192
rect 104820 474774 104848 475186
rect 104808 474768 104860 474774
rect 104808 474710 104860 474716
rect 104256 451376 104308 451382
rect 104256 451318 104308 451324
rect 102612 434330 102640 441586
rect 104164 441584 104216 441590
rect 104164 441526 104216 441532
rect 103704 437436 103756 437442
rect 103704 437378 103756 437384
rect 101232 434302 101568 434330
rect 102152 434302 102304 434330
rect 102612 434302 103040 434330
rect 103716 434058 103744 437378
rect 104176 434330 104204 441526
rect 104268 437442 104296 451318
rect 104820 439550 104848 474710
rect 107028 467945 107056 531966
rect 107014 467936 107070 467945
rect 107014 467871 107070 467880
rect 107566 467936 107622 467945
rect 107566 467871 107622 467880
rect 104900 454708 104952 454714
rect 104900 454650 104952 454656
rect 104912 441614 104940 454650
rect 106924 449200 106976 449206
rect 106924 449142 106976 449148
rect 106936 441614 106964 449142
rect 104912 441586 105400 441614
rect 104808 439544 104860 439550
rect 104808 439486 104860 439492
rect 104256 437436 104308 437442
rect 104256 437378 104308 437384
rect 105372 434330 105400 441586
rect 106660 441586 106964 441614
rect 106660 437073 106688 441586
rect 106646 437064 106702 437073
rect 106646 436999 106702 437008
rect 106660 434330 106688 436999
rect 107384 436756 107436 436762
rect 107384 436698 107436 436704
rect 104176 434302 104328 434330
rect 105372 434302 105800 434330
rect 106352 434302 106688 434330
rect 100208 434036 100260 434042
rect 103592 434030 103744 434058
rect 100208 433978 100260 433984
rect 91466 433800 91522 433809
rect 96710 433800 96766 433809
rect 91522 433758 91816 433786
rect 91466 433735 91522 433744
rect 96710 433735 96766 433744
rect 100482 433800 100538 433809
rect 100538 433758 100832 433786
rect 100482 433735 100538 433744
rect 84714 433622 85252 433650
rect 85946 433664 86002 433673
rect 84658 433599 84714 433608
rect 87234 433664 87290 433673
rect 86002 433622 86296 433650
rect 85946 433599 86002 433608
rect 89994 433664 90050 433673
rect 87290 433622 87584 433650
rect 87234 433599 87290 433608
rect 91190 433664 91246 433673
rect 90050 433622 90344 433650
rect 91080 433622 91190 433650
rect 89994 433599 90050 433608
rect 91190 433599 91246 433608
rect 92938 433664 92994 433673
rect 96342 433664 96398 433673
rect 92994 433622 93288 433650
rect 96048 433622 96342 433650
rect 92938 433599 92994 433608
rect 96724 433650 96752 433735
rect 98182 433664 98238 433673
rect 96600 433622 96752 433650
rect 98072 433622 98182 433650
rect 96342 433599 96398 433608
rect 98182 433599 98238 433608
rect 98458 433664 98514 433673
rect 99838 433664 99894 433673
rect 98514 433622 98808 433650
rect 99544 433622 99838 433650
rect 98458 433599 98514 433608
rect 99838 433599 99894 433608
rect 104714 433664 104770 433673
rect 106738 433664 106794 433673
rect 104770 433622 105064 433650
rect 104714 433599 104770 433608
rect 107396 433650 107424 436698
rect 107580 435470 107608 467871
rect 108316 437442 108344 581062
rect 111064 562964 111116 562970
rect 111064 562906 111116 562912
rect 108488 552084 108540 552090
rect 108488 552026 108540 552032
rect 108396 521620 108448 521626
rect 108396 521562 108448 521568
rect 108408 467906 108436 521562
rect 108500 507006 108528 552026
rect 108488 507000 108540 507006
rect 108488 506942 108540 506948
rect 108488 486464 108540 486470
rect 108488 486406 108540 486412
rect 108500 471306 108528 486406
rect 108488 471300 108540 471306
rect 108488 471242 108540 471248
rect 109684 469872 109736 469878
rect 109684 469814 109736 469820
rect 108396 467900 108448 467906
rect 108396 467842 108448 467848
rect 108304 437436 108356 437442
rect 108304 437378 108356 437384
rect 107658 436112 107714 436121
rect 107658 436047 107714 436056
rect 107568 435464 107620 435470
rect 107568 435406 107620 435412
rect 107672 434330 107700 436047
rect 108316 434330 108344 437378
rect 108408 436121 108436 467842
rect 109696 437345 109724 469814
rect 111076 449177 111104 562906
rect 112456 483682 112484 592010
rect 124404 589348 124456 589354
rect 124404 589290 124456 589296
rect 121460 585812 121512 585818
rect 121460 585754 121512 585760
rect 121472 585274 121500 585754
rect 121460 585268 121512 585274
rect 121460 585210 121512 585216
rect 116584 585200 116636 585206
rect 116584 585142 116636 585148
rect 115204 583772 115256 583778
rect 115204 583714 115256 583720
rect 112720 558952 112772 558958
rect 112720 558894 112772 558900
rect 112536 507000 112588 507006
rect 112536 506942 112588 506948
rect 112444 483676 112496 483682
rect 112444 483618 112496 483624
rect 112548 470594 112576 506942
rect 112456 470566 112576 470594
rect 112456 469266 112484 470566
rect 112444 469260 112496 469266
rect 112444 469202 112496 469208
rect 112456 452606 112484 469202
rect 111800 452600 111852 452606
rect 111800 452542 111852 452548
rect 112444 452600 112496 452606
rect 112444 452542 112496 452548
rect 111812 451314 111840 452542
rect 111800 451308 111852 451314
rect 111800 451250 111852 451256
rect 111062 449168 111118 449177
rect 111062 449103 111118 449112
rect 111076 448633 111104 449103
rect 110418 448624 110474 448633
rect 110418 448559 110474 448568
rect 111062 448624 111118 448633
rect 111062 448559 111118 448568
rect 110432 441614 110460 448559
rect 111812 441614 111840 451250
rect 110432 441586 110920 441614
rect 111812 441586 112208 441614
rect 109682 437336 109738 437345
rect 109682 437271 109738 437280
rect 108394 436112 108450 436121
rect 108394 436047 108450 436056
rect 109696 434330 109724 437271
rect 110892 434330 110920 441586
rect 112180 434330 112208 441586
rect 107672 434302 107824 434330
rect 108316 434302 108560 434330
rect 109696 434302 109848 434330
rect 110892 434302 111320 434330
rect 112180 434302 112608 434330
rect 106794 433622 107424 433650
rect 109038 433664 109094 433673
rect 106738 433599 106794 433608
rect 110694 433664 110750 433673
rect 109094 433622 109296 433650
rect 110584 433622 110694 433650
rect 109038 433599 109094 433608
rect 110694 433599 110750 433608
rect 111798 433664 111854 433673
rect 111854 433622 112056 433650
rect 111798 433599 111854 433608
rect 68652 433288 68704 433294
rect 68652 433230 68704 433236
rect 68664 433129 68692 433230
rect 68650 433120 68706 433129
rect 68650 433055 68706 433064
rect 68572 431926 68692 431954
rect 67822 429856 67878 429865
rect 67822 429791 67878 429800
rect 67732 397520 67784 397526
rect 67730 397488 67732 397497
rect 67784 397488 67786 397497
rect 67786 397446 67864 397474
rect 67730 397423 67786 397432
rect 67744 397397 67772 397423
rect 67730 396400 67786 396409
rect 67730 396335 67786 396344
rect 67546 392048 67602 392057
rect 67546 391983 67602 391992
rect 67546 391232 67602 391241
rect 67546 391167 67602 391176
rect 67560 387433 67588 391167
rect 67640 390176 67692 390182
rect 67640 390118 67692 390124
rect 67546 387424 67602 387433
rect 67546 387359 67602 387368
rect 67652 368422 67680 390118
rect 67744 383042 67772 396335
rect 67836 386374 67864 397446
rect 67824 386368 67876 386374
rect 67824 386310 67876 386316
rect 67732 383036 67784 383042
rect 67732 382978 67784 382984
rect 67640 368416 67692 368422
rect 67640 368358 67692 368364
rect 67456 314696 67508 314702
rect 67456 314638 67508 314644
rect 67364 288448 67416 288454
rect 67364 288390 67416 288396
rect 67086 283792 67142 283801
rect 67086 283727 67142 283736
rect 66812 283008 66864 283014
rect 66810 282976 66812 282985
rect 66864 282976 66866 282985
rect 66810 282911 66866 282920
rect 66168 282260 66220 282266
rect 66168 282202 66220 282208
rect 67100 282198 67128 283727
rect 67088 282192 67140 282198
rect 67086 282160 67088 282169
rect 67272 282192 67324 282198
rect 67140 282160 67142 282169
rect 67272 282134 67324 282140
rect 67086 282095 67142 282104
rect 67284 281625 67312 282134
rect 67270 281616 67326 281625
rect 67270 281551 67326 281560
rect 66534 281480 66590 281489
rect 66534 281415 66590 281424
rect 66548 280226 66576 281415
rect 66902 280528 66958 280537
rect 66902 280463 66958 280472
rect 66916 280294 66944 280463
rect 66904 280288 66956 280294
rect 66904 280230 66956 280236
rect 66536 280220 66588 280226
rect 66536 280162 66588 280168
rect 67180 280220 67232 280226
rect 67180 280162 67232 280168
rect 66628 279472 66680 279478
rect 66628 279414 66680 279420
rect 66640 278905 66668 279414
rect 66626 278896 66682 278905
rect 66626 278831 66682 278840
rect 66810 278080 66866 278089
rect 66810 278015 66812 278024
rect 66864 278015 66866 278024
rect 66812 277986 66864 277992
rect 66088 277366 66208 277394
rect 66180 275641 66208 277366
rect 66904 277364 66956 277370
rect 66904 277306 66956 277312
rect 66916 276457 66944 277306
rect 66902 276448 66958 276457
rect 66902 276383 66958 276392
rect 66166 275632 66222 275641
rect 66166 275567 66222 275576
rect 66074 274816 66130 274825
rect 66074 274751 66130 274760
rect 65982 239864 66038 239873
rect 65982 239799 66038 239808
rect 65904 229066 66024 229094
rect 65800 227044 65852 227050
rect 65800 226986 65852 226992
rect 65812 226409 65840 226986
rect 65798 226400 65854 226409
rect 65798 226335 65854 226344
rect 65812 144945 65840 226335
rect 65996 225622 66024 229066
rect 65984 225616 66036 225622
rect 65984 225558 66036 225564
rect 65798 144936 65854 144945
rect 65798 144871 65854 144880
rect 65812 142154 65840 144871
rect 65812 142126 65932 142154
rect 64788 140072 64840 140078
rect 64788 140014 64840 140020
rect 64694 139632 64750 139641
rect 64694 139567 64750 139576
rect 64708 132394 64736 139567
rect 64696 132388 64748 132394
rect 64696 132330 64748 132336
rect 64604 128308 64656 128314
rect 64604 128250 64656 128256
rect 64512 110424 64564 110430
rect 64512 110366 64564 110372
rect 63408 103488 63460 103494
rect 63408 103430 63460 103436
rect 64604 99476 64656 99482
rect 64604 99418 64656 99424
rect 63316 90976 63368 90982
rect 63316 90918 63368 90924
rect 64616 89593 64644 99418
rect 64696 95260 64748 95266
rect 64696 95202 64748 95208
rect 64602 89584 64658 89593
rect 64602 89519 64658 89528
rect 63224 88324 63276 88330
rect 63224 88266 63276 88272
rect 64708 69018 64736 95202
rect 64800 92410 64828 140014
rect 65524 109064 65576 109070
rect 65524 109006 65576 109012
rect 64788 92404 64840 92410
rect 64788 92346 64840 92352
rect 65536 85542 65564 109006
rect 65904 107817 65932 142126
rect 65996 110265 66024 225558
rect 66088 136678 66116 274751
rect 66534 274000 66590 274009
rect 66534 273935 66536 273944
rect 66588 273935 66590 273944
rect 66536 273906 66588 273912
rect 66626 272368 66682 272377
rect 66626 272303 66682 272312
rect 66640 271930 66668 272303
rect 66628 271924 66680 271930
rect 66628 271866 66680 271872
rect 66258 271552 66314 271561
rect 66258 271487 66314 271496
rect 66272 270570 66300 271487
rect 66260 270564 66312 270570
rect 66260 270506 66312 270512
rect 66902 269104 66958 269113
rect 66902 269039 66958 269048
rect 66916 268462 66944 269039
rect 66904 268456 66956 268462
rect 66904 268398 66956 268404
rect 66812 268388 66864 268394
rect 66812 268330 66864 268336
rect 66824 268297 66852 268330
rect 66810 268288 66866 268297
rect 66810 268223 66866 268232
rect 66626 267472 66682 267481
rect 66626 267407 66682 267416
rect 66640 267034 66668 267407
rect 66628 267028 66680 267034
rect 66628 266970 66680 266976
rect 66442 266656 66498 266665
rect 66442 266591 66498 266600
rect 66456 266422 66484 266591
rect 66444 266416 66496 266422
rect 66444 266358 66496 266364
rect 66810 265840 66866 265849
rect 66810 265775 66866 265784
rect 66824 264994 66852 265775
rect 66812 264988 66864 264994
rect 66812 264930 66864 264936
rect 66260 264240 66312 264246
rect 66260 264182 66312 264188
rect 66810 264208 66866 264217
rect 66272 261769 66300 264182
rect 66810 264143 66866 264152
rect 66824 263634 66852 264143
rect 66812 263628 66864 263634
rect 66812 263570 66864 263576
rect 67086 263392 67142 263401
rect 67086 263327 67142 263336
rect 67100 262886 67128 263327
rect 67088 262880 67140 262886
rect 67088 262822 67140 262828
rect 66902 262576 66958 262585
rect 66902 262511 66958 262520
rect 66258 261760 66314 261769
rect 66258 261695 66314 261704
rect 66272 260166 66300 261695
rect 66916 260914 66944 262511
rect 66904 260908 66956 260914
rect 66904 260850 66956 260856
rect 66260 260160 66312 260166
rect 66260 260102 66312 260108
rect 66810 260128 66866 260137
rect 66810 260063 66866 260072
rect 66444 258732 66496 258738
rect 66444 258674 66496 258680
rect 66456 258058 66484 258674
rect 66824 258505 66852 260063
rect 66810 258496 66866 258505
rect 66810 258431 66866 258440
rect 66260 258052 66312 258058
rect 66260 257994 66312 258000
rect 66444 258052 66496 258058
rect 66444 257994 66496 258000
rect 66272 257961 66300 257994
rect 66258 257952 66314 257961
rect 66258 257887 66314 257896
rect 66628 256896 66680 256902
rect 66626 256864 66628 256873
rect 66680 256864 66682 256873
rect 66626 256799 66682 256808
rect 66812 254584 66864 254590
rect 66812 254526 66864 254532
rect 66824 254425 66852 254526
rect 66810 254416 66866 254425
rect 66810 254351 66866 254360
rect 66916 252550 66944 260850
rect 66994 253600 67050 253609
rect 66994 253535 67050 253544
rect 67008 253230 67036 253535
rect 66996 253224 67048 253230
rect 66996 253166 67048 253172
rect 66904 252544 66956 252550
rect 66904 252486 66956 252492
rect 66810 251968 66866 251977
rect 66810 251903 66866 251912
rect 66824 251870 66852 251903
rect 66812 251864 66864 251870
rect 66812 251806 66864 251812
rect 66812 251184 66864 251190
rect 66442 251152 66498 251161
rect 66812 251126 66864 251132
rect 66442 251087 66498 251096
rect 66456 249830 66484 251087
rect 66824 250345 66852 251126
rect 66810 250336 66866 250345
rect 66810 250271 66866 250280
rect 66444 249824 66496 249830
rect 66444 249766 66496 249772
rect 66626 249520 66682 249529
rect 66626 249455 66682 249464
rect 66640 249082 66668 249455
rect 66628 249076 66680 249082
rect 66628 249018 66680 249024
rect 66166 248704 66222 248713
rect 66166 248639 66222 248648
rect 66076 136672 66128 136678
rect 66076 136614 66128 136620
rect 66088 123865 66116 136614
rect 66074 123856 66130 123865
rect 66074 123791 66130 123800
rect 65982 110256 66038 110265
rect 65982 110191 66038 110200
rect 65996 109070 66024 110191
rect 65984 109064 66036 109070
rect 65984 109006 66036 109012
rect 65890 107808 65946 107817
rect 65890 107743 65946 107752
rect 66076 105596 66128 105602
rect 66076 105538 66128 105544
rect 65984 101448 66036 101454
rect 65984 101390 66036 101396
rect 65524 85536 65576 85542
rect 65524 85478 65576 85484
rect 65996 82822 66024 101390
rect 66088 85513 66116 105538
rect 66180 99634 66208 248639
rect 66812 245608 66864 245614
rect 66812 245550 66864 245556
rect 66824 244633 66852 245550
rect 66810 244624 66866 244633
rect 66810 244559 66866 244568
rect 66812 244248 66864 244254
rect 66812 244190 66864 244196
rect 66626 243808 66682 243817
rect 66626 243743 66682 243752
rect 66640 242962 66668 243743
rect 66824 243001 66852 244190
rect 66810 242992 66866 243001
rect 66628 242956 66680 242962
rect 66810 242927 66866 242936
rect 66628 242898 66680 242904
rect 66260 132456 66312 132462
rect 66260 132398 66312 132404
rect 66272 132025 66300 132398
rect 66352 132388 66404 132394
rect 66352 132330 66404 132336
rect 66258 132016 66314 132025
rect 66258 131951 66314 131960
rect 66364 131209 66392 132330
rect 66350 131200 66406 131209
rect 66350 131135 66406 131144
rect 66260 131096 66312 131102
rect 66260 131038 66312 131044
rect 66272 130665 66300 131038
rect 66258 130656 66314 130665
rect 66258 130591 66314 130600
rect 67192 129849 67220 280162
rect 67376 277273 67404 288390
rect 67362 277264 67418 277273
rect 67362 277199 67418 277208
rect 67468 263401 67496 314638
rect 67548 298784 67600 298790
rect 67548 298726 67600 298732
rect 67560 283801 67588 298726
rect 67546 283792 67602 283801
rect 67546 283727 67602 283736
rect 67548 283076 67600 283082
rect 67548 283018 67600 283024
rect 67560 279721 67588 283018
rect 67546 279712 67602 279721
rect 67546 279647 67602 279656
rect 67454 263392 67510 263401
rect 67454 263327 67510 263336
rect 67272 253224 67324 253230
rect 67272 253166 67324 253172
rect 67284 230450 67312 253166
rect 67454 247072 67510 247081
rect 67454 247007 67510 247016
rect 67362 246256 67418 246265
rect 67362 246191 67418 246200
rect 67272 230444 67324 230450
rect 67272 230386 67324 230392
rect 67284 135318 67312 230386
rect 67376 222154 67404 246191
rect 67468 234598 67496 247007
rect 67652 242962 67680 368358
rect 68664 326398 68692 431926
rect 112732 407017 112760 558894
rect 113180 525088 113232 525094
rect 113180 525030 113232 525036
rect 113192 414905 113220 525030
rect 113364 468512 113416 468518
rect 113364 468454 113416 468460
rect 113272 461644 113324 461650
rect 113272 461586 113324 461592
rect 113284 436801 113312 461586
rect 113270 436792 113326 436801
rect 113270 436727 113326 436736
rect 113270 416800 113326 416809
rect 113270 416735 113326 416744
rect 113178 414896 113234 414905
rect 113178 414831 113234 414840
rect 112718 407008 112774 407017
rect 112718 406943 112774 406952
rect 112718 401840 112774 401849
rect 112718 401775 112774 401784
rect 72514 390960 72570 390969
rect 72514 390895 72570 390904
rect 73986 390960 74042 390969
rect 76654 390960 76710 390969
rect 74042 390918 74488 390946
rect 76360 390918 76654 390946
rect 73986 390895 74042 390904
rect 71134 390824 71190 390833
rect 70688 390782 71134 390810
rect 69664 390584 69716 390590
rect 69368 390532 69664 390538
rect 69368 390526 69716 390532
rect 69368 390510 69704 390526
rect 68802 390182 68830 390388
rect 69584 390374 70104 390402
rect 68790 390176 68842 390182
rect 68790 390118 68842 390124
rect 69584 373994 69612 390374
rect 70688 388249 70716 390782
rect 71134 390759 71190 390768
rect 71240 390374 71576 390402
rect 72128 390374 72464 390402
rect 70674 388240 70730 388249
rect 70674 388175 70730 388184
rect 71240 387841 71268 390374
rect 71688 389156 71740 389162
rect 71688 389098 71740 389104
rect 71226 387832 71282 387841
rect 71226 387767 71282 387776
rect 69662 383752 69718 383761
rect 69662 383687 69718 383696
rect 69032 373966 69612 373994
rect 69032 361554 69060 373966
rect 69020 361548 69072 361554
rect 69020 361490 69072 361496
rect 69032 360534 69060 361490
rect 69020 360528 69072 360534
rect 69020 360470 69072 360476
rect 68652 326392 68704 326398
rect 68652 326334 68704 326340
rect 68664 316034 68692 326334
rect 68296 316006 68692 316034
rect 68296 281489 68324 316006
rect 68652 287768 68704 287774
rect 68652 287710 68704 287716
rect 68558 283520 68614 283529
rect 68558 283455 68614 283464
rect 68282 281480 68338 281489
rect 68282 281415 68338 281424
rect 68190 258768 68246 258777
rect 68190 258703 68246 258712
rect 68204 258058 68232 258703
rect 68192 258052 68244 258058
rect 68192 257994 68244 258000
rect 68284 252544 68336 252550
rect 68284 252486 68336 252492
rect 67640 242956 67692 242962
rect 67640 242898 67692 242904
rect 67456 234592 67508 234598
rect 67456 234534 67508 234540
rect 67364 222148 67416 222154
rect 67364 222090 67416 222096
rect 67272 135312 67324 135318
rect 67272 135254 67324 135260
rect 67178 129840 67234 129849
rect 67178 129775 67234 129784
rect 66258 129024 66314 129033
rect 66258 128959 66314 128968
rect 66272 128722 66300 128959
rect 66260 128716 66312 128722
rect 66260 128658 66312 128664
rect 66904 128308 66956 128314
rect 66904 128250 66956 128256
rect 66916 127673 66944 128250
rect 66902 127664 66958 127673
rect 66902 127599 66958 127608
rect 66904 126948 66956 126954
rect 66904 126890 66956 126896
rect 66812 126880 66864 126886
rect 66810 126848 66812 126857
rect 66864 126848 66866 126857
rect 66810 126783 66866 126792
rect 66916 126041 66944 126890
rect 66902 126032 66958 126041
rect 66902 125967 66958 125976
rect 66812 125384 66864 125390
rect 66812 125326 66864 125332
rect 66824 125225 66852 125326
rect 66810 125216 66866 125225
rect 66810 125151 66866 125160
rect 66812 124908 66864 124914
rect 66812 124850 66864 124856
rect 66824 123049 66852 124850
rect 66810 123040 66866 123049
rect 66810 122975 66866 122984
rect 66352 122800 66404 122806
rect 66352 122742 66404 122748
rect 66364 122233 66392 122742
rect 66350 122224 66406 122233
rect 66350 122159 66406 122168
rect 66812 121440 66864 121446
rect 66810 121408 66812 121417
rect 66864 121408 66866 121417
rect 66810 121343 66866 121352
rect 66904 121372 66956 121378
rect 66904 121314 66956 121320
rect 66916 120601 66944 121314
rect 66902 120592 66958 120601
rect 66902 120527 66958 120536
rect 66812 120080 66864 120086
rect 66810 120048 66812 120057
rect 66864 120048 66866 120057
rect 66810 119983 66866 119992
rect 66904 120012 66956 120018
rect 66904 119954 66956 119960
rect 66916 119241 66944 119954
rect 66902 119232 66958 119241
rect 66902 119167 66958 119176
rect 66812 118652 66864 118658
rect 66812 118594 66864 118600
rect 66824 117609 66852 118594
rect 66904 118584 66956 118590
rect 66904 118526 66956 118532
rect 66916 118425 66944 118526
rect 66902 118416 66958 118425
rect 66902 118351 66958 118360
rect 66810 117600 66866 117609
rect 66810 117535 66866 117544
rect 66628 117292 66680 117298
rect 66628 117234 66680 117240
rect 66640 116249 66668 117234
rect 66626 116240 66682 116249
rect 66626 116175 66682 116184
rect 66812 115932 66864 115938
rect 66812 115874 66864 115880
rect 66824 115433 66852 115874
rect 66904 115456 66956 115462
rect 66810 115424 66866 115433
rect 66904 115398 66956 115404
rect 66810 115359 66866 115368
rect 66916 114617 66944 115398
rect 66902 114608 66958 114617
rect 66902 114543 66958 114552
rect 66812 114504 66864 114510
rect 66812 114446 66864 114452
rect 66824 113801 66852 114446
rect 66904 113824 66956 113830
rect 66810 113792 66866 113801
rect 66904 113766 66956 113772
rect 66810 113727 66866 113736
rect 66916 113257 66944 113766
rect 66902 113248 66958 113257
rect 66902 113183 66958 113192
rect 67180 112464 67232 112470
rect 67180 112406 67232 112412
rect 66904 111784 66956 111790
rect 66904 111726 66956 111732
rect 66916 111625 66944 111726
rect 66902 111616 66958 111625
rect 66902 111551 66958 111560
rect 67192 110809 67220 112406
rect 67178 110800 67234 110809
rect 67178 110735 67234 110744
rect 66812 110424 66864 110430
rect 66812 110366 66864 110372
rect 66824 109449 66852 110366
rect 66810 109440 66866 109449
rect 66810 109375 66866 109384
rect 66810 106992 66866 107001
rect 66810 106927 66866 106936
rect 66824 106350 66852 106927
rect 66812 106344 66864 106350
rect 66812 106286 66864 106292
rect 66626 105632 66682 105641
rect 66626 105567 66628 105576
rect 66680 105567 66682 105576
rect 66628 105538 66680 105544
rect 66812 104848 66864 104854
rect 66810 104816 66812 104825
rect 66864 104816 66866 104825
rect 66810 104751 66866 104760
rect 67284 104009 67312 135254
rect 67270 104000 67326 104009
rect 67270 103935 67326 103944
rect 66812 102808 66864 102814
rect 66812 102750 66864 102756
rect 66824 102649 66852 102750
rect 66810 102640 66866 102649
rect 66810 102575 66866 102584
rect 66534 101824 66590 101833
rect 66534 101759 66590 101768
rect 66548 101454 66576 101759
rect 66536 101448 66588 101454
rect 66536 101390 66588 101396
rect 66810 101008 66866 101017
rect 66810 100943 66866 100952
rect 66824 100774 66852 100943
rect 66812 100768 66864 100774
rect 66812 100710 66864 100716
rect 66718 100192 66774 100201
rect 66718 100127 66774 100136
rect 66258 99648 66314 99657
rect 66180 99606 66258 99634
rect 66074 85504 66130 85513
rect 66074 85439 66130 85448
rect 65984 82816 66036 82822
rect 65984 82758 66036 82764
rect 65996 81462 66024 82758
rect 65524 81456 65576 81462
rect 65524 81398 65576 81404
rect 65984 81456 66036 81462
rect 65984 81398 66036 81404
rect 64696 69012 64748 69018
rect 64696 68954 64748 68960
rect 61844 67584 61896 67590
rect 61844 67526 61896 67532
rect 65536 45558 65564 81398
rect 66180 66162 66208 99606
rect 66258 99583 66314 99592
rect 66732 99482 66760 100127
rect 66720 99476 66772 99482
rect 66720 99418 66772 99424
rect 67376 97209 67404 222090
rect 67468 98025 67496 234534
rect 67546 149152 67602 149161
rect 67546 149087 67548 149096
rect 67600 149087 67602 149096
rect 67548 149058 67600 149064
rect 67652 103514 67680 242898
rect 68296 231130 68324 252486
rect 68284 231124 68336 231130
rect 68284 231066 68336 231072
rect 68572 169794 68600 283455
rect 68664 248414 68692 287710
rect 69676 285802 69704 383687
rect 71700 363662 71728 389098
rect 72436 389065 72464 390374
rect 72422 389056 72478 389065
rect 72422 388991 72478 389000
rect 72528 387569 72556 390895
rect 73804 390652 73856 390658
rect 73804 390594 73856 390600
rect 72620 390374 72864 390402
rect 73172 390374 73600 390402
rect 72620 389162 72648 390374
rect 72608 389156 72660 389162
rect 72608 389098 72660 389104
rect 72974 389056 73030 389065
rect 72974 388991 73030 389000
rect 72514 387560 72570 387569
rect 72514 387495 72570 387504
rect 72988 375290 73016 388991
rect 73172 387002 73200 390374
rect 73080 386974 73200 387002
rect 72976 375284 73028 375290
rect 72976 375226 73028 375232
rect 71688 363656 71740 363662
rect 71688 363598 71740 363604
rect 69756 360528 69808 360534
rect 69756 360470 69808 360476
rect 69112 285796 69164 285802
rect 69112 285738 69164 285744
rect 69664 285796 69716 285802
rect 69664 285738 69716 285744
rect 69124 283370 69152 285738
rect 69386 283520 69442 283529
rect 69442 283478 69552 283506
rect 69386 283455 69442 283464
rect 69768 283393 69796 360470
rect 73080 356697 73108 386974
rect 73816 376650 73844 390594
rect 74460 388929 74488 390918
rect 75058 390130 75086 390388
rect 75196 390374 75624 390402
rect 75058 390102 75132 390130
rect 75104 389298 75132 390102
rect 75092 389292 75144 389298
rect 75092 389234 75144 389240
rect 74446 388920 74502 388929
rect 74446 388855 74502 388864
rect 73804 376644 73856 376650
rect 73804 376586 73856 376592
rect 75196 373994 75224 390374
rect 76576 376038 76604 390918
rect 76654 390895 76710 390904
rect 95252 390782 95864 390810
rect 96600 390782 96936 390810
rect 82082 390688 82138 390697
rect 81452 390646 82082 390674
rect 77096 390374 77248 390402
rect 77220 384985 77248 390374
rect 77404 390374 77832 390402
rect 78048 390374 78384 390402
rect 77300 387048 77352 387054
rect 77300 386990 77352 386996
rect 77206 384976 77262 384985
rect 77206 384911 77262 384920
rect 76564 376032 76616 376038
rect 76564 375974 76616 375980
rect 74552 373966 75224 373994
rect 73066 356688 73122 356697
rect 73066 356623 73122 356632
rect 72422 338192 72478 338201
rect 72422 338127 72478 338136
rect 73066 338192 73122 338201
rect 73066 338127 73068 338136
rect 72436 306374 72464 338127
rect 73120 338127 73122 338136
rect 73068 338098 73120 338104
rect 73066 326360 73122 326369
rect 73066 326295 73122 326304
rect 72436 306346 72648 306374
rect 72620 292574 72648 306346
rect 72528 292546 72648 292574
rect 72424 291236 72476 291242
rect 72424 291178 72476 291184
rect 70492 287700 70544 287706
rect 70492 287642 70544 287648
rect 70308 285796 70360 285802
rect 70308 285738 70360 285744
rect 70320 283506 70348 285738
rect 70104 283478 70348 283506
rect 69000 283342 69152 283370
rect 69754 283384 69810 283393
rect 70504 283370 70532 287642
rect 72054 287056 72110 287065
rect 72054 286991 72110 287000
rect 71318 283520 71374 283529
rect 71208 283492 71318 283506
rect 71194 283478 71318 283492
rect 70504 283356 70656 283370
rect 70504 283342 70670 283356
rect 69754 283319 69810 283328
rect 70642 283098 70670 283342
rect 71042 283112 71098 283121
rect 70642 283084 70992 283098
rect 70656 283082 70992 283084
rect 70656 283076 71004 283082
rect 70656 283070 70952 283076
rect 71194 283098 71222 283478
rect 72068 283506 72096 286991
rect 72436 284345 72464 291178
rect 72528 288522 72556 292546
rect 72516 288516 72568 288522
rect 72516 288458 72568 288464
rect 72422 284336 72478 284345
rect 72422 284271 72478 284280
rect 72436 283506 72464 284271
rect 71760 283478 72096 283506
rect 72312 283478 72464 283506
rect 72528 283506 72556 288458
rect 73080 287065 73108 326295
rect 73252 290488 73304 290494
rect 73252 290430 73304 290436
rect 73158 289912 73214 289921
rect 73158 289847 73214 289856
rect 73066 287056 73122 287065
rect 73066 286991 73122 287000
rect 73172 284209 73200 289847
rect 73158 284200 73214 284209
rect 73158 284135 73214 284144
rect 72528 283478 72864 283506
rect 71318 283455 71374 283464
rect 73172 283370 73200 284135
rect 73264 283490 73292 290430
rect 74552 290057 74580 373966
rect 77312 362914 77340 386990
rect 77404 381546 77432 390374
rect 78048 387054 78076 390374
rect 79106 390130 79134 390388
rect 79244 390374 79856 390402
rect 80072 390374 80592 390402
rect 80992 390374 81328 390402
rect 79106 390102 79180 390130
rect 79152 389065 79180 390102
rect 79138 389056 79194 389065
rect 79138 388991 79194 389000
rect 78036 387048 78088 387054
rect 78036 386990 78088 386996
rect 77392 381540 77444 381546
rect 77392 381482 77444 381488
rect 79244 373994 79272 390374
rect 79966 389056 80022 389065
rect 79966 388991 80022 389000
rect 78692 373966 79272 373994
rect 77300 362908 77352 362914
rect 77300 362850 77352 362856
rect 77390 320240 77446 320249
rect 77390 320175 77446 320184
rect 77300 305040 77352 305046
rect 75182 305008 75238 305017
rect 77300 304982 77352 304988
rect 75182 304943 75238 304952
rect 75196 292574 75224 304943
rect 76012 295996 76064 296002
rect 76012 295938 76064 295944
rect 74920 292546 75224 292574
rect 74538 290048 74594 290057
rect 74538 289983 74594 289992
rect 73620 285728 73672 285734
rect 73620 285670 73672 285676
rect 73632 283506 73660 285670
rect 74920 284345 74948 292546
rect 76024 291242 76052 295938
rect 76012 291236 76064 291242
rect 76012 291178 76064 291184
rect 77024 290488 77076 290494
rect 77024 290430 77076 290436
rect 75828 287020 75880 287026
rect 75828 286962 75880 286968
rect 74906 284336 74962 284345
rect 74906 284271 74962 284280
rect 74920 283506 74948 284271
rect 75840 283506 75868 286962
rect 75918 285832 75974 285841
rect 75918 285767 75974 285776
rect 76012 285796 76064 285802
rect 73252 283484 73304 283490
rect 73632 283478 73968 283506
rect 74520 283478 74948 283506
rect 75624 283478 75868 283506
rect 75932 283506 75960 285767
rect 76012 285738 76064 285744
rect 76024 284889 76052 285738
rect 76010 284880 76066 284889
rect 76010 284815 76066 284824
rect 77036 283506 77064 290430
rect 77312 283778 77340 304982
rect 75932 283478 76176 283506
rect 76728 283478 77064 283506
rect 77266 283750 77340 283778
rect 77266 283492 77294 283750
rect 77404 283506 77432 320175
rect 77944 299600 77996 299606
rect 77944 299542 77996 299548
rect 77956 287026 77984 299542
rect 78692 287774 78720 373966
rect 79980 368393 80008 388991
rect 80072 382974 80100 390374
rect 80992 389065 81020 390374
rect 80150 389056 80206 389065
rect 80150 388991 80206 389000
rect 80978 389056 81034 389065
rect 80978 388991 81034 389000
rect 80060 382968 80112 382974
rect 80060 382910 80112 382916
rect 79966 368384 80022 368393
rect 79966 368319 80022 368328
rect 79324 323604 79376 323610
rect 79324 323546 79376 323552
rect 79336 289241 79364 323546
rect 79966 294536 80022 294545
rect 79966 294471 80022 294480
rect 79322 289232 79378 289241
rect 79322 289167 79378 289176
rect 79690 289096 79746 289105
rect 79690 289031 79746 289040
rect 78680 287768 78732 287774
rect 78680 287710 78732 287716
rect 77944 287020 77996 287026
rect 77944 286962 77996 286968
rect 79232 287020 79284 287026
rect 79232 286962 79284 286968
rect 78588 285796 78640 285802
rect 78588 285738 78640 285744
rect 78600 283506 78628 285738
rect 79244 283506 79272 286962
rect 79704 283506 79732 289031
rect 79980 287026 80008 294471
rect 80164 291825 80192 388991
rect 81452 388906 81480 390646
rect 82082 390623 82138 390632
rect 83200 390646 83352 390674
rect 81268 388878 81480 388906
rect 82004 390374 82616 390402
rect 81268 388385 81296 388878
rect 81254 388376 81310 388385
rect 81254 388311 81310 388320
rect 81268 370530 81296 388311
rect 81346 382936 81402 382945
rect 81346 382871 81402 382880
rect 81256 370524 81308 370530
rect 81256 370466 81308 370472
rect 80150 291816 80206 291825
rect 80150 291751 80206 291760
rect 80886 291272 80942 291281
rect 80886 291207 80942 291216
rect 79968 287020 80020 287026
rect 79968 286962 80020 286968
rect 80152 285660 80204 285666
rect 80152 285602 80204 285608
rect 77404 283478 77832 283506
rect 78384 283478 78628 283506
rect 78936 283478 79272 283506
rect 79488 283478 79732 283506
rect 73252 283426 73304 283432
rect 74724 283416 74776 283422
rect 73172 283342 73416 283370
rect 80164 283370 80192 285602
rect 80900 283506 80928 291207
rect 81360 283506 81388 382871
rect 82004 373994 82032 390374
rect 83200 387569 83228 390646
rect 89258 390552 89314 390561
rect 89314 390524 89608 390538
rect 89314 390510 89622 390524
rect 93840 390510 93992 390538
rect 89258 390487 89314 390496
rect 83476 390374 84088 390402
rect 84304 390374 84824 390402
rect 85040 390374 85376 390402
rect 86112 390374 86632 390402
rect 83186 387560 83242 387569
rect 83186 387495 83242 387504
rect 83476 383654 83504 390374
rect 84200 387048 84252 387054
rect 84200 386990 84252 386996
rect 81452 373966 82032 373994
rect 82832 383626 83504 383654
rect 81452 371890 81480 373966
rect 81440 371884 81492 371890
rect 81440 371826 81492 371832
rect 82832 359514 82860 383626
rect 83464 383036 83516 383042
rect 83464 382978 83516 382984
rect 83476 369753 83504 382978
rect 83462 369744 83518 369753
rect 83462 369679 83518 369688
rect 82820 359508 82872 359514
rect 82820 359450 82872 359456
rect 84212 354006 84240 386990
rect 84304 377466 84332 390374
rect 85040 387054 85068 390374
rect 85028 387048 85080 387054
rect 85028 386990 85080 386996
rect 86604 383654 86632 390374
rect 86834 390130 86862 390388
rect 87064 390374 87584 390402
rect 87800 390374 88136 390402
rect 88872 390374 89208 390402
rect 86834 390102 86908 390130
rect 86776 389836 86828 389842
rect 86776 389778 86828 389784
rect 86788 384826 86816 389778
rect 86880 385014 86908 390102
rect 86868 385008 86920 385014
rect 86868 384950 86920 384956
rect 86788 384798 86908 384826
rect 86604 383626 86816 383654
rect 84292 377460 84344 377466
rect 84292 377402 84344 377408
rect 86788 365022 86816 383626
rect 86776 365016 86828 365022
rect 86776 364958 86828 364964
rect 86880 362234 86908 384798
rect 86868 362228 86920 362234
rect 86868 362170 86920 362176
rect 84200 354000 84252 354006
rect 84200 353942 84252 353948
rect 86866 320784 86922 320793
rect 86866 320719 86922 320728
rect 84842 318744 84898 318753
rect 84842 318679 84898 318688
rect 82726 317520 82782 317529
rect 82726 317455 82728 317464
rect 82780 317455 82782 317464
rect 82728 317426 82780 317432
rect 82726 316840 82782 316849
rect 82726 316775 82782 316784
rect 82740 292574 82768 316775
rect 82910 312488 82966 312497
rect 82910 312423 82966 312432
rect 82924 306374 82952 312423
rect 82924 306346 83412 306374
rect 82648 292546 82768 292574
rect 82648 290057 82676 292546
rect 83094 291952 83150 291961
rect 83094 291887 83150 291896
rect 82634 290048 82690 290057
rect 82634 289983 82690 289992
rect 81992 286476 82044 286482
rect 81992 286418 82044 286424
rect 82004 283506 82032 286418
rect 82648 283506 82676 289983
rect 83108 283506 83136 291887
rect 83186 290456 83242 290465
rect 83186 290391 83242 290400
rect 80592 283478 80928 283506
rect 81144 283478 81388 283506
rect 81696 283478 82032 283506
rect 82248 283478 82676 283506
rect 82800 283478 83136 283506
rect 74724 283358 74776 283364
rect 74736 283234 74764 283358
rect 80040 283342 80192 283370
rect 74736 283206 75072 283234
rect 71098 283084 71222 283098
rect 75366 283112 75422 283121
rect 71098 283070 71208 283084
rect 71042 283047 71098 283056
rect 75366 283047 75422 283056
rect 70952 283018 71004 283024
rect 75380 283014 75408 283047
rect 81268 283014 81296 283478
rect 83200 283370 83228 290391
rect 83384 285818 83412 306346
rect 83462 305008 83518 305017
rect 83462 304943 83518 304952
rect 83476 286482 83504 304943
rect 84200 293276 84252 293282
rect 84200 293218 84252 293224
rect 83464 286476 83516 286482
rect 83464 286418 83516 286424
rect 83384 285790 83504 285818
rect 83476 283506 83504 285790
rect 84212 283506 84240 293218
rect 84856 290494 84884 318679
rect 86222 316704 86278 316713
rect 86222 316639 86278 316648
rect 86236 305046 86264 316639
rect 86224 305040 86276 305046
rect 86224 304982 86276 304988
rect 86776 304360 86828 304366
rect 86776 304302 86828 304308
rect 86788 291281 86816 304302
rect 85854 291272 85910 291281
rect 85854 291207 85910 291216
rect 86774 291272 86830 291281
rect 86774 291207 86830 291216
rect 84844 290488 84896 290494
rect 84844 290430 84896 290436
rect 85868 283506 85896 291207
rect 86880 287473 86908 320719
rect 87064 300801 87092 390374
rect 87800 389842 87828 390374
rect 87788 389836 87840 389842
rect 87788 389778 87840 389784
rect 89180 387569 89208 390374
rect 89594 390130 89622 390510
rect 91926 390416 91982 390425
rect 89548 390102 89622 390130
rect 89732 390374 90344 390402
rect 89166 387560 89222 387569
rect 89166 387495 89222 387504
rect 88982 384296 89038 384305
rect 88982 384231 89038 384240
rect 88248 375352 88300 375358
rect 88248 375294 88300 375300
rect 88260 313342 88288 375294
rect 88996 366994 89024 384231
rect 89548 381585 89576 390102
rect 89628 385076 89680 385082
rect 89628 385018 89680 385024
rect 89534 381576 89590 381585
rect 89534 381511 89590 381520
rect 88984 366988 89036 366994
rect 88984 366930 89036 366936
rect 87604 313336 87656 313342
rect 87604 313278 87656 313284
rect 88248 313336 88300 313342
rect 88248 313278 88300 313284
rect 87050 300792 87106 300801
rect 87050 300727 87106 300736
rect 86406 287464 86462 287473
rect 86406 287399 86462 287408
rect 86866 287464 86922 287473
rect 86866 287399 86922 287408
rect 86420 283506 86448 287399
rect 86868 286340 86920 286346
rect 86868 286282 86920 286288
rect 86880 283506 86908 286282
rect 87510 285696 87566 285705
rect 87510 285631 87566 285640
rect 87524 283506 87552 285631
rect 87616 284209 87644 313278
rect 88982 308000 89038 308009
rect 88982 307935 89038 307944
rect 88616 290488 88668 290494
rect 88616 290430 88668 290436
rect 88064 287156 88116 287162
rect 88064 287098 88116 287104
rect 87602 284200 87658 284209
rect 87602 284135 87658 284144
rect 88076 283506 88104 287098
rect 88628 283529 88656 290430
rect 88996 286346 89024 307935
rect 89534 302832 89590 302841
rect 89534 302767 89590 302776
rect 88984 286340 89036 286346
rect 88984 286282 89036 286288
rect 89166 284472 89222 284481
rect 89166 284407 89222 284416
rect 88614 283520 88670 283529
rect 83476 283478 83904 283506
rect 84212 283478 84456 283506
rect 85560 283478 85896 283506
rect 86112 283478 86448 283506
rect 86664 283478 86908 283506
rect 87216 283478 87552 283506
rect 87768 283478 88104 283506
rect 88320 283478 88614 283506
rect 89180 283506 89208 284407
rect 89548 283506 89576 302767
rect 89640 284481 89668 385018
rect 89732 300801 89760 390374
rect 91066 390130 91094 390388
rect 91204 390374 91632 390402
rect 91066 390102 91140 390130
rect 91112 387025 91140 390102
rect 91098 387016 91154 387025
rect 91098 386951 91154 386960
rect 91006 383752 91062 383761
rect 91006 383687 91062 383696
rect 90914 319424 90970 319433
rect 90914 319359 90970 319368
rect 89718 300792 89774 300801
rect 89718 300727 89774 300736
rect 90928 289921 90956 319359
rect 90914 289912 90970 289921
rect 90914 289847 90970 289856
rect 90272 288516 90324 288522
rect 90272 288458 90324 288464
rect 89626 284472 89682 284481
rect 89626 284407 89682 284416
rect 90284 283506 90312 288458
rect 90824 285796 90876 285802
rect 90824 285738 90876 285744
rect 90836 283506 90864 285738
rect 90928 285705 90956 289847
rect 91020 289134 91048 383687
rect 91204 373994 91232 390374
rect 91982 390374 92368 390402
rect 92492 390374 93104 390402
rect 91926 390351 91982 390360
rect 91940 375358 91968 390351
rect 92492 379438 92520 390374
rect 93964 387802 93992 390510
rect 94392 390374 94728 390402
rect 94700 389230 94728 390374
rect 94792 390374 95128 390402
rect 94688 389224 94740 389230
rect 94688 389166 94740 389172
rect 94318 388240 94374 388249
rect 94318 388175 94374 388184
rect 93952 387796 94004 387802
rect 93952 387738 94004 387744
rect 94332 385082 94360 388175
rect 94792 387977 94820 390374
rect 94778 387968 94834 387977
rect 94778 387903 94834 387912
rect 94504 387796 94556 387802
rect 94504 387738 94556 387744
rect 94320 385076 94372 385082
rect 94320 385018 94372 385024
rect 92480 379432 92532 379438
rect 92480 379374 92532 379380
rect 91928 375352 91980 375358
rect 91928 375294 91980 375300
rect 91112 373966 91232 373994
rect 91112 292641 91140 373966
rect 94516 373318 94544 387738
rect 94504 373312 94556 373318
rect 94504 373254 94556 373260
rect 92480 339516 92532 339522
rect 92480 339458 92532 339464
rect 91192 301504 91244 301510
rect 91192 301446 91244 301452
rect 91098 292632 91154 292641
rect 91098 292567 91154 292576
rect 91008 289128 91060 289134
rect 91008 289070 91060 289076
rect 91020 288522 91048 289070
rect 91008 288516 91060 288522
rect 91008 288458 91060 288464
rect 90914 285696 90970 285705
rect 90914 285631 90970 285640
rect 91204 283506 91232 301446
rect 91926 285832 91982 285841
rect 91926 285767 91982 285776
rect 91940 283506 91968 285767
rect 92388 284368 92440 284374
rect 92388 284310 92440 284316
rect 92400 283506 92428 284310
rect 88872 283478 89208 283506
rect 89424 283478 89576 283506
rect 89976 283478 90312 283506
rect 90528 283478 90864 283506
rect 91080 283478 91232 283506
rect 91632 283478 91968 283506
rect 92184 283478 92428 283506
rect 88614 283455 88670 283464
rect 88628 283395 88656 283455
rect 83462 283384 83518 283393
rect 83200 283342 83462 283370
rect 83462 283319 83518 283328
rect 89548 283014 89576 283478
rect 92492 283422 92520 339458
rect 95146 320240 95202 320249
rect 95146 320175 95202 320184
rect 95054 318064 95110 318073
rect 95054 317999 95110 318008
rect 95068 300218 95096 317999
rect 93952 300212 94004 300218
rect 93952 300154 94004 300160
rect 95056 300212 95108 300218
rect 95056 300154 95108 300160
rect 93766 294536 93822 294545
rect 93766 294471 93822 294480
rect 93124 293344 93176 293350
rect 93124 293286 93176 293292
rect 93136 283506 93164 293286
rect 93780 287162 93808 294471
rect 93768 287156 93820 287162
rect 93768 287098 93820 287104
rect 93858 285696 93914 285705
rect 93858 285631 93914 285640
rect 93872 283778 93900 285631
rect 92736 283478 93164 283506
rect 93826 283750 93900 283778
rect 93826 283492 93854 283750
rect 93964 283506 93992 300154
rect 95068 299538 95096 300154
rect 95056 299532 95108 299538
rect 95056 299474 95108 299480
rect 95160 283506 95188 320175
rect 95252 305017 95280 390782
rect 96724 390697 96752 390782
rect 95330 390688 95386 390697
rect 95330 390623 95386 390632
rect 96710 390688 96766 390697
rect 96710 390623 96766 390632
rect 95238 305008 95294 305017
rect 95238 304943 95294 304952
rect 95344 304366 95372 390623
rect 96712 390516 96764 390522
rect 96712 390458 96764 390464
rect 96724 373994 96752 390458
rect 96908 389065 96936 390782
rect 104254 390688 104310 390697
rect 104144 390646 104254 390674
rect 105082 390688 105138 390697
rect 104310 390646 104572 390674
rect 104880 390646 105082 390674
rect 104254 390623 104310 390632
rect 100942 390552 100998 390561
rect 97552 390522 97888 390538
rect 97540 390516 97888 390522
rect 97592 390510 97888 390516
rect 100832 390510 100942 390538
rect 100942 390487 100998 390496
rect 97540 390458 97592 390464
rect 96986 390416 97042 390425
rect 97042 390374 97764 390402
rect 96986 390351 97042 390360
rect 96894 389056 96950 389065
rect 96894 388991 96950 389000
rect 97630 389056 97686 389065
rect 97630 388991 97686 389000
rect 97644 377466 97672 388991
rect 97736 382226 97764 390374
rect 98012 390374 98624 390402
rect 99360 390374 99512 390402
rect 100096 390374 100432 390402
rect 101384 390374 101720 390402
rect 102120 390374 102456 390402
rect 102856 390374 103192 390402
rect 103592 390374 103928 390402
rect 98012 383654 98040 390374
rect 99484 389337 99512 390374
rect 99470 389328 99526 389337
rect 99470 389263 99526 389272
rect 99484 387802 99512 389263
rect 99562 388512 99618 388521
rect 99562 388447 99618 388456
rect 99472 387796 99524 387802
rect 99472 387738 99524 387744
rect 98000 383648 98052 383654
rect 98000 383590 98052 383596
rect 97724 382220 97776 382226
rect 97724 382162 97776 382168
rect 97264 377460 97316 377466
rect 97264 377402 97316 377408
rect 97632 377460 97684 377466
rect 97632 377402 97684 377408
rect 96632 373966 96752 373994
rect 96526 305688 96582 305697
rect 96526 305623 96582 305632
rect 95332 304360 95384 304366
rect 95332 304302 95384 304308
rect 96540 292574 96568 305623
rect 96632 298761 96660 373966
rect 97276 360126 97304 377402
rect 97264 360120 97316 360126
rect 97264 360062 97316 360068
rect 97906 323640 97962 323649
rect 97906 323575 97962 323584
rect 96618 298752 96674 298761
rect 96618 298687 96674 298696
rect 96620 294636 96672 294642
rect 96620 294578 96672 294584
rect 96448 292546 96568 292574
rect 95790 287192 95846 287201
rect 95790 287127 95846 287136
rect 95804 283506 95832 287127
rect 96448 284442 96476 292546
rect 96436 284436 96488 284442
rect 96436 284378 96488 284384
rect 96448 283506 96476 284378
rect 96632 283778 96660 294578
rect 97920 286618 97948 323575
rect 98000 320204 98052 320210
rect 98000 320146 98052 320152
rect 98012 306374 98040 320146
rect 99286 319424 99342 319433
rect 99286 319359 99342 319368
rect 98012 306346 98592 306374
rect 98460 291236 98512 291242
rect 98460 291178 98512 291184
rect 97448 286612 97500 286618
rect 97448 286554 97500 286560
rect 97908 286612 97960 286618
rect 97908 286554 97960 286560
rect 97460 284345 97488 286554
rect 97446 284336 97502 284345
rect 97446 284271 97502 284280
rect 93964 283478 94392 283506
rect 94944 283478 95188 283506
rect 95496 283478 95832 283506
rect 96048 283478 96476 283506
rect 96586 283750 96660 283778
rect 96586 283492 96614 283750
rect 97460 283506 97488 284271
rect 98472 283506 98500 291178
rect 98564 283778 98592 306346
rect 99300 292534 99328 319359
rect 99288 292528 99340 292534
rect 99288 292470 99340 292476
rect 99300 291242 99328 292470
rect 99288 291236 99340 291242
rect 99288 291178 99340 291184
rect 99576 290494 99604 388447
rect 100404 384946 100432 390374
rect 101692 387734 101720 390374
rect 102046 390280 102102 390289
rect 102046 390215 102102 390224
rect 102060 389201 102088 390215
rect 102428 389473 102456 390374
rect 102414 389464 102470 389473
rect 102414 389399 102470 389408
rect 102046 389192 102102 389201
rect 102046 389127 102102 389136
rect 101680 387728 101732 387734
rect 101680 387670 101732 387676
rect 100392 384940 100444 384946
rect 100392 384882 100444 384888
rect 101494 384296 101550 384305
rect 101494 384231 101550 384240
rect 101404 369164 101456 369170
rect 101404 369106 101456 369112
rect 100758 320240 100814 320249
rect 100758 320175 100814 320184
rect 100772 320074 100800 320175
rect 100760 320068 100812 320074
rect 100760 320010 100812 320016
rect 100022 291952 100078 291961
rect 100022 291887 100078 291896
rect 99564 290488 99616 290494
rect 99564 290430 99616 290436
rect 99012 284368 99064 284374
rect 99012 284310 99064 284316
rect 98564 283750 98638 283778
rect 97152 283478 97488 283506
rect 98256 283478 98500 283506
rect 92480 283416 92532 283422
rect 92480 283358 92532 283364
rect 92940 283416 92992 283422
rect 92992 283364 93288 283370
rect 92940 283358 93288 283364
rect 92952 283342 93288 283358
rect 97906 283112 97962 283121
rect 97704 283070 97906 283098
rect 97906 283047 97962 283056
rect 75368 283008 75420 283014
rect 75368 282950 75420 282956
rect 81256 283008 81308 283014
rect 89536 283008 89588 283014
rect 85302 282976 85358 282985
rect 81256 282950 81308 282956
rect 85008 282934 85302 282962
rect 89536 282950 89588 282956
rect 85302 282911 85358 282920
rect 98000 282872 98052 282878
rect 98610 282826 98638 283750
rect 98828 283076 98880 283082
rect 98828 283018 98880 283024
rect 98000 282814 98052 282820
rect 98012 281586 98040 282814
rect 98380 282812 98638 282826
rect 98380 282798 98624 282812
rect 98000 281580 98052 281586
rect 98000 281522 98052 281528
rect 98380 273254 98408 282798
rect 98840 279478 98868 283018
rect 98918 282840 98974 282849
rect 98918 282775 98974 282784
rect 98932 281654 98960 282775
rect 98920 281648 98972 281654
rect 98920 281590 98972 281596
rect 98828 279472 98880 279478
rect 98828 279414 98880 279420
rect 99024 276010 99052 284310
rect 99104 283280 99156 283286
rect 99104 283222 99156 283228
rect 99116 278730 99144 283222
rect 99104 278724 99156 278730
rect 99104 278666 99156 278672
rect 99012 276004 99064 276010
rect 99012 275946 99064 275952
rect 98196 273226 98408 273254
rect 98090 258496 98146 258505
rect 98090 258431 98146 258440
rect 68664 248386 68968 248414
rect 68652 242956 68704 242962
rect 68652 242898 68704 242904
rect 68664 242298 68692 242898
rect 68664 242270 68816 242298
rect 68940 241398 68968 248386
rect 98000 243568 98052 243574
rect 98000 243510 98052 243516
rect 75368 241800 75420 241806
rect 69478 241768 69534 241777
rect 72698 241768 72754 241777
rect 69534 241726 69736 241754
rect 72496 241726 72698 241754
rect 69478 241703 69534 241712
rect 72698 241703 72754 241712
rect 73250 241768 73306 241777
rect 73250 241703 73306 241712
rect 73802 241768 73858 241777
rect 73858 241726 74152 241754
rect 95976 241800 96028 241806
rect 83738 241768 83794 241777
rect 75368 241742 75420 241748
rect 73802 241703 73858 241712
rect 69184 241590 69520 241618
rect 70288 241590 70348 241618
rect 68928 241392 68980 241398
rect 68928 241334 68980 241340
rect 69492 240106 69520 241590
rect 70320 241505 70348 241590
rect 69662 241496 69718 241505
rect 69662 241431 69718 241440
rect 70306 241496 70362 241505
rect 70306 241431 70362 241440
rect 69480 240100 69532 240106
rect 69480 240042 69532 240048
rect 69202 240000 69258 240009
rect 69202 239935 69258 239944
rect 69216 238814 69244 239935
rect 69204 238808 69256 238814
rect 69204 238750 69256 238756
rect 67824 169788 67876 169794
rect 67824 169730 67876 169736
rect 68560 169788 68612 169794
rect 68560 169730 68612 169736
rect 67732 149728 67784 149734
rect 67732 149670 67784 149676
rect 67744 112441 67772 149670
rect 67836 132841 67864 169730
rect 69294 139496 69350 139505
rect 69294 139431 69350 139440
rect 68652 134836 68704 134842
rect 68652 134778 68704 134784
rect 67822 132832 67878 132841
rect 67822 132767 67878 132776
rect 67730 112432 67786 112441
rect 67730 112367 67786 112376
rect 67730 110800 67786 110809
rect 67730 110735 67786 110744
rect 67560 103486 67680 103514
rect 67454 98016 67510 98025
rect 67454 97951 67510 97960
rect 67362 97200 67418 97209
rect 67362 97135 67418 97144
rect 66902 95840 66958 95849
rect 66902 95775 66958 95784
rect 66916 95266 66944 95775
rect 66904 95260 66956 95266
rect 66904 95202 66956 95208
rect 66812 95192 66864 95198
rect 66812 95134 66864 95140
rect 66824 95033 66852 95134
rect 66810 95024 66866 95033
rect 66810 94959 66866 94968
rect 67270 94208 67326 94217
rect 67270 94143 67326 94152
rect 66168 66156 66220 66162
rect 66168 66098 66220 66104
rect 67284 63481 67312 94143
rect 67376 86737 67404 97135
rect 67468 89010 67496 97951
rect 67560 92886 67588 103486
rect 67548 92880 67600 92886
rect 67548 92822 67600 92828
rect 67546 92576 67602 92585
rect 67546 92511 67548 92520
rect 67600 92511 67602 92520
rect 67548 92482 67600 92488
rect 67456 89004 67508 89010
rect 67456 88946 67508 88952
rect 67362 86728 67418 86737
rect 67362 86663 67418 86672
rect 67744 80034 67772 110735
rect 67824 103488 67876 103494
rect 67824 103430 67876 103436
rect 67836 103193 67864 103430
rect 67822 103184 67878 103193
rect 67822 103119 67878 103128
rect 67732 80028 67784 80034
rect 67732 79970 67784 79976
rect 67836 71738 67864 103119
rect 68664 93854 68692 134778
rect 69308 134722 69336 139431
rect 69572 135040 69624 135046
rect 69570 135008 69572 135017
rect 69624 135008 69626 135017
rect 69570 134943 69626 134952
rect 69676 134842 69704 241431
rect 70826 241369 70854 241604
rect 71332 241590 71392 241618
rect 71944 241590 72280 241618
rect 71332 241369 71360 241590
rect 70812 241360 70868 241369
rect 70812 241295 70868 241304
rect 71318 241360 71374 241369
rect 71318 241295 71374 241304
rect 71332 240145 71360 241295
rect 72252 240145 72280 241590
rect 72620 241590 73048 241618
rect 71318 240136 71374 240145
rect 71318 240071 71374 240080
rect 72238 240136 72294 240145
rect 72238 240071 72294 240080
rect 72620 238754 72648 241590
rect 71792 238726 72648 238754
rect 71686 237552 71742 237561
rect 71686 237487 71742 237496
rect 71044 178084 71096 178090
rect 71044 178026 71096 178032
rect 70584 155304 70636 155310
rect 70584 155246 70636 155252
rect 70030 138272 70086 138281
rect 70030 138207 70086 138216
rect 69846 137320 69902 137329
rect 69846 137255 69902 137264
rect 69664 134836 69716 134842
rect 69664 134778 69716 134784
rect 69860 134722 69888 137255
rect 70044 135028 70072 138207
rect 70596 135028 70624 155246
rect 71056 138417 71084 178026
rect 71700 139369 71728 237487
rect 71792 233238 71820 238726
rect 71780 233232 71832 233238
rect 71780 233174 71832 233180
rect 73068 233232 73120 233238
rect 73068 233174 73120 233180
rect 72976 159384 73028 159390
rect 72976 159326 73028 159332
rect 72882 156496 72938 156505
rect 72882 156431 72938 156440
rect 72896 155990 72924 156431
rect 71780 155984 71832 155990
rect 71780 155926 71832 155932
rect 72884 155984 72936 155990
rect 72884 155926 72936 155932
rect 71686 139360 71742 139369
rect 71686 139295 71742 139304
rect 71228 138712 71280 138718
rect 71228 138654 71280 138660
rect 71134 138544 71190 138553
rect 71134 138479 71190 138488
rect 71042 138408 71098 138417
rect 71042 138343 71098 138352
rect 70044 135000 70118 135028
rect 70596 135000 70670 135028
rect 69000 134694 69336 134722
rect 69552 134694 69888 134722
rect 70090 134708 70118 135000
rect 70642 134708 70670 135000
rect 71148 134722 71176 138479
rect 71024 134694 71176 134722
rect 71240 134722 71268 138654
rect 71700 138553 71728 139295
rect 71686 138544 71742 138553
rect 71686 138479 71742 138488
rect 71792 134722 71820 155926
rect 72332 141432 72384 141438
rect 72332 141374 72384 141380
rect 72344 134722 72372 141374
rect 72988 137970 73016 159326
rect 72976 137964 73028 137970
rect 72976 137906 73028 137912
rect 72988 136746 73016 137906
rect 72976 136740 73028 136746
rect 72976 136682 73028 136688
rect 73080 134745 73108 233174
rect 73264 210458 73292 241703
rect 73600 241590 73936 241618
rect 73908 240038 73936 241590
rect 74690 241466 74718 241604
rect 74920 241590 75256 241618
rect 74678 241460 74730 241466
rect 74678 241402 74730 241408
rect 74920 240145 74948 241590
rect 74906 240136 74962 240145
rect 74906 240071 74962 240080
rect 73896 240032 73948 240038
rect 73896 239974 73948 239980
rect 74814 239864 74870 239873
rect 74814 239799 74870 239808
rect 73436 236768 73488 236774
rect 73436 236710 73488 236716
rect 73252 210452 73304 210458
rect 73252 210394 73304 210400
rect 73160 136740 73212 136746
rect 73160 136682 73212 136688
rect 73172 135028 73200 136682
rect 73172 135000 73246 135028
rect 73066 134736 73122 134745
rect 71240 134694 71576 134722
rect 71792 134694 72128 134722
rect 72344 134694 72680 134722
rect 73218 134708 73246 135000
rect 73448 134722 73476 236710
rect 74828 236706 74856 239799
rect 74632 236700 74684 236706
rect 74632 236642 74684 236648
rect 74816 236700 74868 236706
rect 74816 236642 74868 236648
rect 74538 164384 74594 164393
rect 74538 164319 74594 164328
rect 73804 144220 73856 144226
rect 73804 144162 73856 144168
rect 73816 135046 73844 144162
rect 74448 136740 74500 136746
rect 74448 136682 74500 136688
rect 73804 135040 73856 135046
rect 73804 134982 73856 134988
rect 74460 134722 74488 136682
rect 73448 134694 73600 134722
rect 74152 134694 74488 134722
rect 74552 134722 74580 164319
rect 74644 155310 74672 236642
rect 75380 177410 75408 241742
rect 83536 241726 83738 241754
rect 86590 241768 86646 241777
rect 86296 241726 86590 241754
rect 83738 241703 83794 241712
rect 86590 241703 86646 241712
rect 87142 241768 87198 241777
rect 90362 241768 90418 241777
rect 87198 241726 87552 241754
rect 90160 241726 90362 241754
rect 87142 241703 87198 241712
rect 82636 241664 82688 241670
rect 75472 241590 75808 241618
rect 76024 241590 76360 241618
rect 76576 241590 76912 241618
rect 77464 241590 77524 241618
rect 75472 239873 75500 241590
rect 75920 240168 75972 240174
rect 75920 240110 75972 240116
rect 75458 239864 75514 239873
rect 75458 239799 75514 239808
rect 75932 215393 75960 240110
rect 76024 233170 76052 241590
rect 76576 240174 76604 241590
rect 77496 241398 77524 241590
rect 77588 241590 78016 241618
rect 78140 241590 78568 241618
rect 78692 241590 79120 241618
rect 79336 241590 79672 241618
rect 80164 241590 80224 241618
rect 80348 241590 80776 241618
rect 80992 241590 81328 241618
rect 81880 241590 82216 241618
rect 82432 241612 82636 241618
rect 85946 241632 86002 241641
rect 82432 241606 82688 241612
rect 82432 241604 82676 241606
rect 77484 241392 77536 241398
rect 77484 241334 77536 241340
rect 76564 240168 76616 240174
rect 76564 240110 76616 240116
rect 77496 239970 77524 241334
rect 77484 239964 77536 239970
rect 77484 239906 77536 239912
rect 77588 236745 77616 241590
rect 78140 240122 78168 241590
rect 77680 240094 78168 240122
rect 77680 238746 77708 240094
rect 77944 239964 77996 239970
rect 77944 239906 77996 239912
rect 77668 238740 77720 238746
rect 77668 238682 77720 238688
rect 77680 237454 77708 238682
rect 77668 237448 77720 237454
rect 77668 237390 77720 237396
rect 77574 236736 77630 236745
rect 77574 236671 77630 236680
rect 76012 233164 76064 233170
rect 76012 233106 76064 233112
rect 76564 233164 76616 233170
rect 76564 233106 76616 233112
rect 75918 215384 75974 215393
rect 75918 215319 75974 215328
rect 75368 177404 75420 177410
rect 75368 177346 75420 177352
rect 75920 171828 75972 171834
rect 75920 171770 75972 171776
rect 75182 157448 75238 157457
rect 75182 157383 75238 157392
rect 74632 155304 74684 155310
rect 74632 155246 74684 155252
rect 75196 136746 75224 157383
rect 75932 151814 75960 171770
rect 75932 151786 76328 151814
rect 76196 147688 76248 147694
rect 76196 147630 76248 147636
rect 76208 142769 76236 147630
rect 76194 142760 76250 142769
rect 76194 142695 76250 142704
rect 76196 141500 76248 141506
rect 76196 141442 76248 141448
rect 75828 141432 75880 141438
rect 75828 141374 75880 141380
rect 75550 137728 75606 137737
rect 75550 137663 75606 137672
rect 75184 136740 75236 136746
rect 75184 136682 75236 136688
rect 75564 134722 75592 137663
rect 75840 136785 75868 141374
rect 75826 136776 75882 136785
rect 75826 136711 75882 136720
rect 75840 135028 75868 136711
rect 76208 135028 76236 141442
rect 74552 134694 74704 134722
rect 75256 134694 75592 134722
rect 75794 135000 75868 135028
rect 76162 135000 76236 135028
rect 75794 134708 75822 135000
rect 76162 134708 76190 135000
rect 76300 134722 76328 151786
rect 76576 141574 76604 233106
rect 77484 231124 77536 231130
rect 77484 231066 77536 231072
rect 77496 230518 77524 231066
rect 77484 230512 77536 230518
rect 77484 230454 77536 230460
rect 77300 217320 77352 217326
rect 77300 217262 77352 217268
rect 76654 216064 76710 216073
rect 76654 215999 76710 216008
rect 76668 215393 76696 215999
rect 76654 215384 76710 215393
rect 76654 215319 76710 215328
rect 76564 141568 76616 141574
rect 76564 141510 76616 141516
rect 76668 140078 76696 215319
rect 76656 140072 76708 140078
rect 76656 140014 76708 140020
rect 77312 135028 77340 217262
rect 77392 163600 77444 163606
rect 77392 163542 77444 163548
rect 77404 138106 77432 163542
rect 77496 149734 77524 230454
rect 77956 218822 77984 239906
rect 78036 237448 78088 237454
rect 78036 237390 78088 237396
rect 77944 218816 77996 218822
rect 77944 218758 77996 218764
rect 78048 217297 78076 237390
rect 78034 217288 78090 217297
rect 78034 217223 78090 217232
rect 78692 213217 78720 241590
rect 79336 238754 79364 241590
rect 80060 240168 80112 240174
rect 80060 240110 80112 240116
rect 78784 238726 79364 238754
rect 78784 238649 78812 238726
rect 78770 238640 78826 238649
rect 78770 238575 78826 238584
rect 79968 237448 80020 237454
rect 79968 237390 80020 237396
rect 78678 213208 78734 213217
rect 78678 213143 78734 213152
rect 79980 206310 80008 237390
rect 80072 228410 80100 240110
rect 80164 237454 80192 241590
rect 80152 237448 80204 237454
rect 80152 237390 80204 237396
rect 80348 235929 80376 241590
rect 80992 240174 81020 241590
rect 81440 241528 81492 241534
rect 81440 241470 81492 241476
rect 80980 240168 81032 240174
rect 80980 240110 81032 240116
rect 80334 235920 80390 235929
rect 80334 235855 80390 235864
rect 80060 228404 80112 228410
rect 80060 228346 80112 228352
rect 79968 206304 80020 206310
rect 79968 206246 80020 206252
rect 80796 177336 80848 177342
rect 80796 177278 80848 177284
rect 80704 173188 80756 173194
rect 80704 173130 80756 173136
rect 77484 149728 77536 149734
rect 77484 149670 77536 149676
rect 77576 149184 77628 149190
rect 77576 149126 77628 149132
rect 77392 138100 77444 138106
rect 77392 138042 77444 138048
rect 77266 135000 77340 135028
rect 76300 134694 76728 134722
rect 77266 134708 77294 135000
rect 77588 134722 77616 149126
rect 80058 142896 80114 142905
rect 80058 142831 80114 142840
rect 78678 142760 78734 142769
rect 78678 142695 78734 142704
rect 77944 138100 77996 138106
rect 77944 138042 77996 138048
rect 77956 134722 77984 138042
rect 78692 135028 78720 142695
rect 80072 142154 80100 142831
rect 79704 142126 80100 142154
rect 78692 135000 78766 135028
rect 77588 134694 77832 134722
rect 77956 134694 78200 134722
rect 78738 134708 78766 135000
rect 79704 134722 79732 142126
rect 80610 140856 80666 140865
rect 80610 140791 80666 140800
rect 79874 138000 79930 138009
rect 79874 137935 79930 137944
rect 79888 134858 79916 137935
rect 79304 134694 79732 134722
rect 79842 134830 79916 134858
rect 79842 134708 79870 134830
rect 80624 134722 80652 140791
rect 80716 137329 80744 173130
rect 80808 149190 80836 177278
rect 80796 149184 80848 149190
rect 80796 149126 80848 149132
rect 81346 149152 81402 149161
rect 81346 149087 81402 149096
rect 81360 141409 81388 149087
rect 81346 141400 81402 141409
rect 81346 141335 81402 141344
rect 81360 140865 81388 141335
rect 81346 140856 81402 140865
rect 81346 140791 81402 140800
rect 81452 138825 81480 241470
rect 82188 238921 82216 241590
rect 82418 241590 82676 241604
rect 82832 241590 82984 241618
rect 84088 241590 84148 241618
rect 82418 241534 82446 241590
rect 82406 241528 82458 241534
rect 82406 241470 82458 241476
rect 82174 238912 82230 238921
rect 82174 238847 82230 238856
rect 82832 238678 82860 241590
rect 84120 241233 84148 241590
rect 84212 241590 84640 241618
rect 84764 241590 85192 241618
rect 85744 241590 85946 241618
rect 84106 241224 84162 241233
rect 84106 241159 84162 241168
rect 84106 238776 84162 238785
rect 84106 238711 84162 238720
rect 82820 238672 82872 238678
rect 82820 238614 82872 238620
rect 81532 169040 81584 169046
rect 81532 168982 81584 168988
rect 81438 138816 81494 138825
rect 81438 138751 81494 138760
rect 81438 138680 81494 138689
rect 81438 138615 81494 138624
rect 81452 138038 81480 138615
rect 81440 138032 81492 138038
rect 81440 137974 81492 137980
rect 80702 137320 80758 137329
rect 80702 137255 80758 137264
rect 81346 136912 81402 136921
rect 81346 136847 81402 136856
rect 81072 136740 81124 136746
rect 81072 136682 81124 136688
rect 81084 134722 81112 136682
rect 81360 134858 81388 136847
rect 80408 134694 80652 134722
rect 80776 134694 81112 134722
rect 81314 134830 81388 134858
rect 81314 134708 81342 134830
rect 81544 134722 81572 168982
rect 82912 167680 82964 167686
rect 82912 167622 82964 167628
rect 81990 144120 82046 144129
rect 81990 144055 82046 144064
rect 82004 134722 82032 144055
rect 82924 138106 82952 167622
rect 84120 162178 84148 238711
rect 84212 237386 84240 241590
rect 84764 238754 84792 241590
rect 85946 241567 86002 241576
rect 86604 241590 86848 241618
rect 86604 241505 86632 241590
rect 86590 241496 86646 241505
rect 86590 241431 86646 241440
rect 86788 239873 86816 241590
rect 86866 241496 86922 241505
rect 86866 241431 86922 241440
rect 86774 239864 86830 239873
rect 86774 239799 86830 239808
rect 84842 238912 84898 238921
rect 84842 238847 84898 238856
rect 84304 238746 84792 238754
rect 84292 238740 84792 238746
rect 84344 238726 84792 238740
rect 84292 238682 84344 238688
rect 84200 237380 84252 237386
rect 84200 237322 84252 237328
rect 84856 192574 84884 238847
rect 84936 236700 84988 236706
rect 84936 236642 84988 236648
rect 84948 195294 84976 236642
rect 84936 195288 84988 195294
rect 84936 195230 84988 195236
rect 84844 192568 84896 192574
rect 84844 192510 84896 192516
rect 86880 184278 86908 241431
rect 87524 240009 87552 241726
rect 90362 241703 90418 241712
rect 91558 241768 91614 241777
rect 93766 241768 93822 241777
rect 91614 241726 92244 241754
rect 91558 241703 91614 241712
rect 87616 241590 87952 241618
rect 88352 241590 88504 241618
rect 88720 241590 89056 241618
rect 89608 241590 89668 241618
rect 87510 240000 87566 240009
rect 87510 239935 87566 239944
rect 87616 238754 87644 241590
rect 88062 241496 88118 241505
rect 88062 241431 88118 241440
rect 88076 241233 88104 241431
rect 88062 241224 88118 241233
rect 88062 241159 88118 241168
rect 88246 240136 88302 240145
rect 88246 240071 88302 240080
rect 88154 240000 88210 240009
rect 88154 239935 88210 239944
rect 86972 238726 87644 238754
rect 86972 207738 87000 238726
rect 87604 218816 87656 218822
rect 87604 218758 87656 218764
rect 86960 207732 87012 207738
rect 86960 207674 87012 207680
rect 87616 187066 87644 218758
rect 88168 209098 88196 239935
rect 88260 217326 88288 240071
rect 88352 223582 88380 241590
rect 88720 240145 88748 241590
rect 89640 241233 89668 241590
rect 90376 241590 90712 241618
rect 91204 241590 91264 241618
rect 89626 241224 89682 241233
rect 89626 241159 89682 241168
rect 88706 240136 88762 240145
rect 88706 240071 88762 240080
rect 88982 239864 89038 239873
rect 88982 239799 89038 239808
rect 88340 223576 88392 223582
rect 88340 223518 88392 223524
rect 88248 217320 88300 217326
rect 88248 217262 88300 217268
rect 88248 210452 88300 210458
rect 88248 210394 88300 210400
rect 88156 209092 88208 209098
rect 88156 209034 88208 209040
rect 87604 187060 87656 187066
rect 87604 187002 87656 187008
rect 86868 184272 86920 184278
rect 86868 184214 86920 184220
rect 85580 174548 85632 174554
rect 85580 174490 85632 174496
rect 84842 174040 84898 174049
rect 84842 173975 84898 173984
rect 84200 166320 84252 166326
rect 84200 166262 84252 166268
rect 84108 162172 84160 162178
rect 84108 162114 84160 162120
rect 83462 156088 83518 156097
rect 83462 156023 83518 156032
rect 83002 149288 83058 149297
rect 83002 149223 83058 149232
rect 82912 138100 82964 138106
rect 82912 138042 82964 138048
rect 82910 136776 82966 136785
rect 82910 136711 82966 136720
rect 82924 134722 82952 136711
rect 81544 134694 81880 134722
rect 82004 134694 82432 134722
rect 82800 134694 82952 134722
rect 83016 134722 83044 149223
rect 83476 136746 83504 156023
rect 83554 152552 83610 152561
rect 83554 152487 83610 152496
rect 83568 151814 83596 152487
rect 83568 151786 83688 151814
rect 83556 138100 83608 138106
rect 83556 138042 83608 138048
rect 83464 136740 83516 136746
rect 83464 136682 83516 136688
rect 83568 134722 83596 138042
rect 83660 137737 83688 151786
rect 83646 137728 83702 137737
rect 83646 137663 83702 137672
rect 84212 134722 84240 166262
rect 84856 138009 84884 173975
rect 85592 151814 85620 174490
rect 86958 165744 87014 165753
rect 86958 165679 87014 165688
rect 86222 154592 86278 154601
rect 86222 154527 86278 154536
rect 85592 151786 86080 151814
rect 85948 140072 86000 140078
rect 85948 140014 86000 140020
rect 84842 138000 84898 138009
rect 84842 137935 84898 137944
rect 85486 136776 85542 136785
rect 85212 136740 85264 136746
rect 85486 136711 85542 136720
rect 85212 136682 85264 136688
rect 85224 134722 85252 136682
rect 85500 134722 85528 136711
rect 85960 134994 85988 140014
rect 83016 134694 83352 134722
rect 83568 134694 83904 134722
rect 84212 134694 84456 134722
rect 85008 134694 85252 134722
rect 85376 134694 85528 134722
rect 85914 134966 85988 134994
rect 85914 134708 85942 134966
rect 86052 134722 86080 151786
rect 86236 136921 86264 154527
rect 86316 149184 86368 149190
rect 86316 149126 86368 149132
rect 86222 136912 86278 136921
rect 86222 136847 86278 136856
rect 86328 136746 86356 149126
rect 86316 136740 86368 136746
rect 86316 136682 86368 136688
rect 86972 134994 87000 165679
rect 87142 160168 87198 160177
rect 88260 160138 88288 210394
rect 88996 182850 89024 239799
rect 90376 238754 90404 241590
rect 91006 240272 91062 240281
rect 91006 240207 91062 240216
rect 89732 238726 90404 238754
rect 89732 229770 89760 238726
rect 89720 229764 89772 229770
rect 89720 229706 89772 229712
rect 88984 182844 89036 182850
rect 88984 182786 89036 182792
rect 91020 180130 91048 240207
rect 91100 240168 91152 240174
rect 91100 240110 91152 240116
rect 91112 215286 91140 240110
rect 91204 235278 91232 241590
rect 92216 238754 92244 241726
rect 93766 241703 93822 241712
rect 95344 241748 95976 241754
rect 95344 241742 96028 241748
rect 95344 241726 96016 241742
rect 92308 241590 92368 241618
rect 92920 241602 93256 241618
rect 92920 241596 93268 241602
rect 92920 241590 93216 241596
rect 92308 240174 92336 241590
rect 93216 241538 93268 241544
rect 93320 241590 93472 241618
rect 92296 240168 92348 240174
rect 92296 240110 92348 240116
rect 93320 238754 93348 241590
rect 93780 241233 93808 241703
rect 93872 241590 94024 241618
rect 94148 241590 94576 241618
rect 94792 241590 95128 241618
rect 93766 241224 93822 241233
rect 93766 241159 93822 241168
rect 92216 238726 92336 238754
rect 91192 235272 91244 235278
rect 91192 235214 91244 235220
rect 91100 215280 91152 215286
rect 91100 215222 91152 215228
rect 91100 206304 91152 206310
rect 91100 206246 91152 206252
rect 91112 205698 91140 206246
rect 91100 205692 91152 205698
rect 91100 205634 91152 205640
rect 91008 180124 91060 180130
rect 91008 180066 91060 180072
rect 92308 178702 92336 238726
rect 92492 238726 93348 238754
rect 92492 227730 92520 238726
rect 92480 227724 92532 227730
rect 92480 227666 92532 227672
rect 92492 226370 92520 227666
rect 92480 226364 92532 226370
rect 92480 226306 92532 226312
rect 93124 226364 93176 226370
rect 93124 226306 93176 226312
rect 93136 206310 93164 226306
rect 93872 213314 93900 241590
rect 94148 234025 94176 241590
rect 94792 238754 94820 241590
rect 95240 240168 95292 240174
rect 95240 240110 95292 240116
rect 94240 238726 94820 238754
rect 94240 237561 94268 238726
rect 95148 238672 95200 238678
rect 95148 238614 95200 238620
rect 95160 238105 95188 238614
rect 95146 238096 95202 238105
rect 95146 238031 95202 238040
rect 94226 237552 94282 237561
rect 94226 237487 94282 237496
rect 94688 237448 94740 237454
rect 94688 237390 94740 237396
rect 94134 234016 94190 234025
rect 94134 233951 94190 233960
rect 93860 213308 93912 213314
rect 93860 213250 93912 213256
rect 93124 206304 93176 206310
rect 93124 206246 93176 206252
rect 92388 205692 92440 205698
rect 92388 205634 92440 205640
rect 92296 178696 92348 178702
rect 92296 178638 92348 178644
rect 88982 175944 89038 175953
rect 88982 175879 89038 175888
rect 87142 160103 87198 160112
rect 87604 160132 87656 160138
rect 86972 134966 87046 134994
rect 86052 134694 86480 134722
rect 87018 134708 87046 134966
rect 87156 134722 87184 160103
rect 87604 160074 87656 160080
rect 88248 160132 88300 160138
rect 88248 160074 88300 160080
rect 87616 144906 87644 160074
rect 88340 153944 88392 153950
rect 88340 153886 88392 153892
rect 88352 151814 88380 153886
rect 88352 151786 88656 151814
rect 87604 144900 87656 144906
rect 87604 144842 87656 144848
rect 87616 142154 87644 144842
rect 87616 142126 87736 142154
rect 87708 134722 87736 142126
rect 88524 138712 88576 138718
rect 88524 138654 88576 138660
rect 88340 136604 88392 136610
rect 88340 136546 88392 136552
rect 88352 135930 88380 136546
rect 88340 135924 88392 135930
rect 88340 135866 88392 135872
rect 88536 134994 88564 138654
rect 88628 136066 88656 151786
rect 88996 149190 89024 175879
rect 89720 175296 89772 175302
rect 89720 175238 89772 175244
rect 89628 149796 89680 149802
rect 89628 149738 89680 149744
rect 88984 149184 89036 149190
rect 88984 149126 89036 149132
rect 88708 142180 88760 142186
rect 88708 142122 88760 142128
rect 88720 137290 88748 142122
rect 89166 137320 89222 137329
rect 88708 137284 88760 137290
rect 89166 137255 89222 137264
rect 88708 137226 88760 137232
rect 88616 136060 88668 136066
rect 88616 136002 88668 136008
rect 88490 134966 88564 134994
rect 87156 134694 87584 134722
rect 87708 134694 87952 134722
rect 88490 134708 88518 134966
rect 73066 134671 73122 134680
rect 89180 134586 89208 137255
rect 89640 136610 89668 149738
rect 89732 138106 89760 175238
rect 89810 168464 89866 168473
rect 89810 168399 89866 168408
rect 89720 138100 89772 138106
rect 89720 138042 89772 138048
rect 89628 136604 89680 136610
rect 89628 136546 89680 136552
rect 89260 136060 89312 136066
rect 89260 136002 89312 136008
rect 89272 134722 89300 136002
rect 89824 134722 89852 168399
rect 91744 163532 91796 163538
rect 91744 163474 91796 163480
rect 90180 138100 90232 138106
rect 90180 138042 90232 138048
rect 90192 134722 90220 138042
rect 91192 136604 91244 136610
rect 91192 136546 91244 136552
rect 89272 134694 89608 134722
rect 89824 134694 89976 134722
rect 90192 134694 90528 134722
rect 91204 134586 91232 136546
rect 91756 135425 91784 163474
rect 92400 142154 92428 205634
rect 92478 169824 92534 169833
rect 92478 169759 92534 169768
rect 92308 142126 92428 142154
rect 92308 135425 92336 142126
rect 92388 138100 92440 138106
rect 92388 138042 92440 138048
rect 91742 135416 91798 135425
rect 91742 135351 91798 135360
rect 92294 135416 92350 135425
rect 92294 135351 92350 135360
rect 91756 134722 91784 135351
rect 92400 134722 92428 138042
rect 92492 134994 92520 169759
rect 92664 164892 92716 164898
rect 92664 164834 92716 164840
rect 92572 142860 92624 142866
rect 92572 142802 92624 142808
rect 92584 138106 92612 142802
rect 92572 138100 92624 138106
rect 92572 138042 92624 138048
rect 92492 134966 92566 134994
rect 91632 134694 91784 134722
rect 92184 134694 92428 134722
rect 92538 134708 92566 134966
rect 92676 134722 92704 164834
rect 93136 144809 93164 206246
rect 93860 158772 93912 158778
rect 93860 158714 93912 158720
rect 93872 151814 93900 158714
rect 93872 151786 94360 151814
rect 93122 144800 93178 144809
rect 93122 144735 93178 144744
rect 93216 142248 93268 142254
rect 93216 142190 93268 142196
rect 92676 134694 93104 134722
rect 93228 134638 93256 142190
rect 93768 135992 93820 135998
rect 93768 135934 93820 135940
rect 93780 134722 93808 135934
rect 94228 135924 94280 135930
rect 94228 135866 94280 135872
rect 94240 134858 94268 135866
rect 93656 134694 93808 134722
rect 94194 134830 94268 134858
rect 94194 134708 94222 134830
rect 94332 134722 94360 151786
rect 94332 134694 94576 134722
rect 89056 134558 89208 134586
rect 91080 134558 91232 134586
rect 93216 134632 93268 134638
rect 93216 134574 93268 134580
rect 94700 103514 94728 237390
rect 95148 236020 95200 236026
rect 95148 235962 95200 235968
rect 94780 233708 94832 233714
rect 94780 233650 94832 233656
rect 94792 108769 94820 233650
rect 95160 158778 95188 235962
rect 95252 204950 95280 240110
rect 95344 237454 95372 241726
rect 97722 241632 97778 241641
rect 95896 241590 96232 241618
rect 96784 241590 96936 241618
rect 95896 240174 95924 241590
rect 95884 240168 95936 240174
rect 96908 240145 96936 241590
rect 97000 241590 97336 241618
rect 95884 240110 95936 240116
rect 96894 240136 96950 240145
rect 96894 240071 96950 240080
rect 97000 238754 97028 241590
rect 97888 241590 97948 241618
rect 97722 241567 97724 241576
rect 97776 241567 97778 241576
rect 97724 241538 97776 241544
rect 96632 238726 97028 238754
rect 95332 237448 95384 237454
rect 95332 237390 95384 237396
rect 96528 234660 96580 234666
rect 96528 234602 96580 234608
rect 95240 204944 95292 204950
rect 95240 204886 95292 204892
rect 95884 204944 95936 204950
rect 95884 204886 95936 204892
rect 95148 158772 95200 158778
rect 95148 158714 95200 158720
rect 95700 145580 95752 145586
rect 95700 145522 95752 145528
rect 95712 144974 95740 145522
rect 95424 144968 95476 144974
rect 95424 144910 95476 144916
rect 95700 144968 95752 144974
rect 95700 144910 95752 144916
rect 95238 135552 95294 135561
rect 95238 135487 95294 135496
rect 94872 135312 94924 135318
rect 94872 135254 94924 135260
rect 94884 134570 94912 135254
rect 94872 134564 94924 134570
rect 94872 134506 94924 134512
rect 94778 108760 94834 108769
rect 94778 108695 94834 108704
rect 94700 103486 94820 103514
rect 68664 93826 68968 93854
rect 68388 92886 68416 92917
rect 68376 92880 68428 92886
rect 68428 92828 68816 92834
rect 68376 92822 68816 92828
rect 68388 92806 68816 92822
rect 68388 84194 68416 92806
rect 68940 92750 68968 93826
rect 94688 93560 94740 93566
rect 94392 93508 94688 93514
rect 94392 93502 94740 93508
rect 94392 93486 94728 93502
rect 94792 93242 94820 103486
rect 94872 94512 94924 94518
rect 94872 94454 94924 94460
rect 94700 93214 94820 93242
rect 68928 92744 68980 92750
rect 68928 92686 68980 92692
rect 68296 84166 68416 84194
rect 67824 71732 67876 71738
rect 67824 71674 67876 71680
rect 68296 64802 68324 84166
rect 68284 64796 68336 64802
rect 68284 64738 68336 64744
rect 67270 63472 67326 63481
rect 67270 63407 67326 63416
rect 66904 60036 66956 60042
rect 66904 59978 66956 59984
rect 65524 45552 65576 45558
rect 65524 45494 65576 45500
rect 66168 44872 66220 44878
rect 66168 44814 66220 44820
rect 62028 43444 62080 43450
rect 62028 43386 62080 43392
rect 61660 35216 61712 35222
rect 61660 35158 61712 35164
rect 61936 26920 61988 26926
rect 61936 26862 61988 26868
rect 61948 3534 61976 26862
rect 57244 3528 57296 3534
rect 57244 3470 57296 3476
rect 57888 3528 57940 3534
rect 57888 3470 57940 3476
rect 58440 3528 58492 3534
rect 58440 3470 58492 3476
rect 59268 3528 59320 3534
rect 59268 3470 59320 3476
rect 59636 3528 59688 3534
rect 59636 3470 59688 3476
rect 60648 3528 60700 3534
rect 60648 3470 60700 3476
rect 60832 3528 60884 3534
rect 60832 3470 60884 3476
rect 61936 3528 61988 3534
rect 61936 3470 61988 3476
rect 55128 3052 55180 3058
rect 55128 2994 55180 3000
rect 56048 3052 56100 3058
rect 56048 2994 56100 3000
rect 56060 480 56088 2994
rect 57256 480 57284 3470
rect 58452 480 58480 3470
rect 59648 480 59676 3470
rect 60844 480 60872 3470
rect 62040 480 62068 43386
rect 64788 13116 64840 13122
rect 64788 13058 64840 13064
rect 64800 3534 64828 13058
rect 66180 3534 66208 44814
rect 66720 3596 66772 3602
rect 66720 3538 66772 3544
rect 64328 3528 64380 3534
rect 64328 3470 64380 3476
rect 64788 3528 64840 3534
rect 64788 3470 64840 3476
rect 65524 3528 65576 3534
rect 65524 3470 65576 3476
rect 66168 3528 66220 3534
rect 66168 3470 66220 3476
rect 63222 3360 63278 3369
rect 63222 3295 63278 3304
rect 63236 480 63264 3295
rect 64340 480 64368 3470
rect 65536 480 65564 3470
rect 66732 480 66760 3538
rect 66916 3466 66944 59978
rect 68940 57934 68968 92686
rect 69170 92562 69198 92820
rect 69722 92721 69750 92820
rect 70274 92750 70302 92820
rect 70262 92744 70314 92750
rect 69708 92712 69764 92721
rect 70262 92686 70314 92692
rect 69708 92647 69764 92656
rect 69722 92562 69750 92647
rect 69170 92534 69244 92562
rect 69216 89758 69244 92534
rect 69676 92534 69750 92562
rect 69846 92576 69902 92585
rect 69204 89752 69256 89758
rect 69204 89694 69256 89700
rect 69676 84194 69704 92534
rect 70826 92562 70854 92820
rect 71194 92721 71222 92820
rect 71180 92712 71236 92721
rect 71746 92698 71774 92820
rect 71746 92670 71820 92698
rect 71180 92647 71236 92656
rect 69846 92511 69902 92520
rect 70412 92534 70854 92562
rect 69216 84166 69704 84194
rect 69216 70378 69244 84166
rect 69860 73166 69888 92511
rect 70306 77888 70362 77897
rect 70306 77823 70362 77832
rect 69848 73160 69900 73166
rect 69848 73102 69900 73108
rect 69204 70372 69256 70378
rect 69204 70314 69256 70320
rect 68928 57928 68980 57934
rect 68928 57870 68980 57876
rect 70216 32428 70268 32434
rect 70216 32370 70268 32376
rect 68928 15904 68980 15910
rect 68928 15846 68980 15852
rect 68940 3534 68968 15846
rect 70228 3534 70256 32370
rect 67916 3528 67968 3534
rect 67916 3470 67968 3476
rect 68928 3528 68980 3534
rect 68928 3470 68980 3476
rect 69112 3528 69164 3534
rect 69112 3470 69164 3476
rect 70216 3528 70268 3534
rect 70216 3470 70268 3476
rect 66904 3460 66956 3466
rect 66904 3402 66956 3408
rect 67928 480 67956 3470
rect 69124 480 69152 3470
rect 70320 480 70348 77823
rect 70412 56574 70440 92534
rect 71792 91089 71820 92670
rect 72298 92562 72326 92820
rect 72850 92721 72878 92820
rect 72836 92712 72892 92721
rect 72836 92647 72892 92656
rect 73402 92562 73430 92820
rect 73770 92698 73798 92820
rect 72298 92534 72372 92562
rect 71778 91080 71834 91089
rect 71778 91015 71834 91024
rect 71044 89752 71096 89758
rect 71044 89694 71096 89700
rect 71056 84182 71084 89694
rect 71792 86601 71820 91015
rect 72344 88262 72372 92534
rect 73356 92534 73430 92562
rect 73724 92670 73798 92698
rect 73066 90400 73122 90409
rect 73066 90335 73122 90344
rect 73080 89758 73108 90335
rect 73068 89752 73120 89758
rect 73068 89694 73120 89700
rect 72332 88256 72384 88262
rect 72332 88198 72384 88204
rect 71778 86592 71834 86601
rect 71778 86527 71834 86536
rect 71044 84176 71096 84182
rect 71044 84118 71096 84124
rect 73080 78033 73108 89694
rect 73160 89684 73212 89690
rect 73160 89626 73212 89632
rect 73172 89078 73200 89626
rect 73160 89072 73212 89078
rect 73160 89014 73212 89020
rect 73066 78024 73122 78033
rect 73066 77959 73122 77968
rect 71688 76560 71740 76566
rect 71688 76502 71740 76508
rect 70400 56568 70452 56574
rect 70400 56510 70452 56516
rect 71700 6914 71728 76502
rect 73356 60722 73384 92534
rect 73724 89690 73752 92670
rect 74322 92562 74350 92820
rect 74874 92562 74902 92820
rect 74276 92534 74350 92562
rect 74736 92534 74902 92562
rect 74276 89758 74304 92534
rect 74736 92478 74764 92534
rect 75426 92528 75454 92820
rect 75794 92528 75822 92820
rect 76346 92698 76374 92820
rect 75426 92500 75500 92528
rect 74724 92472 74776 92478
rect 74724 92414 74776 92420
rect 74264 89752 74316 89758
rect 74264 89694 74316 89700
rect 73712 89684 73764 89690
rect 73712 89626 73764 89632
rect 75472 85474 75500 92500
rect 75748 92500 75822 92528
rect 76300 92670 76374 92698
rect 75748 90914 75776 92500
rect 76300 92410 76328 92670
rect 76898 92528 76926 92820
rect 77450 92528 77478 92820
rect 78002 92528 78030 92820
rect 76668 92500 76926 92528
rect 77312 92500 77478 92528
rect 77588 92500 78030 92528
rect 78370 92528 78398 92820
rect 78922 92528 78950 92820
rect 79474 92528 79502 92820
rect 80026 92528 80054 92820
rect 80578 92528 80606 92820
rect 78370 92500 78444 92528
rect 78922 92500 78996 92528
rect 79474 92500 79548 92528
rect 80026 92500 80100 92528
rect 76288 92404 76340 92410
rect 76288 92346 76340 92352
rect 75736 90908 75788 90914
rect 75736 90850 75788 90856
rect 75460 85468 75512 85474
rect 75460 85410 75512 85416
rect 76668 84194 76696 92500
rect 76024 84166 76696 84194
rect 76024 82754 76052 84166
rect 76012 82748 76064 82754
rect 76012 82690 76064 82696
rect 77312 80073 77340 92500
rect 77588 81297 77616 92500
rect 78416 89729 78444 92500
rect 78968 90982 78996 92500
rect 78956 90976 79008 90982
rect 78956 90918 79008 90924
rect 78402 89720 78458 89729
rect 78402 89655 78458 89664
rect 77944 89072 77996 89078
rect 77944 89014 77996 89020
rect 77574 81288 77630 81297
rect 77574 81223 77630 81232
rect 77298 80064 77354 80073
rect 77298 79999 77354 80008
rect 77956 75886 77984 89014
rect 79520 85377 79548 92500
rect 79506 85368 79562 85377
rect 79506 85303 79562 85312
rect 80072 84114 80100 92500
rect 80164 92500 80606 92528
rect 80946 92528 80974 92820
rect 81498 92528 81526 92820
rect 81624 92608 81676 92614
rect 81624 92550 81676 92556
rect 80946 92500 81020 92528
rect 80060 84108 80112 84114
rect 80060 84050 80112 84056
rect 80164 81326 80192 92500
rect 80992 86970 81020 92500
rect 81452 92500 81526 92528
rect 81452 92449 81480 92500
rect 81438 92440 81494 92449
rect 81438 92375 81494 92384
rect 80980 86964 81032 86970
rect 80980 86906 81032 86912
rect 80152 81320 80204 81326
rect 80152 81262 80204 81268
rect 81636 77246 81664 92550
rect 82050 92528 82078 92820
rect 82602 92614 82630 92820
rect 82590 92608 82642 92614
rect 82590 92550 82642 92556
rect 82970 92528 82998 92820
rect 81728 92500 82078 92528
rect 82832 92500 82998 92528
rect 83522 92528 83550 92820
rect 84074 92528 84102 92820
rect 84626 92698 84654 92820
rect 84626 92670 84700 92698
rect 83522 92500 83596 92528
rect 84074 92500 84148 92528
rect 81728 79966 81756 92500
rect 82832 82521 82860 92500
rect 83568 92313 83596 92500
rect 83554 92304 83610 92313
rect 83554 92239 83610 92248
rect 84120 89457 84148 92500
rect 84672 91050 84700 92670
rect 85178 92528 85206 92820
rect 84948 92500 85206 92528
rect 85546 92528 85574 92820
rect 86098 92528 86126 92820
rect 86650 92528 86678 92820
rect 87202 92698 87230 92820
rect 87202 92670 87276 92698
rect 85546 92500 85620 92528
rect 86098 92500 86172 92528
rect 86650 92500 86724 92528
rect 84660 91044 84712 91050
rect 84660 90986 84712 90992
rect 84106 89448 84162 89457
rect 84106 89383 84162 89392
rect 84948 84194 84976 92500
rect 85592 92410 85620 92500
rect 85580 92404 85632 92410
rect 85580 92346 85632 92352
rect 86144 86873 86172 92500
rect 86696 88097 86724 92500
rect 86682 88088 86738 88097
rect 86682 88023 86738 88032
rect 86130 86864 86186 86873
rect 86130 86799 86186 86808
rect 87248 85542 87276 92670
rect 87570 92528 87598 92820
rect 87340 92500 87598 92528
rect 88122 92528 88150 92820
rect 88674 92750 88702 92820
rect 88662 92744 88714 92750
rect 88662 92686 88714 92692
rect 88674 92562 88702 92686
rect 88674 92534 88748 92562
rect 88122 92500 88196 92528
rect 87236 85536 87288 85542
rect 87236 85478 87288 85484
rect 87340 84194 87368 92500
rect 88168 92410 88196 92500
rect 88156 92404 88208 92410
rect 88156 92346 88208 92352
rect 88720 89622 88748 92534
rect 89226 92528 89254 92820
rect 89778 92528 89806 92820
rect 89904 92608 89956 92614
rect 89904 92550 89956 92556
rect 89226 92500 89300 92528
rect 89778 92500 89852 92528
rect 89272 89690 89300 92500
rect 89260 89684 89312 89690
rect 89260 89626 89312 89632
rect 88708 89616 88760 89622
rect 88708 89558 88760 89564
rect 89536 89616 89588 89622
rect 89536 89558 89588 89564
rect 87604 89004 87656 89010
rect 87604 88946 87656 88952
rect 84212 84166 84976 84194
rect 86972 84166 87368 84194
rect 82818 82512 82874 82521
rect 82818 82447 82874 82456
rect 81716 79960 81768 79966
rect 81716 79902 81768 79908
rect 81624 77240 81676 77246
rect 81624 77182 81676 77188
rect 77944 75880 77996 75886
rect 77944 75822 77996 75828
rect 75826 75168 75882 75177
rect 75826 75103 75882 75112
rect 73344 60716 73396 60722
rect 73344 60658 73396 60664
rect 73068 53100 73120 53106
rect 73068 53042 73120 53048
rect 71516 6886 71728 6914
rect 71516 480 71544 6886
rect 73080 3534 73108 53042
rect 73802 6216 73858 6225
rect 73802 6151 73858 6160
rect 72608 3528 72660 3534
rect 72608 3470 72660 3476
rect 73068 3528 73120 3534
rect 73068 3470 73120 3476
rect 72620 480 72648 3470
rect 73816 480 73844 6151
rect 75840 3534 75868 75103
rect 84212 74526 84240 84166
rect 84200 74520 84252 74526
rect 84200 74462 84252 74468
rect 76562 73808 76618 73817
rect 76562 73743 76618 73752
rect 76576 3602 76604 73743
rect 86868 68332 86920 68338
rect 86868 68274 86920 68280
rect 84106 61432 84162 61441
rect 84106 61367 84162 61376
rect 79968 42084 80020 42090
rect 79968 42026 80020 42032
rect 77208 40724 77260 40730
rect 77208 40666 77260 40672
rect 76564 3596 76616 3602
rect 76564 3538 76616 3544
rect 77220 3534 77248 40666
rect 78588 17264 78640 17270
rect 78588 17206 78640 17212
rect 75000 3528 75052 3534
rect 75000 3470 75052 3476
rect 75828 3528 75880 3534
rect 75828 3470 75880 3476
rect 76196 3528 76248 3534
rect 76196 3470 76248 3476
rect 77208 3528 77260 3534
rect 77208 3470 77260 3476
rect 75012 480 75040 3470
rect 76208 480 76236 3470
rect 77392 3392 77444 3398
rect 77392 3334 77444 3340
rect 77404 480 77432 3334
rect 78600 480 78628 17206
rect 79980 6914 80008 42026
rect 84016 24132 84068 24138
rect 84016 24074 84068 24080
rect 81346 14512 81402 14521
rect 81346 14447 81402 14456
rect 79704 6886 80008 6914
rect 79704 480 79732 6886
rect 81360 3534 81388 14447
rect 82084 8968 82136 8974
rect 82084 8910 82136 8916
rect 80888 3528 80940 3534
rect 80888 3470 80940 3476
rect 81348 3528 81400 3534
rect 81348 3470 81400 3476
rect 80900 480 80928 3470
rect 82096 480 82124 8910
rect 84028 3466 84056 24074
rect 83280 3460 83332 3466
rect 83280 3402 83332 3408
rect 84016 3460 84068 3466
rect 84016 3402 84068 3408
rect 83292 480 83320 3402
rect 84120 2802 84148 61367
rect 86776 21412 86828 21418
rect 86776 21354 86828 21360
rect 86788 16574 86816 21354
rect 86696 16546 86816 16574
rect 85672 3596 85724 3602
rect 85672 3538 85724 3544
rect 84120 2774 84516 2802
rect 84488 480 84516 2774
rect 85684 480 85712 3538
rect 86696 3482 86724 16546
rect 86880 6914 86908 68274
rect 86972 66230 87000 84166
rect 87616 81394 87644 88946
rect 87604 81388 87656 81394
rect 87604 81330 87656 81336
rect 86960 66224 87012 66230
rect 86960 66166 87012 66172
rect 89548 62082 89576 89558
rect 89824 86902 89852 92500
rect 89812 86896 89864 86902
rect 89812 86838 89864 86844
rect 89916 77217 89944 92550
rect 90146 92528 90174 92820
rect 90698 92614 90726 92820
rect 90686 92608 90738 92614
rect 90686 92550 90738 92556
rect 91250 92528 91278 92820
rect 91802 92721 91830 92820
rect 91788 92712 91844 92721
rect 91788 92647 91844 92656
rect 90008 92500 90174 92528
rect 91112 92500 91278 92528
rect 92354 92528 92382 92820
rect 92722 92528 92750 92820
rect 93274 92721 93302 92820
rect 93260 92712 93316 92721
rect 93260 92647 93316 92656
rect 93274 92528 93302 92647
rect 93826 92562 93854 92820
rect 94700 92562 94728 93214
rect 94778 93120 94834 93129
rect 94778 93055 94834 93064
rect 93826 92534 94728 92562
rect 92354 92500 92428 92528
rect 92722 92500 92796 92528
rect 93274 92500 93348 92528
rect 90008 82657 90036 92500
rect 91112 84153 91140 92500
rect 92400 92177 92428 92500
rect 92386 92168 92442 92177
rect 92386 92103 92442 92112
rect 92768 88233 92796 92500
rect 93122 91760 93178 91769
rect 93122 91695 93178 91704
rect 92754 88224 92810 88233
rect 92754 88159 92810 88168
rect 91098 84144 91154 84153
rect 91098 84079 91154 84088
rect 89994 82648 90050 82657
rect 89994 82583 90050 82592
rect 89902 77208 89958 77217
rect 89902 77143 89958 77152
rect 91006 72448 91062 72457
rect 91006 72383 91062 72392
rect 89628 71052 89680 71058
rect 89628 70994 89680 71000
rect 89536 62076 89588 62082
rect 89536 62018 89588 62024
rect 88246 48920 88302 48929
rect 88246 48855 88302 48864
rect 88260 6914 88288 48855
rect 86788 6886 86908 6914
rect 87984 6886 88288 6914
rect 86788 3602 86816 6886
rect 86776 3596 86828 3602
rect 86776 3538 86828 3544
rect 86696 3454 86908 3482
rect 86880 480 86908 3454
rect 87984 480 88012 6886
rect 89640 3534 89668 70994
rect 90916 11756 90968 11762
rect 90916 11698 90968 11704
rect 90928 3534 90956 11698
rect 91020 3534 91048 72383
rect 93136 20670 93164 91695
rect 93320 84194 93348 92500
rect 93872 84194 93900 92534
rect 94792 87961 94820 93055
rect 94884 92410 94912 94454
rect 95148 93152 95200 93158
rect 95148 93094 95200 93100
rect 95160 92478 95188 93094
rect 95252 92818 95280 135487
rect 95436 127673 95464 144910
rect 95422 127664 95478 127673
rect 95422 127599 95478 127608
rect 95330 120320 95386 120329
rect 95330 120255 95386 120264
rect 95240 92812 95292 92818
rect 95240 92754 95292 92760
rect 95148 92472 95200 92478
rect 95148 92414 95200 92420
rect 94872 92404 94924 92410
rect 94872 92346 94924 92352
rect 95148 91112 95200 91118
rect 95148 91054 95200 91060
rect 94778 87952 94834 87961
rect 94778 87887 94834 87896
rect 95160 86873 95188 91054
rect 95146 86864 95202 86873
rect 95146 86799 95202 86808
rect 93320 84166 93808 84194
rect 93872 84166 94544 84194
rect 93780 64870 93808 84166
rect 94516 67522 94544 84166
rect 95344 83473 95372 120255
rect 95896 93566 95924 204886
rect 96540 98297 96568 234602
rect 96632 211138 96660 238726
rect 97920 231810 97948 241590
rect 97264 231804 97316 231810
rect 97264 231746 97316 231752
rect 97908 231804 97960 231810
rect 97908 231746 97960 231752
rect 97276 230586 97304 231746
rect 97264 230580 97316 230586
rect 97264 230522 97316 230528
rect 96620 211132 96672 211138
rect 96620 211074 96672 211080
rect 97276 207670 97304 230522
rect 97264 207664 97316 207670
rect 97264 207606 97316 207612
rect 96804 137284 96856 137290
rect 96804 137226 96856 137232
rect 96710 135960 96766 135969
rect 96710 135895 96766 135904
rect 96620 133204 96672 133210
rect 96620 133146 96672 133152
rect 96632 132297 96660 133146
rect 96724 133113 96752 135895
rect 96710 133104 96766 133113
rect 96710 133039 96766 133048
rect 96712 132388 96764 132394
rect 96712 132330 96764 132336
rect 96618 132288 96674 132297
rect 96618 132223 96674 132232
rect 96724 131481 96752 132330
rect 96710 131472 96766 131481
rect 96710 131407 96766 131416
rect 96710 130928 96766 130937
rect 96710 130863 96766 130872
rect 96620 130620 96672 130626
rect 96620 130562 96672 130568
rect 96632 130121 96660 130562
rect 96724 130422 96752 130863
rect 96712 130416 96764 130422
rect 96712 130358 96764 130364
rect 96618 130112 96674 130121
rect 96618 130047 96674 130056
rect 96724 129826 96752 130358
rect 96632 129798 96752 129826
rect 96526 98288 96582 98297
rect 96526 98223 96582 98232
rect 95884 93560 95936 93566
rect 95884 93502 95936 93508
rect 96632 91769 96660 129798
rect 96712 129736 96764 129742
rect 96712 129678 96764 129684
rect 96724 129305 96752 129678
rect 96710 129296 96766 129305
rect 96710 129231 96766 129240
rect 96816 128354 96844 137226
rect 96724 128326 96844 128354
rect 96724 125497 96752 128326
rect 96710 125488 96766 125497
rect 96710 125423 96766 125432
rect 97172 120080 97224 120086
rect 97172 120022 97224 120028
rect 97184 119513 97212 120022
rect 97170 119504 97226 119513
rect 97170 119439 97226 119448
rect 97172 115728 97224 115734
rect 97170 115696 97172 115705
rect 97224 115696 97226 115705
rect 97170 115631 97226 115640
rect 96712 111920 96764 111926
rect 96710 111888 96712 111897
rect 96764 111888 96766 111897
rect 96710 111823 96766 111832
rect 96712 111784 96764 111790
rect 96712 111726 96764 111732
rect 96724 111081 96752 111726
rect 96710 111072 96766 111081
rect 96710 111007 96766 111016
rect 97080 110288 97132 110294
rect 97078 110256 97080 110265
rect 97132 110256 97134 110265
rect 97078 110191 97134 110200
rect 96804 106276 96856 106282
rect 96804 106218 96856 106224
rect 96816 105097 96844 106218
rect 96802 105088 96858 105097
rect 96802 105023 96858 105032
rect 96712 102128 96764 102134
rect 96710 102096 96712 102105
rect 96764 102096 96766 102105
rect 96710 102031 96766 102040
rect 96712 101856 96764 101862
rect 96712 101798 96764 101804
rect 96724 101289 96752 101798
rect 96710 101280 96766 101289
rect 96710 101215 96766 101224
rect 96712 96892 96764 96898
rect 96712 96834 96764 96840
rect 96724 96665 96752 96834
rect 96710 96656 96766 96665
rect 96710 96591 96766 96600
rect 97276 95033 97304 207606
rect 97356 184272 97408 184278
rect 97356 184214 97408 184220
rect 97368 137358 97396 184214
rect 97448 144900 97500 144906
rect 97448 144842 97500 144848
rect 97356 137352 97408 137358
rect 97356 137294 97408 137300
rect 97460 123321 97488 144842
rect 97632 128308 97684 128314
rect 97632 128250 97684 128256
rect 97644 127129 97672 128250
rect 97630 127120 97686 127129
rect 97630 127055 97686 127064
rect 97908 126948 97960 126954
rect 97908 126890 97960 126896
rect 97920 126313 97948 126890
rect 97906 126304 97962 126313
rect 97906 126239 97962 126248
rect 97816 125588 97868 125594
rect 97816 125530 97868 125536
rect 97828 124681 97856 125530
rect 97908 125520 97960 125526
rect 97906 125488 97908 125497
rect 97960 125488 97962 125497
rect 97906 125423 97962 125432
rect 97814 124672 97870 124681
rect 97814 124607 97870 124616
rect 97908 124160 97960 124166
rect 97906 124128 97908 124137
rect 97960 124128 97962 124137
rect 97906 124063 97962 124072
rect 97722 123448 97778 123457
rect 97722 123383 97778 123392
rect 97446 123312 97502 123321
rect 97446 123247 97502 123256
rect 97448 122732 97500 122738
rect 97448 122674 97500 122680
rect 97460 121689 97488 122674
rect 97446 121680 97502 121689
rect 97446 121615 97502 121624
rect 97540 121440 97592 121446
rect 97540 121382 97592 121388
rect 97552 120329 97580 121382
rect 97632 121100 97684 121106
rect 97632 121042 97684 121048
rect 97644 120873 97672 121042
rect 97630 120864 97686 120873
rect 97630 120799 97686 120808
rect 97538 120320 97594 120329
rect 97538 120255 97594 120264
rect 97354 116648 97410 116657
rect 97354 116583 97410 116592
rect 97368 114073 97396 116583
rect 97736 116521 97764 123383
rect 97908 122800 97960 122806
rect 97908 122742 97960 122748
rect 97920 122505 97948 122742
rect 97906 122496 97962 122505
rect 97906 122431 97962 122440
rect 97906 118688 97962 118697
rect 97816 118652 97868 118658
rect 97906 118623 97962 118632
rect 97816 118594 97868 118600
rect 97828 117881 97856 118594
rect 97920 118590 97948 118623
rect 97908 118584 97960 118590
rect 97908 118526 97960 118532
rect 97814 117872 97870 117881
rect 97814 117807 97870 117816
rect 97908 117292 97960 117298
rect 97908 117234 97960 117240
rect 97920 117065 97948 117234
rect 97906 117056 97962 117065
rect 97906 116991 97962 117000
rect 97722 116512 97778 116521
rect 97722 116447 97778 116456
rect 97540 115932 97592 115938
rect 97540 115874 97592 115880
rect 97552 114889 97580 115874
rect 97538 114880 97594 114889
rect 97538 114815 97594 114824
rect 97354 114064 97410 114073
rect 97354 113999 97410 114008
rect 97262 95024 97318 95033
rect 97262 94959 97318 94968
rect 96986 94480 97042 94489
rect 96986 94415 97042 94424
rect 96618 91760 96674 91769
rect 96618 91695 96674 91704
rect 97000 88262 97028 94415
rect 96988 88256 97040 88262
rect 96988 88198 97040 88204
rect 95330 83464 95386 83473
rect 95330 83399 95386 83408
rect 97368 78606 97396 113999
rect 97538 113520 97594 113529
rect 97538 113455 97594 113464
rect 97552 113218 97580 113455
rect 97540 113212 97592 113218
rect 97540 113154 97592 113160
rect 97906 112704 97962 112713
rect 97906 112639 97962 112648
rect 97920 111858 97948 112639
rect 97908 111852 97960 111858
rect 97908 111794 97960 111800
rect 97908 110424 97960 110430
rect 97908 110366 97960 110372
rect 97920 109721 97948 110366
rect 97906 109712 97962 109721
rect 97906 109647 97962 109656
rect 98012 108118 98040 243510
rect 98104 213926 98132 258431
rect 98196 236026 98224 273226
rect 100036 269793 100064 291887
rect 100114 287464 100170 287473
rect 100114 287399 100170 287408
rect 100022 269784 100078 269793
rect 100022 269719 100078 269728
rect 100128 267889 100156 287399
rect 100298 284880 100354 284889
rect 100298 284815 100354 284824
rect 100312 268433 100340 284815
rect 100760 282736 100812 282742
rect 100758 282704 100760 282713
rect 100812 282704 100814 282713
rect 100758 282639 100814 282648
rect 100760 281512 100812 281518
rect 100760 281454 100812 281460
rect 100772 280265 100800 281454
rect 100850 281072 100906 281081
rect 100850 281007 100906 281016
rect 100758 280256 100814 280265
rect 100864 280226 100892 281007
rect 100758 280191 100814 280200
rect 100852 280220 100904 280226
rect 100852 280162 100904 280168
rect 100760 280152 100812 280158
rect 100760 280094 100812 280100
rect 100772 279449 100800 280094
rect 100758 279440 100814 279449
rect 100758 279375 100814 279384
rect 100760 278656 100812 278662
rect 100760 278598 100812 278604
rect 100772 277817 100800 278598
rect 100758 277808 100814 277817
rect 100758 277743 100814 277752
rect 100760 277296 100812 277302
rect 100760 277238 100812 277244
rect 100772 276185 100800 277238
rect 100850 276720 100906 276729
rect 100850 276655 100906 276664
rect 100758 276176 100814 276185
rect 100758 276111 100814 276120
rect 100760 274644 100812 274650
rect 100760 274586 100812 274592
rect 100772 273737 100800 274586
rect 100758 273728 100814 273737
rect 100758 273663 100814 273672
rect 100760 273216 100812 273222
rect 100760 273158 100812 273164
rect 100772 272921 100800 273158
rect 100758 272912 100814 272921
rect 100758 272847 100814 272856
rect 100864 272105 100892 276655
rect 100850 272096 100906 272105
rect 100850 272031 100906 272040
rect 100760 271856 100812 271862
rect 100760 271798 100812 271804
rect 100772 271289 100800 271798
rect 100758 271280 100814 271289
rect 100680 271238 100758 271266
rect 100298 268424 100354 268433
rect 100298 268359 100354 268368
rect 100114 267880 100170 267889
rect 100114 267815 100170 267824
rect 99286 258224 99342 258233
rect 99286 258159 99342 258168
rect 99196 249756 99248 249762
rect 99196 249698 99248 249704
rect 99208 248441 99236 249698
rect 99194 248432 99250 248441
rect 99194 248367 99250 248376
rect 98274 248296 98330 248305
rect 98274 248231 98330 248240
rect 98288 243574 98316 248231
rect 98276 243568 98328 243574
rect 98276 243510 98328 243516
rect 98440 241590 98776 241618
rect 98748 240145 98776 241590
rect 98734 240136 98790 240145
rect 98734 240071 98790 240080
rect 98184 236020 98236 236026
rect 98184 235962 98236 235968
rect 98092 213920 98144 213926
rect 98092 213862 98144 213868
rect 98736 213920 98788 213926
rect 98736 213862 98788 213868
rect 98748 213246 98776 213862
rect 98736 213240 98788 213246
rect 98736 213182 98788 213188
rect 98644 208412 98696 208418
rect 98644 208354 98696 208360
rect 98000 108112 98052 108118
rect 98000 108054 98052 108060
rect 97906 107264 97962 107273
rect 97906 107199 97962 107208
rect 97920 106418 97948 107199
rect 97908 106412 97960 106418
rect 97908 106354 97960 106360
rect 98000 105596 98052 105602
rect 98000 105538 98052 105544
rect 97906 104272 97962 104281
rect 98012 104258 98040 105538
rect 97962 104230 98040 104258
rect 97906 104207 97962 104216
rect 97908 103488 97960 103494
rect 97814 103456 97870 103465
rect 97908 103430 97960 103436
rect 97814 103391 97816 103400
rect 97868 103391 97870 103400
rect 97816 103362 97868 103368
rect 97920 102921 97948 103430
rect 97906 102912 97962 102921
rect 97906 102847 97962 102856
rect 97446 100464 97502 100473
rect 97446 100399 97502 100408
rect 97460 78674 97488 100399
rect 97906 99648 97962 99657
rect 97906 99583 97962 99592
rect 97920 99414 97948 99583
rect 97908 99408 97960 99414
rect 97908 99350 97960 99356
rect 97906 99104 97962 99113
rect 97906 99039 97908 99048
rect 97960 99039 97962 99048
rect 97908 99010 97960 99016
rect 97906 98288 97962 98297
rect 97906 98223 97962 98232
rect 97920 98190 97948 98223
rect 97908 98184 97960 98190
rect 97908 98126 97960 98132
rect 98656 96898 98684 208354
rect 98748 111926 98776 213182
rect 99194 179480 99250 179489
rect 99194 179415 99196 179424
rect 99248 179415 99250 179424
rect 99196 179386 99248 179392
rect 99300 146334 99328 258159
rect 100114 257408 100170 257417
rect 100114 257343 100170 257352
rect 100022 251152 100078 251161
rect 100022 251087 100078 251096
rect 99380 202836 99432 202842
rect 99380 202778 99432 202784
rect 99392 202162 99420 202778
rect 99380 202156 99432 202162
rect 99380 202098 99432 202104
rect 98828 146328 98880 146334
rect 98828 146270 98880 146276
rect 99288 146328 99340 146334
rect 99288 146270 99340 146276
rect 98736 111920 98788 111926
rect 98736 111862 98788 111868
rect 98840 111790 98868 146270
rect 98828 111784 98880 111790
rect 98828 111726 98880 111732
rect 98736 111172 98788 111178
rect 98736 111114 98788 111120
rect 98644 96892 98696 96898
rect 98644 96834 98696 96840
rect 97814 96112 97870 96121
rect 97814 96047 97870 96056
rect 97828 95334 97856 96047
rect 97816 95328 97868 95334
rect 97816 95270 97868 95276
rect 97906 95296 97962 95305
rect 97906 95231 97908 95240
rect 97960 95231 97962 95240
rect 97908 95202 97960 95208
rect 97908 93696 97960 93702
rect 97906 93664 97908 93673
rect 97960 93664 97962 93673
rect 97906 93599 97962 93608
rect 98748 82657 98776 111114
rect 98920 108112 98972 108118
rect 98920 108054 98972 108060
rect 98932 107710 98960 108054
rect 98920 107704 98972 107710
rect 98920 107646 98972 107652
rect 98932 102134 98960 107646
rect 98920 102128 98972 102134
rect 98920 102070 98972 102076
rect 99392 101862 99420 202098
rect 100036 106282 100064 251087
rect 100128 220114 100156 257343
rect 100206 247616 100262 247625
rect 100206 247551 100262 247560
rect 100116 220108 100168 220114
rect 100116 220050 100168 220056
rect 100128 110294 100156 220050
rect 100220 214606 100248 247551
rect 100208 214600 100260 214606
rect 100208 214542 100260 214548
rect 100220 202842 100248 214542
rect 100208 202836 100260 202842
rect 100208 202778 100260 202784
rect 100680 164286 100708 271238
rect 100758 271215 100814 271224
rect 100760 270496 100812 270502
rect 100758 270464 100760 270473
rect 100812 270464 100814 270473
rect 100758 270399 100814 270408
rect 100760 269068 100812 269074
rect 100760 269010 100812 269016
rect 100772 268841 100800 269010
rect 100758 268832 100814 268841
rect 100758 268767 100814 268776
rect 100760 268388 100812 268394
rect 100760 268330 100812 268336
rect 100772 268025 100800 268330
rect 100758 268016 100814 268025
rect 100758 267951 100814 267960
rect 100758 267200 100814 267209
rect 100758 267135 100814 267144
rect 100772 267034 100800 267135
rect 100760 267028 100812 267034
rect 100760 266970 100812 266976
rect 100942 266384 100998 266393
rect 100942 266319 100998 266328
rect 100758 265568 100814 265577
rect 100758 265503 100814 265512
rect 100772 264994 100800 265503
rect 100760 264988 100812 264994
rect 100760 264930 100812 264936
rect 100850 264752 100906 264761
rect 100850 264687 100906 264696
rect 100758 263936 100814 263945
rect 100758 263871 100814 263880
rect 100772 263634 100800 263871
rect 100864 263702 100892 264687
rect 100852 263696 100904 263702
rect 100852 263638 100904 263644
rect 100760 263628 100812 263634
rect 100760 263570 100812 263576
rect 100758 263120 100814 263129
rect 100758 263055 100814 263064
rect 100772 262886 100800 263055
rect 100760 262880 100812 262886
rect 100956 262857 100984 266319
rect 100760 262822 100812 262828
rect 100942 262848 100998 262857
rect 100772 262426 100800 262822
rect 100942 262783 100998 262792
rect 100772 262398 100984 262426
rect 100758 262304 100814 262313
rect 100758 262239 100760 262248
rect 100812 262239 100814 262248
rect 100760 262210 100812 262216
rect 100852 262200 100904 262206
rect 100852 262142 100904 262148
rect 100864 261497 100892 262142
rect 100850 261488 100906 261497
rect 100850 261423 100906 261432
rect 100850 260672 100906 260681
rect 100850 260607 100906 260616
rect 100758 259856 100814 259865
rect 100758 259791 100814 259800
rect 100772 259554 100800 259791
rect 100760 259548 100812 259554
rect 100760 259490 100812 259496
rect 100864 259486 100892 260607
rect 100852 259480 100904 259486
rect 100852 259422 100904 259428
rect 100956 258074 100984 262398
rect 101416 258233 101444 369106
rect 101508 277001 101536 384231
rect 102060 371210 102088 389127
rect 102782 388512 102838 388521
rect 102782 388447 102838 388456
rect 102048 371204 102100 371210
rect 102048 371146 102100 371152
rect 102690 320240 102746 320249
rect 102690 320175 102746 320184
rect 102704 320074 102732 320175
rect 102692 320068 102744 320074
rect 102692 320010 102744 320016
rect 101588 316736 101640 316742
rect 101588 316678 101640 316684
rect 101494 276992 101550 277001
rect 101494 276927 101550 276936
rect 101494 274544 101550 274553
rect 101494 274479 101550 274488
rect 101508 265674 101536 274479
rect 101600 269657 101628 316678
rect 101678 304192 101734 304201
rect 101678 304127 101734 304136
rect 101692 278633 101720 304127
rect 102796 293962 102824 388447
rect 103164 385694 103192 390374
rect 103900 389337 103928 390374
rect 103886 389328 103942 389337
rect 103886 389263 103942 389272
rect 104164 387796 104216 387802
rect 104164 387738 104216 387744
rect 103152 385688 103204 385694
rect 103152 385630 103204 385636
rect 103520 359508 103572 359514
rect 103520 359450 103572 359456
rect 102876 329860 102928 329866
rect 102876 329802 102928 329808
rect 102140 293956 102192 293962
rect 102140 293898 102192 293904
rect 102784 293956 102836 293962
rect 102784 293898 102836 293904
rect 102152 293350 102180 293898
rect 102140 293344 102192 293350
rect 102140 293286 102192 293292
rect 102138 285696 102194 285705
rect 102138 285631 102194 285640
rect 101678 278624 101734 278633
rect 101678 278559 101734 278568
rect 101586 269648 101642 269657
rect 101586 269583 101642 269592
rect 101496 265668 101548 265674
rect 101496 265610 101548 265616
rect 101680 258732 101732 258738
rect 101680 258674 101732 258680
rect 101402 258224 101458 258233
rect 101402 258159 101458 258168
rect 100772 258046 100984 258074
rect 100208 164280 100260 164286
rect 100208 164222 100260 164228
rect 100668 164280 100720 164286
rect 100668 164222 100720 164228
rect 100220 144906 100248 164222
rect 100208 144900 100260 144906
rect 100208 144842 100260 144848
rect 100772 115734 100800 258046
rect 100850 256592 100906 256601
rect 100850 256527 100906 256536
rect 100864 255406 100892 256527
rect 101402 255776 101458 255785
rect 101402 255711 101458 255720
rect 100852 255400 100904 255406
rect 100852 255342 100904 255348
rect 100852 254992 100904 254998
rect 100850 254960 100852 254969
rect 100904 254960 100906 254969
rect 100850 254895 100906 254904
rect 100850 254144 100906 254153
rect 100850 254079 100906 254088
rect 100864 253978 100892 254079
rect 100852 253972 100904 253978
rect 100852 253914 100904 253920
rect 100850 253328 100906 253337
rect 100850 253263 100906 253272
rect 100864 252618 100892 253263
rect 100852 252612 100904 252618
rect 100852 252554 100904 252560
rect 100852 251048 100904 251054
rect 100852 250990 100904 250996
rect 100864 250889 100892 250990
rect 100850 250880 100906 250889
rect 100850 250815 100906 250824
rect 100850 249248 100906 249257
rect 100850 249183 100906 249192
rect 100864 249082 100892 249183
rect 100852 249076 100904 249082
rect 100852 249018 100904 249024
rect 100850 246800 100906 246809
rect 100850 246735 100906 246744
rect 100864 246362 100892 246735
rect 100852 246356 100904 246362
rect 100852 246298 100904 246304
rect 100850 245984 100906 245993
rect 100850 245919 100906 245928
rect 100864 245682 100892 245919
rect 100852 245676 100904 245682
rect 100852 245618 100904 245624
rect 100850 245168 100906 245177
rect 100850 245103 100906 245112
rect 100864 245002 100892 245103
rect 100852 244996 100904 245002
rect 100852 244938 100904 244944
rect 100942 244352 100998 244361
rect 100942 244287 100998 244296
rect 100850 243536 100906 243545
rect 100850 243471 100906 243480
rect 100864 242962 100892 243471
rect 100852 242956 100904 242962
rect 100852 242898 100904 242904
rect 100956 238754 100984 244287
rect 101416 240174 101444 255711
rect 101692 252521 101720 258674
rect 101678 252512 101734 252521
rect 101678 252447 101734 252456
rect 101956 250504 102008 250510
rect 101956 250446 102008 250452
rect 101968 250073 101996 250446
rect 101954 250064 102010 250073
rect 101954 249999 102010 250008
rect 101968 248414 101996 249999
rect 101968 248386 102088 248414
rect 101404 240168 101456 240174
rect 101404 240110 101456 240116
rect 100864 238726 100984 238754
rect 100864 234666 100892 238726
rect 100852 234660 100904 234666
rect 100852 234602 100904 234608
rect 101416 233714 101444 240110
rect 101404 233708 101456 233714
rect 101404 233650 101456 233656
rect 100852 137352 100904 137358
rect 100852 137294 100904 137300
rect 100760 115728 100812 115734
rect 100760 115670 100812 115676
rect 100116 110288 100168 110294
rect 100116 110230 100168 110236
rect 100116 106956 100168 106962
rect 100116 106898 100168 106904
rect 100024 106276 100076 106282
rect 100024 106218 100076 106224
rect 99380 101856 99432 101862
rect 99380 101798 99432 101804
rect 98828 100768 98880 100774
rect 98828 100710 98880 100716
rect 98840 89593 98868 100710
rect 100024 97300 100076 97306
rect 100024 97242 100076 97248
rect 98826 89584 98882 89593
rect 98826 89519 98882 89528
rect 100036 86737 100064 97242
rect 100128 88097 100156 106898
rect 100760 99068 100812 99074
rect 100760 99010 100812 99016
rect 100772 98705 100800 99010
rect 100758 98696 100814 98705
rect 100758 98631 100814 98640
rect 100864 91050 100892 137294
rect 101404 111104 101456 111110
rect 101404 111046 101456 111052
rect 100852 91044 100904 91050
rect 100852 90986 100904 90992
rect 101416 88330 101444 111046
rect 102060 103562 102088 248386
rect 102152 210458 102180 285631
rect 102888 282742 102916 329802
rect 102968 294092 103020 294098
rect 102968 294034 103020 294040
rect 102980 285705 103008 294034
rect 102966 285696 103022 285705
rect 102966 285631 103022 285640
rect 102876 282736 102928 282742
rect 102876 282678 102928 282684
rect 102784 247104 102836 247110
rect 102784 247046 102836 247052
rect 102322 242720 102378 242729
rect 102322 242655 102378 242664
rect 102230 241632 102286 241641
rect 102230 241567 102232 241576
rect 102284 241567 102286 241576
rect 102232 241538 102284 241544
rect 102336 238754 102364 242655
rect 102244 238726 102364 238754
rect 102140 210452 102192 210458
rect 102140 210394 102192 210400
rect 102244 209778 102272 238726
rect 102796 238649 102824 247046
rect 102782 238640 102838 238649
rect 102782 238575 102838 238584
rect 103532 235929 103560 359450
rect 104176 358766 104204 387738
rect 104544 383654 104572 390646
rect 107750 390688 107806 390697
rect 105138 390646 105216 390674
rect 107640 390646 107750 390674
rect 105082 390623 105138 390632
rect 105188 389065 105216 390646
rect 111982 390688 112038 390697
rect 107806 390646 107976 390674
rect 107750 390623 107806 390632
rect 105266 390552 105322 390561
rect 105322 390510 105952 390538
rect 105266 390487 105322 390496
rect 105174 389056 105230 389065
rect 105174 388991 105230 389000
rect 104806 385656 104862 385665
rect 104806 385591 104862 385600
rect 104544 383626 104756 383654
rect 104164 358760 104216 358766
rect 104164 358702 104216 358708
rect 104728 357406 104756 383626
rect 104716 357400 104768 357406
rect 104716 357342 104768 357348
rect 104164 320884 104216 320890
rect 104164 320826 104216 320832
rect 104176 294098 104204 320826
rect 104164 294092 104216 294098
rect 104164 294034 104216 294040
rect 104162 291272 104218 291281
rect 104162 291207 104218 291216
rect 103612 249076 103664 249082
rect 103612 249018 103664 249024
rect 103624 244934 103652 249018
rect 103612 244928 103664 244934
rect 103612 244870 103664 244876
rect 104176 236065 104204 291207
rect 104256 269136 104308 269142
rect 104256 269078 104308 269084
rect 104268 251054 104296 269078
rect 104820 267034 104848 385591
rect 105924 383625 105952 390510
rect 106338 390130 106366 390388
rect 106292 390102 106366 390130
rect 106476 390374 107088 390402
rect 106094 389056 106150 389065
rect 106094 388991 106150 389000
rect 105910 383616 105966 383625
rect 105910 383551 105966 383560
rect 106002 382936 106058 382945
rect 106002 382871 106058 382880
rect 105544 376032 105596 376038
rect 105544 375974 105596 375980
rect 104898 290048 104954 290057
rect 104898 289983 104954 289992
rect 104808 267028 104860 267034
rect 104808 266970 104860 266976
rect 104820 266422 104848 266970
rect 104808 266416 104860 266422
rect 104808 266358 104860 266364
rect 104256 251048 104308 251054
rect 104256 250990 104308 250996
rect 104808 248600 104860 248606
rect 104808 248542 104860 248548
rect 104254 241904 104310 241913
rect 104254 241839 104310 241848
rect 104162 236056 104218 236065
rect 104162 235991 104218 236000
rect 103518 235920 103574 235929
rect 103518 235855 103574 235864
rect 103428 218816 103480 218822
rect 103428 218758 103480 218764
rect 102324 211132 102376 211138
rect 102324 211074 102376 211080
rect 102336 209846 102364 211074
rect 102324 209840 102376 209846
rect 102324 209782 102376 209788
rect 102232 209772 102284 209778
rect 102232 209714 102284 209720
rect 102244 208418 102272 209714
rect 102232 208412 102284 208418
rect 102232 208354 102284 208360
rect 102048 103556 102100 103562
rect 102048 103498 102100 103504
rect 102060 103426 102088 103498
rect 102048 103420 102100 103426
rect 102048 103362 102100 103368
rect 101496 101448 101548 101454
rect 101496 101390 101548 101396
rect 101404 88324 101456 88330
rect 101404 88266 101456 88272
rect 100114 88088 100170 88097
rect 100114 88023 100170 88032
rect 100022 86728 100078 86737
rect 100022 86663 100078 86672
rect 101508 85474 101536 101390
rect 101588 98116 101640 98122
rect 101588 98058 101640 98064
rect 101496 85468 101548 85474
rect 101496 85410 101548 85416
rect 101600 84182 101628 98058
rect 102336 93702 102364 209782
rect 102782 149288 102838 149297
rect 102782 149223 102838 149232
rect 102796 130626 102824 149223
rect 102784 130620 102836 130626
rect 102784 130562 102836 130568
rect 102784 129056 102836 129062
rect 102784 128998 102836 129004
rect 102796 121106 102824 128998
rect 102784 121100 102836 121106
rect 102784 121042 102836 121048
rect 102324 93696 102376 93702
rect 102324 93638 102376 93644
rect 101588 84176 101640 84182
rect 101588 84118 101640 84124
rect 98734 82648 98790 82657
rect 98734 82583 98790 82592
rect 97448 78668 97500 78674
rect 97448 78610 97500 78616
rect 97356 78600 97408 78606
rect 97356 78542 97408 78548
rect 94504 67516 94556 67522
rect 94504 67458 94556 67464
rect 97368 64874 97396 78542
rect 101402 78024 101458 78033
rect 101402 77959 101458 77968
rect 98642 69592 98698 69601
rect 98642 69527 98698 69536
rect 93768 64864 93820 64870
rect 93768 64806 93820 64812
rect 97276 64846 97396 64874
rect 95146 54496 95202 54505
rect 95146 54431 95202 54440
rect 93124 20664 93176 20670
rect 93124 20606 93176 20612
rect 93768 19984 93820 19990
rect 93768 19926 93820 19932
rect 93780 3534 93808 19926
rect 95056 18624 95108 18630
rect 95056 18566 95108 18572
rect 95068 3534 95096 18566
rect 89168 3528 89220 3534
rect 89168 3470 89220 3476
rect 89628 3528 89680 3534
rect 89628 3470 89680 3476
rect 90364 3528 90416 3534
rect 90364 3470 90416 3476
rect 90916 3528 90968 3534
rect 90916 3470 90968 3476
rect 91008 3528 91060 3534
rect 91008 3470 91060 3476
rect 91560 3528 91612 3534
rect 91560 3470 91612 3476
rect 92756 3528 92808 3534
rect 92756 3470 92808 3476
rect 93768 3528 93820 3534
rect 93768 3470 93820 3476
rect 93952 3528 94004 3534
rect 93952 3470 94004 3476
rect 95056 3528 95108 3534
rect 95056 3470 95108 3476
rect 89180 480 89208 3470
rect 90376 480 90404 3470
rect 91572 480 91600 3470
rect 92768 480 92796 3470
rect 93964 480 93992 3470
rect 95160 480 95188 54431
rect 96252 4888 96304 4894
rect 96252 4830 96304 4836
rect 96264 480 96292 4830
rect 97276 4826 97304 64846
rect 97908 10396 97960 10402
rect 97908 10338 97960 10344
rect 97264 4820 97316 4826
rect 97264 4762 97316 4768
rect 97920 3534 97948 10338
rect 98656 6914 98684 69527
rect 101416 59362 101444 77959
rect 101404 59356 101456 59362
rect 101404 59298 101456 59304
rect 101404 51740 101456 51746
rect 101404 51682 101456 51688
rect 100668 25560 100720 25566
rect 100668 25502 100720 25508
rect 99288 17332 99340 17338
rect 99288 17274 99340 17280
rect 98564 6886 98684 6914
rect 97448 3528 97500 3534
rect 97448 3470 97500 3476
rect 97908 3528 97960 3534
rect 97908 3470 97960 3476
rect 97460 480 97488 3470
rect 98564 3466 98592 6886
rect 99300 3534 99328 17274
rect 100300 7608 100352 7614
rect 100300 7550 100352 7556
rect 98644 3528 98696 3534
rect 98644 3470 98696 3476
rect 99288 3528 99340 3534
rect 99288 3470 99340 3476
rect 99840 3528 99892 3534
rect 99840 3470 99892 3476
rect 98552 3460 98604 3466
rect 98552 3402 98604 3408
rect 98656 480 98684 3470
rect 99852 480 99880 3470
rect 100312 3369 100340 7550
rect 100680 3534 100708 25502
rect 101416 10334 101444 51682
rect 102048 22772 102100 22778
rect 102048 22714 102100 22720
rect 101404 10328 101456 10334
rect 101404 10270 101456 10276
rect 102060 3534 102088 22714
rect 103440 6914 103468 218758
rect 104268 218006 104296 241839
rect 104820 240145 104848 248542
rect 104806 240136 104862 240145
rect 104806 240071 104862 240080
rect 104714 236736 104770 236745
rect 104714 236671 104770 236680
rect 104624 236020 104676 236026
rect 104624 235962 104676 235968
rect 104256 218000 104308 218006
rect 104256 217942 104308 217948
rect 104164 187060 104216 187066
rect 104164 187002 104216 187008
rect 104176 90545 104204 187002
rect 104636 171154 104664 235962
rect 104624 171148 104676 171154
rect 104624 171090 104676 171096
rect 104636 161474 104664 171090
rect 104268 161446 104664 161474
rect 104268 141545 104296 161446
rect 104254 141536 104310 141545
rect 104254 141471 104310 141480
rect 104256 139460 104308 139466
rect 104256 139402 104308 139408
rect 104268 120766 104296 139402
rect 104256 120760 104308 120766
rect 104256 120702 104308 120708
rect 104728 93854 104756 236671
rect 104806 211848 104862 211857
rect 104806 211783 104862 211792
rect 104360 93826 104756 93854
rect 104162 90536 104218 90545
rect 104162 90471 104218 90480
rect 104176 82754 104204 90471
rect 104360 90409 104388 93826
rect 104346 90400 104402 90409
rect 104346 90335 104402 90344
rect 104164 82748 104216 82754
rect 104164 82690 104216 82696
rect 104360 80073 104388 90335
rect 104346 80064 104402 80073
rect 104346 79999 104402 80008
rect 104820 6914 104848 211783
rect 104912 143449 104940 289983
rect 104990 267880 105046 267889
rect 104990 267815 105046 267824
rect 105004 236026 105032 267815
rect 105556 254998 105584 375974
rect 105636 299464 105688 299470
rect 105636 299406 105688 299412
rect 105648 271862 105676 299406
rect 106016 287054 106044 382871
rect 106108 372570 106136 388991
rect 106096 372564 106148 372570
rect 106096 372506 106148 372512
rect 106016 287026 106136 287054
rect 105636 271856 105688 271862
rect 105636 271798 105688 271804
rect 106108 270609 106136 287026
rect 106188 271176 106240 271182
rect 106188 271118 106240 271124
rect 106094 270600 106150 270609
rect 106094 270535 106150 270544
rect 106108 270502 106136 270535
rect 106096 270496 106148 270502
rect 106096 270438 106148 270444
rect 106200 262206 106228 271118
rect 106188 262200 106240 262206
rect 106188 262142 106240 262148
rect 105544 254992 105596 254998
rect 105544 254934 105596 254940
rect 105544 252612 105596 252618
rect 105544 252554 105596 252560
rect 104992 236020 105044 236026
rect 104992 235962 105044 235968
rect 105556 221649 105584 252554
rect 106292 248606 106320 390102
rect 106372 382968 106424 382974
rect 106372 382910 106424 382916
rect 106280 248600 106332 248606
rect 106280 248542 106332 248548
rect 106384 236745 106412 382910
rect 106476 380769 106504 390374
rect 107948 389065 107976 390646
rect 111982 390623 112038 390632
rect 111996 390538 112024 390623
rect 111872 390524 112024 390538
rect 111858 390510 112024 390524
rect 108376 390374 108712 390402
rect 107934 389056 107990 389065
rect 107934 388991 107990 389000
rect 108684 387705 108712 390374
rect 109098 390130 109126 390388
rect 109512 390374 109848 390402
rect 109098 390102 109172 390130
rect 108854 389056 108910 389065
rect 108854 388991 108910 389000
rect 108670 387696 108726 387705
rect 108670 387631 108726 387640
rect 106462 380760 106518 380769
rect 106462 380695 106518 380704
rect 108868 365702 108896 388991
rect 108948 387796 109000 387802
rect 108948 387738 109000 387744
rect 108856 365696 108908 365702
rect 108856 365638 108908 365644
rect 107568 322176 107620 322182
rect 107568 322118 107620 322124
rect 107580 299470 107608 322118
rect 108856 304020 108908 304026
rect 108856 303962 108908 303968
rect 107568 299464 107620 299470
rect 107568 299406 107620 299412
rect 106462 291816 106518 291825
rect 106462 291751 106518 291760
rect 106370 236736 106426 236745
rect 106370 236671 106426 236680
rect 105542 221640 105598 221649
rect 105542 221575 105598 221584
rect 105542 217288 105598 217297
rect 105542 217223 105598 217232
rect 104898 143440 104954 143449
rect 104898 143375 104954 143384
rect 105556 90681 105584 217223
rect 106280 195288 106332 195294
rect 106280 195230 106332 195236
rect 105636 149116 105688 149122
rect 105636 149058 105688 149064
rect 105648 110362 105676 149058
rect 105636 110356 105688 110362
rect 105636 110298 105688 110304
rect 106292 102134 106320 195230
rect 106476 177342 106504 291751
rect 108396 289876 108448 289882
rect 108396 289818 108448 289824
rect 108304 274712 108356 274718
rect 108304 274654 108356 274660
rect 106924 251864 106976 251870
rect 106924 251806 106976 251812
rect 106936 241369 106964 251806
rect 107844 251184 107896 251190
rect 107844 251126 107896 251132
rect 107856 248414 107884 251126
rect 107764 248386 107884 248414
rect 107764 245002 107792 248386
rect 108316 246362 108344 274654
rect 108408 262886 108436 289818
rect 108396 262880 108448 262886
rect 108396 262822 108448 262828
rect 108396 253224 108448 253230
rect 108396 253166 108448 253172
rect 108304 246356 108356 246362
rect 108304 246298 108356 246304
rect 107752 244996 107804 245002
rect 107752 244938 107804 244944
rect 107016 242956 107068 242962
rect 107016 242898 107068 242904
rect 106922 241360 106978 241369
rect 106922 241295 106978 241304
rect 106554 236056 106610 236065
rect 106554 235991 106610 236000
rect 106464 177336 106516 177342
rect 106464 177278 106516 177284
rect 106568 144129 106596 235991
rect 106922 231160 106978 231169
rect 106922 231095 106978 231104
rect 106554 144120 106610 144129
rect 106554 144055 106610 144064
rect 106280 102128 106332 102134
rect 106280 102070 106332 102076
rect 106292 101454 106320 102070
rect 106280 101448 106332 101454
rect 106280 101390 106332 101396
rect 105542 90672 105598 90681
rect 105542 90607 105598 90616
rect 105556 81297 105584 90607
rect 105542 81288 105598 81297
rect 105542 81223 105598 81232
rect 106936 6914 106964 231095
rect 107028 219201 107056 242898
rect 107658 235920 107714 235929
rect 107658 235855 107714 235864
rect 107014 219192 107070 219201
rect 107014 219127 107070 219136
rect 107014 161528 107070 161537
rect 107014 161463 107070 161472
rect 107028 135969 107056 161463
rect 107566 144120 107622 144129
rect 107566 144055 107622 144064
rect 107014 135960 107070 135969
rect 107014 135895 107070 135904
rect 107016 130484 107068 130490
rect 107016 130426 107068 130432
rect 107028 118590 107056 130426
rect 107016 118584 107068 118590
rect 107016 118526 107068 118532
rect 103348 6886 103468 6914
rect 104544 6886 104848 6914
rect 106844 6886 106964 6914
rect 100668 3528 100720 3534
rect 100668 3470 100720 3476
rect 101036 3528 101088 3534
rect 101036 3470 101088 3476
rect 102048 3528 102100 3534
rect 102048 3470 102100 3476
rect 102232 3528 102284 3534
rect 102232 3470 102284 3476
rect 100298 3360 100354 3369
rect 100298 3295 100354 3304
rect 101048 480 101076 3470
rect 102244 480 102272 3470
rect 103348 480 103376 6886
rect 104544 480 104572 6886
rect 106844 3534 106872 6886
rect 107580 3534 107608 144055
rect 107672 84182 107700 235855
rect 107764 98705 107792 244938
rect 108316 195974 108344 246298
rect 108408 230450 108436 253166
rect 108868 252550 108896 303962
rect 108960 273222 108988 387738
rect 109040 387048 109092 387054
rect 109040 386990 109092 386996
rect 109052 379409 109080 386990
rect 109144 380186 109172 390102
rect 109512 387054 109540 390374
rect 110386 390130 110414 390388
rect 110524 390374 111136 390402
rect 110386 390102 110460 390130
rect 110432 389201 110460 390102
rect 110418 389192 110474 389201
rect 110418 389127 110474 389136
rect 109500 387048 109552 387054
rect 109500 386990 109552 386996
rect 109132 380180 109184 380186
rect 109132 380122 109184 380128
rect 109038 379400 109094 379409
rect 109038 379335 109094 379344
rect 109682 379400 109738 379409
rect 109682 379335 109738 379344
rect 108948 273216 109000 273222
rect 108948 273158 109000 273164
rect 108960 272542 108988 273158
rect 108948 272536 109000 272542
rect 108948 272478 109000 272484
rect 108488 252544 108540 252550
rect 108488 252486 108540 252492
rect 108856 252544 108908 252550
rect 108856 252486 108908 252492
rect 108500 250510 108528 252486
rect 109696 251190 109724 379335
rect 110524 373994 110552 390374
rect 111858 390130 111886 390510
rect 111996 390374 112608 390402
rect 111858 390102 111932 390130
rect 111904 389162 111932 390102
rect 111892 389156 111944 389162
rect 111892 389098 111944 389104
rect 111996 383654 112024 390374
rect 110432 373966 110552 373994
rect 111812 383626 112024 383654
rect 110432 274718 110460 373966
rect 111062 320784 111118 320793
rect 111062 320719 111118 320728
rect 110420 274712 110472 274718
rect 110420 274654 110472 274660
rect 111076 268394 111104 320719
rect 111154 284472 111210 284481
rect 111154 284407 111210 284416
rect 111064 268388 111116 268394
rect 111064 268330 111116 268336
rect 109776 266416 109828 266422
rect 109776 266358 109828 266364
rect 109684 251184 109736 251190
rect 109684 251126 109736 251132
rect 108488 250504 108540 250510
rect 108488 250446 108540 250452
rect 108396 230444 108448 230450
rect 108396 230386 108448 230392
rect 108304 195968 108356 195974
rect 108304 195910 108356 195916
rect 109040 162172 109092 162178
rect 109040 162114 109092 162120
rect 108302 145616 108358 145625
rect 108302 145551 108358 145560
rect 108316 128489 108344 145551
rect 108302 128480 108358 128489
rect 108302 128415 108358 128424
rect 107750 98696 107806 98705
rect 107750 98631 107806 98640
rect 108302 98696 108358 98705
rect 108302 98631 108358 98640
rect 108316 91769 108344 98631
rect 108302 91760 108358 91769
rect 108302 91695 108358 91704
rect 107660 84176 107712 84182
rect 107660 84118 107712 84124
rect 109052 77246 109080 162114
rect 109788 161474 109816 266358
rect 110972 247716 111024 247722
rect 110972 247658 111024 247664
rect 110984 247110 111012 247658
rect 110420 247104 110472 247110
rect 110420 247046 110472 247052
rect 110972 247104 111024 247110
rect 110972 247046 111024 247052
rect 110326 226944 110382 226953
rect 110326 226879 110382 226888
rect 109696 161446 109816 161474
rect 109696 160313 109724 161446
rect 109682 160304 109738 160313
rect 109682 160239 109738 160248
rect 109696 120086 109724 160239
rect 109684 120080 109736 120086
rect 109684 120022 109736 120028
rect 109040 77240 109092 77246
rect 109040 77182 109092 77188
rect 108948 33788 109000 33794
rect 108948 33730 109000 33736
rect 108960 3534 108988 33730
rect 110340 3534 110368 226879
rect 110432 90982 110460 247046
rect 111076 236706 111104 268330
rect 111168 260137 111196 284407
rect 111154 260128 111210 260137
rect 111154 260063 111210 260072
rect 111156 257372 111208 257378
rect 111156 257314 111208 257320
rect 111064 236700 111116 236706
rect 111064 236642 111116 236648
rect 111168 234598 111196 257314
rect 111812 249762 111840 383626
rect 112732 381750 112760 401775
rect 111892 381744 111944 381750
rect 111892 381686 111944 381692
rect 112720 381744 112772 381750
rect 112720 381686 112772 381692
rect 111904 380934 111932 381686
rect 111892 380928 111944 380934
rect 111892 380870 111944 380876
rect 111904 369850 111932 380870
rect 111892 369844 111944 369850
rect 111892 369786 111944 369792
rect 111904 369170 111932 369786
rect 111892 369164 111944 369170
rect 111892 369106 111944 369112
rect 113284 316742 113312 416735
rect 113376 402393 113404 468454
rect 114652 439544 114704 439550
rect 114652 439486 114704 439492
rect 114664 429321 114692 439486
rect 115020 434716 115072 434722
rect 115020 434658 115072 434664
rect 115032 433401 115060 434658
rect 115018 433392 115074 433401
rect 115018 433327 115074 433336
rect 115216 431954 115244 583714
rect 115296 569968 115348 569974
rect 115296 569910 115348 569916
rect 115308 458561 115336 569910
rect 115940 550656 115992 550662
rect 115940 550598 115992 550604
rect 115294 458552 115350 458561
rect 115294 458487 115350 458496
rect 115032 431926 115244 431954
rect 114650 429312 114706 429321
rect 114650 429247 114706 429256
rect 113454 426048 113510 426057
rect 113454 425983 113510 425992
rect 113362 402384 113418 402393
rect 113362 402319 113418 402328
rect 113468 384305 113496 425983
rect 114652 423768 114704 423774
rect 114652 423710 114704 423716
rect 114664 421977 114692 423710
rect 114650 421968 114706 421977
rect 114650 421903 114706 421912
rect 114558 420880 114614 420889
rect 114558 420815 114614 420824
rect 114572 402974 114600 420815
rect 115032 414089 115060 431926
rect 115308 431610 115336 458487
rect 115388 434036 115440 434042
rect 115388 433978 115440 433984
rect 115124 431582 115336 431610
rect 115124 424153 115152 431582
rect 115296 431316 115348 431322
rect 115296 431258 115348 431264
rect 115308 431225 115336 431258
rect 115294 431216 115350 431225
rect 115294 431151 115350 431160
rect 115296 426148 115348 426154
rect 115296 426090 115348 426096
rect 115308 426057 115336 426090
rect 115294 426048 115350 426057
rect 115294 425983 115350 425992
rect 115296 424992 115348 424998
rect 115294 424960 115296 424969
rect 115348 424960 115350 424969
rect 115294 424895 115350 424904
rect 115110 424144 115166 424153
rect 115110 424079 115166 424088
rect 115202 418976 115258 418985
rect 115202 418911 115258 418920
rect 115216 418130 115244 418911
rect 115204 418124 115256 418130
rect 115204 418066 115256 418072
rect 115018 414080 115074 414089
rect 115018 414015 115074 414024
rect 115032 412729 115060 414015
rect 115018 412720 115074 412729
rect 115018 412655 115074 412664
rect 115216 412634 115244 418066
rect 115216 412606 115336 412634
rect 115202 406464 115258 406473
rect 115202 406399 115258 406408
rect 114572 402946 114692 402974
rect 113824 397520 113876 397526
rect 113824 397462 113876 397468
rect 113836 387433 113864 397462
rect 114664 387802 114692 402946
rect 114744 401396 114796 401402
rect 114744 401338 114796 401344
rect 114756 400489 114784 401338
rect 114742 400480 114798 400489
rect 114742 400415 114798 400424
rect 114834 391232 114890 391241
rect 114834 391167 114890 391176
rect 114848 390794 114876 391167
rect 114836 390788 114888 390794
rect 114836 390730 114888 390736
rect 114652 387796 114704 387802
rect 114652 387738 114704 387744
rect 113822 387424 113878 387433
rect 113822 387359 113878 387368
rect 113454 384296 113510 384305
rect 113454 384231 113510 384240
rect 115216 349110 115244 406399
rect 115204 349104 115256 349110
rect 115204 349046 115256 349052
rect 113272 316736 113324 316742
rect 113272 316678 113324 316684
rect 113822 298208 113878 298217
rect 113822 298143 113878 298152
rect 112444 285796 112496 285802
rect 112444 285738 112496 285744
rect 111800 249756 111852 249762
rect 111800 249698 111852 249704
rect 111892 238740 111944 238746
rect 111892 238682 111944 238688
rect 111156 234592 111208 234598
rect 111156 234534 111208 234540
rect 111064 229764 111116 229770
rect 111064 229706 111116 229712
rect 110512 207732 110564 207738
rect 110512 207674 110564 207680
rect 110524 207058 110552 207674
rect 110512 207052 110564 207058
rect 110512 206994 110564 207000
rect 110524 106962 110552 206994
rect 110972 123480 111024 123486
rect 110972 123422 111024 123428
rect 110984 121446 111012 123422
rect 110972 121440 111024 121446
rect 110972 121382 111024 121388
rect 110512 106956 110564 106962
rect 110512 106898 110564 106904
rect 110420 90976 110472 90982
rect 110420 90918 110472 90924
rect 110432 89758 110460 90918
rect 110420 89752 110472 89758
rect 110420 89694 110472 89700
rect 111076 89690 111104 229706
rect 111800 228404 111852 228410
rect 111800 228346 111852 228352
rect 111812 89758 111840 228346
rect 111904 108361 111932 238682
rect 112456 229090 112484 285738
rect 113836 285569 113864 298143
rect 113822 285560 113878 285569
rect 113822 285495 113878 285504
rect 113822 281616 113878 281625
rect 113822 281551 113878 281560
rect 112536 249824 112588 249830
rect 112536 249766 112588 249772
rect 112548 238746 112576 249766
rect 112536 238740 112588 238746
rect 112536 238682 112588 238688
rect 112444 229084 112496 229090
rect 112444 229026 112496 229032
rect 113836 220794 113864 281551
rect 115216 271182 115244 349046
rect 115308 322182 115336 412606
rect 115400 405657 115428 433978
rect 115848 430296 115900 430302
rect 115848 430238 115900 430244
rect 115860 430137 115888 430238
rect 115846 430128 115902 430137
rect 115846 430063 115902 430072
rect 115848 428460 115900 428466
rect 115848 428402 115900 428408
rect 115860 428233 115888 428402
rect 115846 428224 115902 428233
rect 115846 428159 115902 428168
rect 115848 427780 115900 427786
rect 115848 427722 115900 427728
rect 115860 427145 115888 427722
rect 115846 427136 115902 427145
rect 115846 427071 115902 427080
rect 115848 423632 115900 423638
rect 115848 423574 115900 423580
rect 115860 423065 115888 423574
rect 115846 423056 115902 423065
rect 115846 422991 115902 423000
rect 115846 420064 115902 420073
rect 115846 419999 115902 420008
rect 115860 419558 115888 419999
rect 115848 419552 115900 419558
rect 115848 419494 115900 419500
rect 115848 418056 115900 418062
rect 115848 417998 115900 418004
rect 115860 416809 115888 417998
rect 115846 416800 115902 416809
rect 115846 416735 115902 416744
rect 115846 415712 115902 415721
rect 115846 415647 115902 415656
rect 115860 415478 115888 415647
rect 115848 415472 115900 415478
rect 115848 415414 115900 415420
rect 115848 413840 115900 413846
rect 115846 413808 115848 413817
rect 115900 413808 115902 413817
rect 115846 413743 115902 413752
rect 115846 410544 115902 410553
rect 115846 410479 115902 410488
rect 115860 409902 115888 410479
rect 115848 409896 115900 409902
rect 115848 409838 115900 409844
rect 115846 409728 115902 409737
rect 115846 409663 115902 409672
rect 115860 409154 115888 409663
rect 115848 409148 115900 409154
rect 115848 409090 115900 409096
rect 115846 408640 115902 408649
rect 115846 408575 115902 408584
rect 115860 408542 115888 408575
rect 115848 408536 115900 408542
rect 115848 408478 115900 408484
rect 115846 407552 115902 407561
rect 115846 407487 115902 407496
rect 115860 407182 115888 407487
rect 115848 407176 115900 407182
rect 115848 407118 115900 407124
rect 115756 405748 115808 405754
rect 115756 405690 115808 405696
rect 115768 405657 115796 405690
rect 115848 405680 115900 405686
rect 115386 405648 115442 405657
rect 115386 405583 115442 405592
rect 115754 405648 115810 405657
rect 115848 405622 115900 405628
rect 115754 405583 115810 405592
rect 115860 404569 115888 405622
rect 115846 404560 115902 404569
rect 115846 404495 115902 404504
rect 115846 403472 115902 403481
rect 115846 403407 115902 403416
rect 115860 403034 115888 403407
rect 115848 403028 115900 403034
rect 115848 402970 115900 402976
rect 115662 401296 115718 401305
rect 115662 401231 115718 401240
rect 115676 400246 115704 401231
rect 115664 400240 115716 400246
rect 115664 400182 115716 400188
rect 115846 399392 115902 399401
rect 115846 399327 115902 399336
rect 115860 398886 115888 399327
rect 115848 398880 115900 398886
rect 115848 398822 115900 398828
rect 115570 398304 115626 398313
rect 115570 398239 115626 398248
rect 115584 397594 115612 398239
rect 115572 397588 115624 397594
rect 115572 397530 115624 397536
rect 115846 396400 115902 396409
rect 115846 396335 115848 396344
rect 115900 396335 115902 396344
rect 115848 396306 115900 396312
rect 115846 395312 115902 395321
rect 115846 395247 115902 395256
rect 115860 394738 115888 395247
rect 115848 394732 115900 394738
rect 115848 394674 115900 394680
rect 115846 394224 115902 394233
rect 115846 394159 115902 394168
rect 115860 393378 115888 394159
rect 115848 393372 115900 393378
rect 115848 393314 115900 393320
rect 115846 393136 115902 393145
rect 115846 393071 115902 393080
rect 115860 392630 115888 393071
rect 115848 392624 115900 392630
rect 115848 392566 115900 392572
rect 115386 392048 115442 392057
rect 115386 391983 115442 391992
rect 115400 353258 115428 391983
rect 115952 382974 115980 550598
rect 116032 435464 116084 435470
rect 116032 435406 116084 435412
rect 116044 423774 116072 435406
rect 116032 423768 116084 423774
rect 116032 423710 116084 423716
rect 116122 418296 116178 418305
rect 116122 418231 116178 418240
rect 116030 414896 116086 414905
rect 116030 414831 116086 414840
rect 115940 382968 115992 382974
rect 115940 382910 115992 382916
rect 115940 371884 115992 371890
rect 115940 371826 115992 371832
rect 115388 353252 115440 353258
rect 115388 353194 115440 353200
rect 115296 322176 115348 322182
rect 115296 322118 115348 322124
rect 115400 304026 115428 353194
rect 115388 304020 115440 304026
rect 115388 303962 115440 303968
rect 115296 302252 115348 302258
rect 115296 302194 115348 302200
rect 115204 271176 115256 271182
rect 115204 271118 115256 271124
rect 115204 264988 115256 264994
rect 115204 264930 115256 264936
rect 115216 224913 115244 264930
rect 115308 238105 115336 302194
rect 115848 284368 115900 284374
rect 115848 284310 115900 284316
rect 115860 282198 115888 284310
rect 115848 282192 115900 282198
rect 115848 282134 115900 282140
rect 115952 247722 115980 371826
rect 116044 321570 116072 414831
rect 116136 411641 116164 418231
rect 116122 411632 116178 411641
rect 116122 411567 116178 411576
rect 116596 397497 116624 585142
rect 119342 583808 119398 583817
rect 119342 583743 119398 583752
rect 117320 561740 117372 561746
rect 117320 561682 117372 561688
rect 116676 454096 116728 454102
rect 116676 454038 116728 454044
rect 116688 436762 116716 454038
rect 116766 451344 116822 451353
rect 116766 451279 116822 451288
rect 116780 437345 116808 451279
rect 116766 437336 116822 437345
rect 116766 437271 116822 437280
rect 116676 436756 116728 436762
rect 116676 436698 116728 436704
rect 117332 413846 117360 561682
rect 118700 472660 118752 472666
rect 118700 472602 118752 472608
rect 118712 472054 118740 472602
rect 118700 472048 118752 472054
rect 118700 471990 118752 471996
rect 117412 471300 117464 471306
rect 117412 471242 117464 471248
rect 117424 470626 117452 471242
rect 117412 470620 117464 470626
rect 117412 470562 117464 470568
rect 117424 424998 117452 470562
rect 118712 431322 118740 471990
rect 119356 459610 119384 583743
rect 120080 573368 120132 573374
rect 120080 573310 120132 573316
rect 119344 459604 119396 459610
rect 119344 459546 119396 459552
rect 118700 431316 118752 431322
rect 118700 431258 118752 431264
rect 119356 426154 119384 459546
rect 119434 455560 119490 455569
rect 119434 455495 119490 455504
rect 119448 430302 119476 455495
rect 119436 430296 119488 430302
rect 119436 430238 119488 430244
rect 119344 426148 119396 426154
rect 119344 426090 119396 426096
rect 117412 424992 117464 424998
rect 117412 424934 117464 424940
rect 118700 416084 118752 416090
rect 118700 416026 118752 416032
rect 118712 415478 118740 416026
rect 118700 415472 118752 415478
rect 118700 415414 118752 415420
rect 117320 413840 117372 413846
rect 117320 413782 117372 413788
rect 116674 406328 116730 406337
rect 116674 406263 116730 406272
rect 116688 401402 116716 406263
rect 116676 401396 116728 401402
rect 116676 401338 116728 401344
rect 116582 397488 116638 397497
rect 116582 397423 116638 397432
rect 116584 390788 116636 390794
rect 116584 390730 116636 390736
rect 116596 364342 116624 390730
rect 117332 385665 117360 413782
rect 117964 397588 118016 397594
rect 117964 397530 118016 397536
rect 117318 385656 117374 385665
rect 117318 385591 117374 385600
rect 117976 376582 118004 397530
rect 118712 386345 118740 415414
rect 118792 400920 118844 400926
rect 118792 400862 118844 400868
rect 118804 397594 118832 400862
rect 118792 397588 118844 397594
rect 118792 397530 118844 397536
rect 119342 397488 119398 397497
rect 119342 397423 119398 397432
rect 118792 387796 118844 387802
rect 118792 387738 118844 387744
rect 118698 386336 118754 386345
rect 118698 386271 118754 386280
rect 118804 385014 118832 387738
rect 118792 385008 118844 385014
rect 118792 384950 118844 384956
rect 118700 377460 118752 377466
rect 118700 377402 118752 377408
rect 117964 376576 118016 376582
rect 117964 376518 118016 376524
rect 117976 376038 118004 376518
rect 117964 376032 118016 376038
rect 117964 375974 118016 375980
rect 117226 371920 117282 371929
rect 117226 371855 117228 371864
rect 117280 371855 117282 371864
rect 117228 371826 117280 371832
rect 116584 364336 116636 364342
rect 116584 364278 116636 364284
rect 116584 322244 116636 322250
rect 116584 322186 116636 322192
rect 116032 321564 116084 321570
rect 116032 321506 116084 321512
rect 116044 320793 116072 321506
rect 116030 320784 116086 320793
rect 116030 320719 116086 320728
rect 116596 307086 116624 322186
rect 116584 307080 116636 307086
rect 116584 307022 116636 307028
rect 117228 306400 117280 306406
rect 117228 306342 117280 306348
rect 116676 248464 116728 248470
rect 116676 248406 116728 248412
rect 115940 247716 115992 247722
rect 115940 247658 115992 247664
rect 115294 238096 115350 238105
rect 115294 238031 115350 238040
rect 115202 224904 115258 224913
rect 115202 224839 115258 224848
rect 115202 222864 115258 222873
rect 115202 222799 115258 222808
rect 113824 220788 113876 220794
rect 113824 220730 113876 220736
rect 114466 217288 114522 217297
rect 114466 217223 114522 217232
rect 113822 213208 113878 213217
rect 113822 213143 113878 213152
rect 113086 208992 113142 209001
rect 113086 208927 113142 208936
rect 111890 108352 111946 108361
rect 111890 108287 111946 108296
rect 111156 89752 111208 89758
rect 111156 89694 111208 89700
rect 111248 89752 111300 89758
rect 111248 89694 111300 89700
rect 111800 89752 111852 89758
rect 111800 89694 111852 89700
rect 111064 89684 111116 89690
rect 111064 89626 111116 89632
rect 111168 79801 111196 89694
rect 111260 81326 111288 89694
rect 111248 81320 111300 81326
rect 111248 81262 111300 81268
rect 111154 79792 111210 79801
rect 111154 79727 111210 79736
rect 111260 64874 111288 81262
rect 111076 64846 111288 64874
rect 111076 57866 111104 64846
rect 111064 57860 111116 57866
rect 111064 57802 111116 57808
rect 111708 36576 111760 36582
rect 111708 36518 111760 36524
rect 111720 6914 111748 36518
rect 113100 6914 113128 208927
rect 113836 89729 113864 213143
rect 113822 89720 113878 89729
rect 113822 89655 113878 89664
rect 114374 89720 114430 89729
rect 114374 89655 114430 89664
rect 114388 89622 114416 89655
rect 114376 89616 114428 89622
rect 114376 89558 114428 89564
rect 111628 6886 111748 6914
rect 112824 6886 113128 6914
rect 106832 3528 106884 3534
rect 106832 3470 106884 3476
rect 106924 3528 106976 3534
rect 106924 3470 106976 3476
rect 107568 3528 107620 3534
rect 107568 3470 107620 3476
rect 108120 3528 108172 3534
rect 108120 3470 108172 3476
rect 108948 3528 109000 3534
rect 108948 3470 109000 3476
rect 109316 3528 109368 3534
rect 109316 3470 109368 3476
rect 110328 3528 110380 3534
rect 110328 3470 110380 3476
rect 110510 3496 110566 3505
rect 105728 3460 105780 3466
rect 105728 3402 105780 3408
rect 105740 480 105768 3402
rect 106936 480 106964 3470
rect 108132 480 108160 3470
rect 109328 480 109356 3470
rect 110510 3431 110566 3440
rect 110524 480 110552 3431
rect 111628 480 111656 6886
rect 112824 480 112852 6886
rect 114480 3534 114508 217223
rect 115216 6914 115244 222799
rect 115308 89729 115336 238031
rect 116584 235272 116636 235278
rect 116584 235214 116636 235220
rect 115388 192568 115440 192574
rect 115388 192510 115440 192516
rect 115400 109002 115428 192510
rect 115938 181384 115994 181393
rect 115938 181319 115994 181328
rect 115388 108996 115440 109002
rect 115388 108938 115440 108944
rect 115294 89720 115350 89729
rect 115294 89655 115350 89664
rect 115308 79966 115336 89655
rect 115400 86970 115428 108938
rect 115388 86964 115440 86970
rect 115388 86906 115440 86912
rect 115296 79960 115348 79966
rect 115296 79902 115348 79908
rect 115952 74526 115980 181319
rect 116596 86902 116624 235214
rect 116688 233170 116716 248406
rect 116676 233164 116728 233170
rect 116676 233106 116728 233112
rect 116584 86896 116636 86902
rect 116584 86838 116636 86844
rect 115940 74520 115992 74526
rect 115940 74462 115992 74468
rect 115848 46300 115900 46306
rect 115848 46242 115900 46248
rect 115124 6886 115244 6914
rect 114008 3528 114060 3534
rect 114008 3470 114060 3476
rect 114468 3528 114520 3534
rect 114468 3470 114520 3476
rect 114020 480 114048 3470
rect 115124 3466 115152 6886
rect 115860 3534 115888 46242
rect 117240 3534 117268 306342
rect 118056 288448 118108 288454
rect 118056 288390 118108 288396
rect 117962 283112 118018 283121
rect 117962 283047 118018 283056
rect 117976 197334 118004 283047
rect 118068 277370 118096 288390
rect 118056 277364 118108 277370
rect 118056 277306 118108 277312
rect 118712 229770 118740 377402
rect 118804 302258 118832 384950
rect 119356 382265 119384 397423
rect 120092 388362 120120 573310
rect 120170 440328 120226 440337
rect 120170 440263 120226 440272
rect 120000 388334 120120 388362
rect 120000 387569 120028 388334
rect 119986 387560 120042 387569
rect 119986 387495 120042 387504
rect 120000 384334 120028 387495
rect 119988 384328 120040 384334
rect 119988 384270 120040 384276
rect 119342 382256 119398 382265
rect 119342 382191 119398 382200
rect 118792 302252 118844 302258
rect 118792 302194 118844 302200
rect 119344 296744 119396 296750
rect 119344 296686 119396 296692
rect 118976 289196 119028 289202
rect 118976 289138 119028 289144
rect 118988 281518 119016 289138
rect 118976 281512 119028 281518
rect 118976 281454 119028 281460
rect 119356 252550 119384 296686
rect 120184 289105 120212 440263
rect 120724 388068 120776 388074
rect 120724 388010 120776 388016
rect 120736 383654 120764 388010
rect 121472 387870 121500 585210
rect 122840 576904 122892 576910
rect 122840 576846 122892 576852
rect 122852 527882 122880 576846
rect 122840 527876 122892 527882
rect 122840 527818 122892 527824
rect 121552 475380 121604 475386
rect 121552 475322 121604 475328
rect 121564 388074 121592 475322
rect 122104 451308 122156 451314
rect 122104 451250 122156 451256
rect 122116 437442 122144 451250
rect 122104 437436 122156 437442
rect 122104 437378 122156 437384
rect 122104 396364 122156 396370
rect 122104 396306 122156 396312
rect 121552 388068 121604 388074
rect 121552 388010 121604 388016
rect 121460 387864 121512 387870
rect 121460 387806 121512 387812
rect 120724 383648 120776 383654
rect 120724 383590 120776 383596
rect 120736 364993 120764 383590
rect 121460 373312 121512 373318
rect 121460 373254 121512 373260
rect 120722 364984 120778 364993
rect 120722 364919 120778 364928
rect 120722 294536 120778 294545
rect 120722 294471 120778 294480
rect 120170 289096 120226 289105
rect 120170 289031 120226 289040
rect 119436 265736 119488 265742
rect 119436 265678 119488 265684
rect 119344 252544 119396 252550
rect 119344 252486 119396 252492
rect 119342 234016 119398 234025
rect 119342 233951 119398 233960
rect 118700 229764 118752 229770
rect 118700 229706 118752 229712
rect 118608 216028 118660 216034
rect 118608 215970 118660 215976
rect 117964 197328 118016 197334
rect 117964 197270 118016 197276
rect 117320 180124 117372 180130
rect 117320 180066 117372 180072
rect 117332 94518 117360 180066
rect 117320 94512 117372 94518
rect 117320 94454 117372 94460
rect 118620 3534 118648 215970
rect 118700 178696 118752 178702
rect 118700 178638 118752 178644
rect 118712 111790 118740 178638
rect 118700 111784 118752 111790
rect 118700 111726 118752 111732
rect 118712 111178 118740 111726
rect 118700 111172 118752 111178
rect 118700 111114 118752 111120
rect 119356 88233 119384 233951
rect 119448 228410 119476 265678
rect 119436 228404 119488 228410
rect 119436 228346 119488 228352
rect 119986 225720 120042 225729
rect 119986 225655 120042 225664
rect 119342 88224 119398 88233
rect 119342 88159 119398 88168
rect 119896 39364 119948 39370
rect 119896 39306 119948 39312
rect 119908 16574 119936 39306
rect 119816 16546 119936 16574
rect 115204 3528 115256 3534
rect 115204 3470 115256 3476
rect 115848 3528 115900 3534
rect 115848 3470 115900 3476
rect 116400 3528 116452 3534
rect 116400 3470 116452 3476
rect 117228 3528 117280 3534
rect 117228 3470 117280 3476
rect 117596 3528 117648 3534
rect 117596 3470 117648 3476
rect 118608 3528 118660 3534
rect 118608 3470 118660 3476
rect 115112 3460 115164 3466
rect 115112 3402 115164 3408
rect 115216 480 115244 3470
rect 116412 480 116440 3470
rect 117608 480 117636 3470
rect 119816 3126 119844 16546
rect 120000 6914 120028 225655
rect 120080 209092 120132 209098
rect 120080 209034 120132 209040
rect 120092 91118 120120 209034
rect 120736 196654 120764 294471
rect 121472 223582 121500 373254
rect 122116 367033 122144 396306
rect 122852 392630 122880 527818
rect 124312 498840 124364 498846
rect 124312 498782 124364 498788
rect 123484 496120 123536 496126
rect 123484 496062 123536 496068
rect 123496 462913 123524 496062
rect 123482 462904 123538 462913
rect 123482 462839 123538 462848
rect 123496 428466 123524 462839
rect 122932 428460 122984 428466
rect 122932 428402 122984 428408
rect 123484 428460 123536 428466
rect 123484 428402 123536 428408
rect 122840 392624 122892 392630
rect 122840 392566 122892 392572
rect 122102 367024 122158 367033
rect 122102 366959 122158 366968
rect 122746 310720 122802 310729
rect 122746 310655 122802 310664
rect 121460 223576 121512 223582
rect 121460 223518 121512 223524
rect 120724 196648 120776 196654
rect 120724 196590 120776 196596
rect 120172 182844 120224 182850
rect 120172 182786 120224 182792
rect 120184 93158 120212 182786
rect 120172 93152 120224 93158
rect 120172 93094 120224 93100
rect 120080 91112 120132 91118
rect 120080 91054 120132 91060
rect 120092 88330 120120 91054
rect 120080 88324 120132 88330
rect 120080 88266 120132 88272
rect 121472 85542 121500 223518
rect 121552 213308 121604 213314
rect 121552 213250 121604 213256
rect 121564 212566 121592 213250
rect 121552 212560 121604 212566
rect 121552 212502 121604 212508
rect 121564 104145 121592 212502
rect 121550 104136 121606 104145
rect 121550 104071 121606 104080
rect 121460 85536 121512 85542
rect 121460 85478 121512 85484
rect 121368 28280 121420 28286
rect 121368 28222 121420 28228
rect 121380 6914 121408 28222
rect 119908 6886 120028 6914
rect 121104 6886 121408 6914
rect 118792 3120 118844 3126
rect 118792 3062 118844 3068
rect 119804 3120 119856 3126
rect 119804 3062 119856 3068
rect 118804 480 118832 3062
rect 119908 480 119936 6886
rect 121104 480 121132 6886
rect 122760 3534 122788 310655
rect 122944 304201 122972 428402
rect 123484 392624 123536 392630
rect 123484 392566 123536 392572
rect 123496 360874 123524 392566
rect 124220 382220 124272 382226
rect 124220 382162 124272 382168
rect 123484 360868 123536 360874
rect 123484 360810 123536 360816
rect 122930 304192 122986 304201
rect 122930 304127 122986 304136
rect 122838 301472 122894 301481
rect 122838 301407 122894 301416
rect 122852 143313 122880 301407
rect 123496 269142 123524 360810
rect 123484 269136 123536 269142
rect 123484 269078 123536 269084
rect 122838 143304 122894 143313
rect 122838 143239 122894 143248
rect 122852 142769 122880 143239
rect 122838 142760 122894 142769
rect 122838 142695 122894 142704
rect 123496 113174 123524 269078
rect 124128 256012 124180 256018
rect 124128 255954 124180 255960
rect 123496 113146 123616 113174
rect 123588 106350 123616 113146
rect 123576 106344 123628 106350
rect 123576 106286 123628 106292
rect 123588 105602 123616 106286
rect 123576 105596 123628 105602
rect 123576 105538 123628 105544
rect 124140 3534 124168 255954
rect 124232 235278 124260 382162
rect 124324 380769 124352 498782
rect 124310 380760 124366 380769
rect 124310 380695 124366 380704
rect 124416 379409 124444 589290
rect 128360 587920 128412 587926
rect 128360 587862 128412 587868
rect 125600 576156 125652 576162
rect 125600 576098 125652 576104
rect 124862 417480 124918 417489
rect 124862 417415 124918 417424
rect 124876 409154 124904 417415
rect 124864 409148 124916 409154
rect 124864 409090 124916 409096
rect 124876 400897 124904 409090
rect 124862 400888 124918 400897
rect 124862 400823 124918 400832
rect 125612 387734 125640 576098
rect 125784 501628 125836 501634
rect 125784 501570 125836 501576
rect 125692 483676 125744 483682
rect 125692 483618 125744 483624
rect 125600 387728 125652 387734
rect 125600 387670 125652 387676
rect 125508 382968 125560 382974
rect 125508 382910 125560 382916
rect 125520 382226 125548 382910
rect 125508 382220 125560 382226
rect 125508 382162 125560 382168
rect 124862 380760 124918 380769
rect 124862 380695 124918 380704
rect 124402 379400 124458 379409
rect 124402 379335 124458 379344
rect 124876 360194 124904 380695
rect 125704 379438 125732 483618
rect 125796 406337 125824 501570
rect 126980 465724 127032 465730
rect 126980 465666 127032 465672
rect 126888 408604 126940 408610
rect 126888 408546 126940 408552
rect 125782 406328 125838 406337
rect 125782 406263 125838 406272
rect 126900 405686 126928 408546
rect 126888 405680 126940 405686
rect 126888 405622 126940 405628
rect 126992 388226 127020 465666
rect 128372 400926 128400 587862
rect 133142 582720 133198 582729
rect 133142 582655 133198 582664
rect 129740 554804 129792 554810
rect 129740 554746 129792 554752
rect 128452 478168 128504 478174
rect 128452 478110 128504 478116
rect 128464 417489 128492 478110
rect 128450 417480 128506 417489
rect 128450 417415 128506 417424
rect 128360 400920 128412 400926
rect 128360 400862 128412 400868
rect 127624 396092 127676 396098
rect 127624 396034 127676 396040
rect 126900 388198 127020 388226
rect 126244 387728 126296 387734
rect 126244 387670 126296 387676
rect 126256 383654 126284 387670
rect 126900 386345 126928 388198
rect 126886 386336 126942 386345
rect 126886 386271 126942 386280
rect 126900 384946 126928 386271
rect 126888 384940 126940 384946
rect 126888 384882 126940 384888
rect 126256 383626 126376 383654
rect 125692 379432 125744 379438
rect 125692 379374 125744 379380
rect 126348 370569 126376 383626
rect 127636 380905 127664 396034
rect 129004 393440 129056 393446
rect 129004 393382 129056 393388
rect 127622 380896 127678 380905
rect 127622 380831 127678 380840
rect 126428 379432 126480 379438
rect 126428 379374 126480 379380
rect 126334 370560 126390 370569
rect 126334 370495 126390 370504
rect 124864 360188 124916 360194
rect 124864 360130 124916 360136
rect 126242 298752 126298 298761
rect 126242 298687 126298 298696
rect 124864 262268 124916 262274
rect 124864 262210 124916 262216
rect 124220 235272 124272 235278
rect 124220 235214 124272 235220
rect 124876 149734 124904 262210
rect 126256 262206 126284 298687
rect 126244 262200 126296 262206
rect 126244 262142 126296 262148
rect 126244 258120 126296 258126
rect 126244 258062 126296 258068
rect 125508 238128 125560 238134
rect 125508 238070 125560 238076
rect 124954 153232 125010 153241
rect 124954 153167 125010 153176
rect 124864 149728 124916 149734
rect 124864 149670 124916 149676
rect 124876 115938 124904 149670
rect 124968 122738 124996 153167
rect 124956 122732 125008 122738
rect 124956 122674 125008 122680
rect 124864 115932 124916 115938
rect 124864 115874 124916 115880
rect 125520 3534 125548 238070
rect 125600 35216 125652 35222
rect 125600 35158 125652 35164
rect 125612 16574 125640 35158
rect 126256 17270 126284 258062
rect 126348 234025 126376 370495
rect 126440 368490 126468 379374
rect 126428 368484 126480 368490
rect 126428 368426 126480 368432
rect 129016 368422 129044 393382
rect 129752 387870 129780 554746
rect 130384 541000 130436 541006
rect 130384 540942 130436 540948
rect 130396 414730 130424 540942
rect 133156 461009 133184 582655
rect 134524 578264 134576 578270
rect 134524 578206 134576 578212
rect 133142 461000 133198 461009
rect 133142 460935 133198 460944
rect 132498 434752 132554 434761
rect 132498 434687 132554 434696
rect 130384 414724 130436 414730
rect 130384 414666 130436 414672
rect 129096 387864 129148 387870
rect 129096 387806 129148 387812
rect 129740 387864 129792 387870
rect 129740 387806 129792 387812
rect 129108 384985 129136 387806
rect 129094 384976 129150 384985
rect 129094 384911 129150 384920
rect 129108 379438 129136 384911
rect 130396 379506 130424 414666
rect 130384 379500 130436 379506
rect 130384 379442 130436 379448
rect 129096 379432 129148 379438
rect 129096 379374 129148 379380
rect 129096 370524 129148 370530
rect 129096 370466 129148 370472
rect 129004 368416 129056 368422
rect 129004 368358 129056 368364
rect 129004 365016 129056 365022
rect 129004 364958 129056 364964
rect 129016 354074 129044 364958
rect 129108 356046 129136 370466
rect 129096 356040 129148 356046
rect 129096 355982 129148 355988
rect 129004 354068 129056 354074
rect 129004 354010 129056 354016
rect 130476 336796 130528 336802
rect 130476 336738 130528 336744
rect 129004 329112 129056 329118
rect 129004 329054 129056 329060
rect 126888 325712 126940 325718
rect 126888 325654 126940 325660
rect 126900 320074 126928 325654
rect 126888 320068 126940 320074
rect 126888 320010 126940 320016
rect 127624 320068 127676 320074
rect 127624 320010 127676 320016
rect 126428 236700 126480 236706
rect 126428 236642 126480 236648
rect 126334 234016 126390 234025
rect 126334 233951 126390 233960
rect 126440 151814 126468 236642
rect 126348 151786 126468 151814
rect 126348 147801 126376 151786
rect 127636 150482 127664 320010
rect 128360 295384 128412 295390
rect 128360 295326 128412 295332
rect 128372 293962 128400 295326
rect 128360 293956 128412 293962
rect 128360 293898 128412 293904
rect 129016 276729 129044 329054
rect 129094 320240 129150 320249
rect 129094 320175 129150 320184
rect 129108 294642 129136 320175
rect 130384 304360 130436 304366
rect 130384 304302 130436 304308
rect 129096 294636 129148 294642
rect 129096 294578 129148 294584
rect 129094 287736 129150 287745
rect 129094 287671 129150 287680
rect 129108 287201 129136 287671
rect 129094 287192 129150 287201
rect 129094 287127 129150 287136
rect 129002 276720 129058 276729
rect 129002 276655 129058 276664
rect 129004 177404 129056 177410
rect 129004 177346 129056 177352
rect 127624 150476 127676 150482
rect 127624 150418 127676 150424
rect 127636 149802 127664 150418
rect 127624 149796 127676 149802
rect 127624 149738 127676 149744
rect 126334 147792 126390 147801
rect 126334 147727 126390 147736
rect 127624 147756 127676 147762
rect 126348 123486 126376 147727
rect 127624 147698 127676 147704
rect 126336 123480 126388 123486
rect 126336 123422 126388 123428
rect 127636 115938 127664 147698
rect 127624 115932 127676 115938
rect 127624 115874 127676 115880
rect 126244 17264 126296 17270
rect 126244 17206 126296 17212
rect 125612 16546 125916 16574
rect 122288 3528 122340 3534
rect 122288 3470 122340 3476
rect 122748 3528 122800 3534
rect 122748 3470 122800 3476
rect 123484 3528 123536 3534
rect 123484 3470 123536 3476
rect 124128 3528 124180 3534
rect 124128 3470 124180 3476
rect 124680 3528 124732 3534
rect 124680 3470 124732 3476
rect 125508 3528 125560 3534
rect 125508 3470 125560 3476
rect 122300 480 122328 3470
rect 123496 480 123524 3470
rect 124692 480 124720 3470
rect 125888 480 125916 16546
rect 129016 490 129044 177346
rect 129108 163538 129136 287127
rect 129186 270600 129242 270609
rect 129186 270535 129242 270544
rect 129096 163532 129148 163538
rect 129096 163474 129148 163480
rect 129200 161498 129228 270535
rect 129740 244928 129792 244934
rect 129740 244870 129792 244876
rect 129188 161492 129240 161498
rect 129188 161434 129240 161440
rect 129200 142154 129228 161434
rect 129108 142126 129228 142154
rect 129108 122806 129136 142126
rect 129096 122800 129148 122806
rect 129096 122742 129148 122748
rect 129752 103494 129780 244870
rect 129740 103488 129792 103494
rect 129740 103430 129792 103436
rect 129752 102814 129780 103430
rect 129740 102808 129792 102814
rect 129740 102750 129792 102756
rect 130396 18630 130424 304302
rect 130488 278662 130516 336738
rect 131762 302424 131818 302433
rect 131762 302359 131818 302368
rect 130568 283620 130620 283626
rect 130568 283562 130620 283568
rect 130476 278656 130528 278662
rect 130476 278598 130528 278604
rect 130580 241670 130608 283562
rect 130568 241664 130620 241670
rect 130568 241606 130620 241612
rect 131776 60042 131804 302359
rect 131764 60036 131816 60042
rect 131764 59978 131816 59984
rect 130384 18624 130436 18630
rect 130384 18566 130436 18572
rect 132512 16574 132540 434687
rect 133156 418062 133184 460935
rect 133144 418056 133196 418062
rect 133144 417998 133196 418004
rect 133142 300928 133198 300937
rect 133142 300863 133198 300872
rect 133156 192506 133184 300863
rect 133236 278044 133288 278050
rect 133236 277986 133288 277992
rect 133248 269074 133276 277986
rect 133236 269068 133288 269074
rect 133236 269010 133288 269016
rect 133236 259548 133288 259554
rect 133236 259490 133288 259496
rect 133248 230450 133276 259490
rect 133236 230444 133288 230450
rect 133236 230386 133288 230392
rect 133144 192500 133196 192506
rect 133144 192442 133196 192448
rect 133144 181484 133196 181490
rect 133144 181426 133196 181432
rect 133156 32434 133184 181426
rect 133144 32428 133196 32434
rect 133144 32370 133196 32376
rect 132512 16546 133000 16574
rect 129200 598 129412 626
rect 129200 490 129228 598
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129016 462 129228 490
rect 129384 480 129412 598
rect 132972 480 133000 16546
rect 134536 4214 134564 578206
rect 136652 538218 136680 703582
rect 137664 703474 137692 703582
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 137848 703474 137876 703520
rect 137664 703446 137876 703474
rect 154132 702846 154160 703520
rect 154120 702840 154172 702846
rect 154120 702782 154172 702788
rect 170324 702574 170352 703520
rect 191748 703384 191800 703390
rect 191748 703326 191800 703332
rect 173808 702772 173860 702778
rect 173808 702714 173860 702720
rect 170312 702568 170364 702574
rect 170312 702510 170364 702516
rect 143540 587240 143592 587246
rect 143540 587182 143592 587188
rect 136640 538212 136692 538218
rect 136640 538154 136692 538160
rect 136638 536072 136694 536081
rect 136638 536007 136694 536016
rect 136652 389042 136680 536007
rect 141424 530596 141476 530602
rect 141424 530538 141476 530544
rect 137284 465112 137336 465118
rect 137284 465054 137336 465060
rect 137296 451382 137324 465054
rect 141436 463826 141464 530538
rect 142896 469260 142948 469266
rect 142896 469202 142948 469208
rect 141424 463820 141476 463826
rect 141424 463762 141476 463768
rect 137284 451376 137336 451382
rect 137284 451318 137336 451324
rect 136560 389014 136680 389042
rect 136560 387705 136588 389014
rect 136546 387696 136602 387705
rect 136546 387631 136602 387640
rect 137296 335374 137324 451318
rect 141436 434926 141464 463762
rect 142066 451888 142122 451897
rect 142066 451823 142122 451832
rect 142080 451314 142108 451823
rect 142068 451308 142120 451314
rect 142068 451250 142120 451256
rect 137376 434920 137428 434926
rect 137376 434862 137428 434868
rect 141424 434920 141476 434926
rect 141424 434862 141476 434868
rect 137388 423638 137416 434862
rect 137376 423632 137428 423638
rect 137376 423574 137428 423580
rect 137928 422952 137980 422958
rect 137928 422894 137980 422900
rect 137940 416090 137968 422894
rect 137928 416084 137980 416090
rect 137928 416026 137980 416032
rect 137284 335368 137336 335374
rect 137284 335310 137336 335316
rect 135902 328536 135958 328545
rect 135902 328471 135958 328480
rect 134614 291816 134670 291825
rect 134614 291751 134670 291760
rect 134628 51746 134656 291751
rect 134616 51740 134668 51746
rect 134616 51682 134668 51688
rect 135916 46238 135944 328471
rect 137296 320890 137324 335310
rect 138664 331288 138716 331294
rect 138664 331230 138716 331236
rect 137466 326360 137522 326369
rect 137466 326295 137522 326304
rect 137284 320884 137336 320890
rect 137284 320826 137336 320832
rect 135996 316736 136048 316742
rect 135996 316678 136048 316684
rect 136008 301510 136036 316678
rect 135996 301504 136048 301510
rect 135996 301446 136048 301452
rect 135996 272536 136048 272542
rect 135996 272478 136048 272484
rect 136008 241534 136036 272478
rect 137374 267200 137430 267209
rect 137374 267135 137430 267144
rect 137282 261488 137338 261497
rect 137282 261423 137338 261432
rect 135996 241528 136048 241534
rect 135996 241470 136048 241476
rect 135904 46232 135956 46238
rect 135904 46174 135956 46180
rect 137296 21418 137324 261423
rect 137388 43450 137416 267135
rect 137480 251161 137508 326295
rect 137466 251152 137522 251161
rect 137466 251087 137522 251096
rect 138676 53106 138704 331230
rect 142080 321638 142108 451250
rect 142804 329928 142856 329934
rect 142804 329870 142856 329876
rect 141516 321632 141568 321638
rect 141516 321574 141568 321580
rect 142068 321632 142120 321638
rect 142068 321574 142120 321580
rect 141424 305108 141476 305114
rect 141424 305050 141476 305056
rect 140136 294636 140188 294642
rect 140136 294578 140188 294584
rect 140042 268560 140098 268569
rect 140042 268495 140098 268504
rect 138756 145036 138808 145042
rect 138756 144978 138808 144984
rect 138768 132462 138796 144978
rect 138756 132456 138808 132462
rect 138756 132398 138808 132404
rect 138664 53100 138716 53106
rect 138664 53042 138716 53048
rect 140056 44878 140084 268495
rect 140148 243574 140176 294578
rect 140136 243568 140188 243574
rect 140136 243510 140188 243516
rect 140044 44872 140096 44878
rect 140044 44814 140096 44820
rect 137376 43444 137428 43450
rect 137376 43386 137428 43392
rect 141436 22778 141464 305050
rect 141528 287745 141556 321574
rect 141514 287736 141570 287745
rect 141514 287671 141570 287680
rect 141514 273864 141570 273873
rect 141514 273799 141570 273808
rect 141528 36582 141556 273799
rect 141608 167068 141660 167074
rect 141608 167010 141660 167016
rect 141620 135998 141648 167010
rect 141700 136672 141752 136678
rect 141700 136614 141752 136620
rect 141608 135992 141660 135998
rect 141608 135934 141660 135940
rect 141712 123486 141740 136614
rect 141700 123480 141752 123486
rect 141700 123422 141752 123428
rect 142816 40730 142844 329870
rect 142908 320142 142936 469202
rect 143552 408610 143580 587182
rect 148324 581052 148376 581058
rect 148324 580994 148376 581000
rect 148336 458250 148364 580994
rect 159364 469328 159416 469334
rect 159364 469270 159416 469276
rect 148324 458244 148376 458250
rect 148324 458186 148376 458192
rect 147586 454200 147642 454209
rect 147586 454135 147642 454144
rect 143540 408604 143592 408610
rect 143540 408546 143592 408552
rect 144184 408604 144236 408610
rect 144184 408546 144236 408552
rect 144196 380905 144224 408546
rect 144182 380896 144238 380905
rect 144182 380831 144238 380840
rect 146942 331256 146998 331265
rect 146942 331191 146998 331200
rect 144276 324964 144328 324970
rect 144276 324906 144328 324912
rect 142896 320136 142948 320142
rect 142896 320078 142948 320084
rect 143448 320136 143500 320142
rect 143448 320078 143500 320084
rect 143460 319462 143488 320078
rect 143448 319456 143500 319462
rect 143448 319398 143500 319404
rect 144182 316160 144238 316169
rect 144182 316095 144238 316104
rect 142896 305040 142948 305046
rect 142896 304982 142948 304988
rect 142908 46306 142936 304982
rect 142986 269784 143042 269793
rect 142986 269719 143042 269728
rect 143000 247722 143028 269719
rect 142988 247716 143040 247722
rect 142988 247658 143040 247664
rect 144196 185638 144224 316095
rect 144288 265742 144316 324906
rect 145562 317520 145618 317529
rect 145562 317455 145618 317464
rect 144828 269816 144880 269822
rect 144828 269758 144880 269764
rect 144276 265736 144328 265742
rect 144276 265678 144328 265684
rect 144184 185632 144236 185638
rect 144184 185574 144236 185580
rect 144182 156224 144238 156233
rect 144182 156159 144238 156168
rect 144196 125526 144224 156159
rect 144184 125520 144236 125526
rect 144184 125462 144236 125468
rect 142988 62824 143040 62830
rect 142988 62766 143040 62772
rect 142896 46300 142948 46306
rect 142896 46242 142948 46248
rect 142804 40724 142856 40730
rect 142804 40666 142856 40672
rect 141516 36576 141568 36582
rect 141516 36518 141568 36524
rect 141424 22772 141476 22778
rect 141424 22714 141476 22720
rect 137284 21412 137336 21418
rect 137284 21354 137336 21360
rect 134524 4208 134576 4214
rect 134524 4150 134576 4156
rect 136456 4208 136508 4214
rect 136456 4150 136508 4156
rect 136468 480 136496 4150
rect 143000 2786 143028 62766
rect 144840 3534 144868 269758
rect 145576 37942 145604 317455
rect 145656 269884 145708 269890
rect 145656 269826 145708 269832
rect 145668 253230 145696 269826
rect 145748 259480 145800 259486
rect 145748 259422 145800 259428
rect 145656 253224 145708 253230
rect 145656 253166 145708 253172
rect 145760 243574 145788 259422
rect 145748 243568 145800 243574
rect 145748 243510 145800 243516
rect 146956 47598 146984 331191
rect 147036 299532 147088 299538
rect 147036 299474 147088 299480
rect 147048 244934 147076 299474
rect 147128 245676 147180 245682
rect 147128 245618 147180 245624
rect 147036 244928 147088 244934
rect 147036 244870 147088 244876
rect 147140 202842 147168 245618
rect 147128 202836 147180 202842
rect 147128 202778 147180 202784
rect 147034 164384 147090 164393
rect 147034 164319 147090 164328
rect 147048 128314 147076 164319
rect 147128 134632 147180 134638
rect 147128 134574 147180 134580
rect 147036 128308 147088 128314
rect 147036 128250 147088 128256
rect 147140 125526 147168 134574
rect 147128 125520 147180 125526
rect 147128 125462 147180 125468
rect 146944 47592 146996 47598
rect 146944 47534 146996 47540
rect 145564 37936 145616 37942
rect 145564 37878 145616 37884
rect 147600 3534 147628 454135
rect 148336 422958 148364 458186
rect 157340 456884 157392 456890
rect 157340 456826 157392 456832
rect 151084 454164 151136 454170
rect 151084 454106 151136 454112
rect 151096 429146 151124 454106
rect 151084 429140 151136 429146
rect 151084 429082 151136 429088
rect 157248 424380 157300 424386
rect 157248 424322 157300 424328
rect 148324 422952 148376 422958
rect 148324 422894 148376 422900
rect 155224 409896 155276 409902
rect 155224 409838 155276 409844
rect 152464 400240 152516 400246
rect 152464 400182 152516 400188
rect 151084 398880 151136 398886
rect 151084 398822 151136 398828
rect 151096 369782 151124 398822
rect 151084 369776 151136 369782
rect 151084 369718 151136 369724
rect 152476 368422 152504 400182
rect 155236 376553 155264 409838
rect 155222 376544 155278 376553
rect 155222 376479 155278 376488
rect 152464 368416 152516 368422
rect 152464 368358 152516 368364
rect 152556 354068 152608 354074
rect 152556 354010 152608 354016
rect 151176 323060 151228 323066
rect 151176 323002 151228 323008
rect 151084 307828 151136 307834
rect 151084 307770 151136 307776
rect 148324 306468 148376 306474
rect 148324 306410 148376 306416
rect 148336 10402 148364 306410
rect 148414 301472 148470 301481
rect 148414 301407 148470 301416
rect 148428 188358 148456 301407
rect 149796 299532 149848 299538
rect 149796 299474 149848 299480
rect 149704 282192 149756 282198
rect 149704 282134 149756 282140
rect 148508 263696 148560 263702
rect 148508 263638 148560 263644
rect 148520 227118 148548 263638
rect 148508 227112 148560 227118
rect 148508 227054 148560 227060
rect 148416 188352 148468 188358
rect 148416 188294 148468 188300
rect 148416 161560 148468 161566
rect 148416 161502 148468 161508
rect 148428 132394 148456 161502
rect 149716 142866 149744 282134
rect 149808 193866 149836 299474
rect 149886 274816 149942 274825
rect 149886 274751 149942 274760
rect 149900 228410 149928 274751
rect 149888 228404 149940 228410
rect 149888 228346 149940 228352
rect 149796 193860 149848 193866
rect 149796 193802 149848 193808
rect 149794 153368 149850 153377
rect 149794 153303 149850 153312
rect 149704 142860 149756 142866
rect 149704 142802 149756 142808
rect 148416 132388 148468 132394
rect 148416 132330 148468 132336
rect 149808 117298 149836 153303
rect 149796 117292 149848 117298
rect 149796 117234 149848 117240
rect 151096 39370 151124 307770
rect 151188 289202 151216 323002
rect 152462 303920 152518 303929
rect 152462 303855 152518 303864
rect 151176 289196 151228 289202
rect 151176 289138 151228 289144
rect 151174 280800 151230 280809
rect 151174 280735 151230 280744
rect 151188 42090 151216 280735
rect 151268 265668 151320 265674
rect 151268 265610 151320 265616
rect 151280 241466 151308 265610
rect 151360 244996 151412 245002
rect 151360 244938 151412 244944
rect 151268 241460 151320 241466
rect 151268 241402 151320 241408
rect 151372 233238 151400 244938
rect 151360 233232 151412 233238
rect 151360 233174 151412 233180
rect 151266 157584 151322 157593
rect 151266 157519 151322 157528
rect 151280 135930 151308 157519
rect 151268 135924 151320 135930
rect 151268 135866 151320 135872
rect 151176 42084 151228 42090
rect 151176 42026 151228 42032
rect 151084 39364 151136 39370
rect 151084 39306 151136 39312
rect 152476 24138 152504 303855
rect 152568 287054 152596 354010
rect 155406 327176 155462 327185
rect 155406 327111 155462 327120
rect 153844 314764 153896 314770
rect 153844 314706 153896 314712
rect 153108 302932 153160 302938
rect 153108 302874 153160 302880
rect 152568 287026 152688 287054
rect 152660 284306 152688 287026
rect 152648 284300 152700 284306
rect 152648 284242 152700 284248
rect 152660 283626 152688 284242
rect 152648 283620 152700 283626
rect 152648 283562 152700 283568
rect 152554 271144 152610 271153
rect 152554 271079 152610 271088
rect 152568 222970 152596 271079
rect 152556 222964 152608 222970
rect 152556 222906 152608 222912
rect 152554 154728 152610 154737
rect 152554 154663 152610 154672
rect 152568 130490 152596 154663
rect 152646 135960 152702 135969
rect 152646 135895 152702 135904
rect 152556 130484 152608 130490
rect 152556 130426 152608 130432
rect 152660 126954 152688 135895
rect 152648 126948 152700 126954
rect 152648 126890 152700 126896
rect 152556 107704 152608 107710
rect 152556 107646 152608 107652
rect 152568 75818 152596 107646
rect 153120 94761 153148 302874
rect 153106 94752 153162 94761
rect 153106 94687 153162 94696
rect 152556 75812 152608 75818
rect 152556 75754 152608 75760
rect 152464 24132 152516 24138
rect 152464 24074 152516 24080
rect 153856 11762 153884 314706
rect 155224 309188 155276 309194
rect 155224 309130 155276 309136
rect 153936 253972 153988 253978
rect 153936 253914 153988 253920
rect 153948 234025 153976 253914
rect 153934 234016 153990 234025
rect 153934 233951 153990 233960
rect 154488 217320 154540 217326
rect 154488 217262 154540 217268
rect 154500 211138 154528 217262
rect 154488 211132 154540 211138
rect 154488 211074 154540 211080
rect 154028 175364 154080 175370
rect 154028 175306 154080 175312
rect 153936 173936 153988 173942
rect 153936 173878 153988 173884
rect 153948 164898 153976 173878
rect 154040 169046 154068 175306
rect 154028 169040 154080 169046
rect 154028 168982 154080 168988
rect 154488 169040 154540 169046
rect 154488 168982 154540 168988
rect 153936 164892 153988 164898
rect 153936 164834 153988 164840
rect 154500 163606 154528 168982
rect 154488 163600 154540 163606
rect 154488 163542 154540 163548
rect 153936 162920 153988 162926
rect 153936 162862 153988 162868
rect 153948 153950 153976 162862
rect 153936 153944 153988 153950
rect 153936 153886 153988 153892
rect 155236 33794 155264 309130
rect 155314 293176 155370 293185
rect 155314 293111 155370 293120
rect 155328 186998 155356 293111
rect 155420 258738 155448 327111
rect 156602 289096 156658 289105
rect 156602 289031 156658 289040
rect 155958 267064 156014 267073
rect 155958 266999 156014 267008
rect 156418 267064 156474 267073
rect 156418 266999 156420 267008
rect 155408 258732 155460 258738
rect 155408 258674 155460 258680
rect 155316 186992 155368 186998
rect 155316 186934 155368 186940
rect 155314 149424 155370 149433
rect 155314 149359 155370 149368
rect 155328 118658 155356 149359
rect 155972 144809 156000 266999
rect 156472 266999 156474 267008
rect 156420 266970 156472 266976
rect 156616 171834 156644 289031
rect 157260 287065 157288 424322
rect 157246 287056 157302 287065
rect 157246 286991 157302 287000
rect 157260 285841 157288 286991
rect 157246 285832 157302 285841
rect 157246 285767 157302 285776
rect 156696 280220 156748 280226
rect 156696 280162 156748 280168
rect 156708 233170 156736 280162
rect 157352 278730 157380 456826
rect 159376 427786 159404 469270
rect 166908 461032 166960 461038
rect 166908 460974 166960 460980
rect 166262 453112 166318 453121
rect 166262 453047 166318 453056
rect 166276 443698 166304 453047
rect 166264 443692 166316 443698
rect 166264 443634 166316 443640
rect 162124 441652 162176 441658
rect 162124 441594 162176 441600
rect 161388 440904 161440 440910
rect 161388 440846 161440 440852
rect 159364 427780 159416 427786
rect 159364 427722 159416 427728
rect 159456 416084 159508 416090
rect 159456 416026 159508 416032
rect 159364 403096 159416 403102
rect 159364 403038 159416 403044
rect 158718 376680 158774 376689
rect 159376 376650 159404 403038
rect 159468 376689 159496 416026
rect 159454 376680 159510 376689
rect 158718 376615 158774 376624
rect 159364 376644 159416 376650
rect 158732 322250 158760 376615
rect 159454 376615 159510 376624
rect 159364 376586 159416 376592
rect 159376 332625 159404 376586
rect 159362 332616 159418 332625
rect 159362 332551 159418 332560
rect 159376 323610 159404 332551
rect 159364 323604 159416 323610
rect 159364 323546 159416 323552
rect 158720 322244 158772 322250
rect 158720 322186 158772 322192
rect 159546 321600 159602 321609
rect 159546 321535 159602 321544
rect 159456 300892 159508 300898
rect 159456 300834 159508 300840
rect 157984 287768 158036 287774
rect 157984 287710 158036 287716
rect 157996 287162 158024 287710
rect 159364 287700 159416 287706
rect 159364 287642 159416 287648
rect 157984 287156 158036 287162
rect 157984 287098 158036 287104
rect 157340 278724 157392 278730
rect 157340 278666 157392 278672
rect 157352 272610 157380 278666
rect 157340 272604 157392 272610
rect 157340 272546 157392 272552
rect 156696 233164 156748 233170
rect 156696 233106 156748 233112
rect 156696 218748 156748 218754
rect 156696 218690 156748 218696
rect 156604 171828 156656 171834
rect 156604 171770 156656 171776
rect 156708 151201 156736 218690
rect 157996 166326 158024 287098
rect 159376 287094 159404 287642
rect 159364 287088 159416 287094
rect 159364 287030 159416 287036
rect 158626 269784 158682 269793
rect 158626 269719 158682 269728
rect 158074 235376 158130 235385
rect 158074 235311 158130 235320
rect 158088 204270 158116 235311
rect 158640 217938 158668 269719
rect 158628 217932 158680 217938
rect 158628 217874 158680 217880
rect 158076 204264 158128 204270
rect 158076 204206 158128 204212
rect 157984 166320 158036 166326
rect 157984 166262 158036 166268
rect 156694 151192 156750 151201
rect 156694 151127 156750 151136
rect 155958 144800 156014 144809
rect 155958 144735 156014 144744
rect 156694 144800 156750 144809
rect 156694 144735 156750 144744
rect 156604 143608 156656 143614
rect 156708 143585 156736 144735
rect 156604 143550 156656 143556
rect 156694 143576 156750 143585
rect 156616 129062 156644 143550
rect 156694 143511 156750 143520
rect 156708 131102 156736 143511
rect 158088 142154 158116 204206
rect 157996 142126 158116 142154
rect 157996 138689 158024 142126
rect 157982 138680 158038 138689
rect 157982 138615 158038 138624
rect 156696 131096 156748 131102
rect 156696 131038 156748 131044
rect 156604 129056 156656 129062
rect 156604 128998 156656 129004
rect 155316 118652 155368 118658
rect 155316 118594 155368 118600
rect 157996 113150 158024 138615
rect 157984 113144 158036 113150
rect 157984 113086 158036 113092
rect 158640 108934 158668 217874
rect 159376 141506 159404 287030
rect 159468 256018 159496 300834
rect 159560 280158 159588 321535
rect 160926 285832 160982 285841
rect 160926 285767 160928 285776
rect 160980 285767 160982 285776
rect 160928 285738 160980 285744
rect 159548 280152 159600 280158
rect 159548 280094 159600 280100
rect 159546 268424 159602 268433
rect 159546 268359 159602 268368
rect 159456 256012 159508 256018
rect 159456 255954 159508 255960
rect 159560 234598 159588 268359
rect 160744 253972 160796 253978
rect 160744 253914 160796 253920
rect 160008 251184 160060 251190
rect 160008 251126 160060 251132
rect 160020 249830 160048 251126
rect 160008 249824 160060 249830
rect 160008 249766 160060 249772
rect 160020 235278 160048 249766
rect 160008 235272 160060 235278
rect 160008 235214 160060 235220
rect 159548 234592 159600 234598
rect 159548 234534 159600 234540
rect 159456 222896 159508 222902
rect 159456 222838 159508 222844
rect 159468 217977 159496 222838
rect 159454 217968 159510 217977
rect 159454 217903 159510 217912
rect 159468 147694 159496 217903
rect 159560 178090 159588 234534
rect 159548 178084 159600 178090
rect 159548 178026 159600 178032
rect 159456 147688 159508 147694
rect 159456 147630 159508 147636
rect 159364 141500 159416 141506
rect 159364 141442 159416 141448
rect 159364 135924 159416 135930
rect 159364 135866 159416 135872
rect 155316 108928 155368 108934
rect 155316 108870 155368 108876
rect 158628 108928 158680 108934
rect 158628 108870 158680 108876
rect 155328 93129 155356 108870
rect 157984 106412 158036 106418
rect 157984 106354 158036 106360
rect 155314 93120 155370 93129
rect 155314 93055 155370 93064
rect 155498 93120 155554 93129
rect 155498 93055 155554 93064
rect 155512 82822 155540 93055
rect 155500 82816 155552 82822
rect 155500 82758 155552 82764
rect 157996 82657 158024 106354
rect 157982 82648 158038 82657
rect 157982 82583 158038 82592
rect 155224 33788 155276 33794
rect 155224 33730 155276 33736
rect 153844 11756 153896 11762
rect 153844 11698 153896 11704
rect 148324 10396 148376 10402
rect 148324 10338 148376 10344
rect 159376 7614 159404 135866
rect 159468 117298 159496 147630
rect 159560 145761 159588 178026
rect 159546 145752 159602 145761
rect 159546 145687 159602 145696
rect 159456 117292 159508 117298
rect 159456 117234 159508 117240
rect 160756 26926 160784 253914
rect 160836 249824 160888 249830
rect 160836 249766 160888 249772
rect 160848 31074 160876 249766
rect 160940 173194 160968 285738
rect 161400 282849 161428 440846
rect 162136 412078 162164 441594
rect 162124 412072 162176 412078
rect 162124 412014 162176 412020
rect 162768 412072 162820 412078
rect 162768 412014 162820 412020
rect 162780 411942 162808 412014
rect 162768 411936 162820 411942
rect 162768 411878 162820 411884
rect 162124 405816 162176 405822
rect 162124 405758 162176 405764
rect 162136 378146 162164 405758
rect 162124 378140 162176 378146
rect 162124 378082 162176 378088
rect 162136 322998 162164 378082
rect 161940 322992 161992 322998
rect 161940 322934 161992 322940
rect 162124 322992 162176 322998
rect 162124 322934 162176 322940
rect 161952 322153 161980 322934
rect 161938 322144 161994 322153
rect 161938 322079 161994 322088
rect 162780 313449 162808 411878
rect 166262 406328 166318 406337
rect 166262 406263 166318 406272
rect 163596 390584 163648 390590
rect 163596 390526 163648 390532
rect 163504 380180 163556 380186
rect 163504 380122 163556 380128
rect 163516 372502 163544 380122
rect 163504 372496 163556 372502
rect 163504 372438 163556 372444
rect 163502 318880 163558 318889
rect 163502 318815 163558 318824
rect 162122 313440 162178 313449
rect 162122 313375 162178 313384
rect 162766 313440 162822 313449
rect 162766 313375 162822 313384
rect 161386 282840 161442 282849
rect 161386 282775 161442 282784
rect 161110 272504 161166 272513
rect 161110 272439 161166 272448
rect 161020 253224 161072 253230
rect 161020 253166 161072 253172
rect 160928 173188 160980 173194
rect 160928 173130 160980 173136
rect 161032 146946 161060 253166
rect 161124 251190 161152 272439
rect 162136 269890 162164 313375
rect 162306 282840 162362 282849
rect 162306 282775 162362 282784
rect 162320 281625 162348 282775
rect 162306 281616 162362 281625
rect 162306 281551 162362 281560
rect 162216 272536 162268 272542
rect 162216 272478 162268 272484
rect 162124 269884 162176 269890
rect 162124 269826 162176 269832
rect 162122 265160 162178 265169
rect 162122 265095 162178 265104
rect 161112 251184 161164 251190
rect 161112 251126 161164 251132
rect 161020 146940 161072 146946
rect 161020 146882 161072 146888
rect 161032 142154 161060 146882
rect 160940 142126 161060 142154
rect 160940 120086 160968 142126
rect 160928 120080 160980 120086
rect 160928 120022 160980 120028
rect 160836 31068 160888 31074
rect 160836 31010 160888 31016
rect 160744 26920 160796 26926
rect 160744 26862 160796 26868
rect 162136 25566 162164 265095
rect 162228 156058 162256 272478
rect 162320 169046 162348 281551
rect 163516 277302 163544 318815
rect 163504 277296 163556 277302
rect 163504 277238 163556 277244
rect 163504 262268 163556 262274
rect 163504 262210 163556 262216
rect 162308 169040 162360 169046
rect 162308 168982 162360 168988
rect 162216 156052 162268 156058
rect 162216 155994 162268 156000
rect 162228 151814 162256 155994
rect 162228 151786 162348 151814
rect 162216 148368 162268 148374
rect 162216 148310 162268 148316
rect 162228 106321 162256 148310
rect 162320 122806 162348 151786
rect 162308 122800 162360 122806
rect 162308 122742 162360 122748
rect 162214 106312 162270 106321
rect 162214 106247 162270 106256
rect 163516 71058 163544 262210
rect 163608 240106 163636 390526
rect 164976 389292 165028 389298
rect 164976 389234 165028 389240
rect 164884 354000 164936 354006
rect 164884 353942 164936 353948
rect 164896 271862 164924 353942
rect 164148 271856 164200 271862
rect 164148 271798 164200 271804
rect 164884 271856 164936 271862
rect 164884 271798 164936 271804
rect 163686 262848 163742 262857
rect 163686 262783 163742 262792
rect 163596 240100 163648 240106
rect 163596 240042 163648 240048
rect 163700 222902 163728 262783
rect 164056 240100 164108 240106
rect 164056 240042 164108 240048
rect 164068 239426 164096 240042
rect 164056 239420 164108 239426
rect 164056 239362 164108 239368
rect 163688 222896 163740 222902
rect 163688 222838 163740 222844
rect 164160 109002 164188 271798
rect 164884 260908 164936 260914
rect 164884 260850 164936 260856
rect 164148 108996 164200 109002
rect 164148 108938 164200 108944
rect 164160 108322 164188 108938
rect 164148 108316 164200 108322
rect 164148 108258 164200 108264
rect 163504 71052 163556 71058
rect 163504 70994 163556 71000
rect 164896 68338 164924 260850
rect 164988 240038 165016 389234
rect 166276 377369 166304 406263
rect 166354 388920 166410 388929
rect 166354 388855 166410 388864
rect 166262 377360 166318 377369
rect 166262 377295 166318 377304
rect 165528 279472 165580 279478
rect 165528 279414 165580 279420
rect 164976 240032 165028 240038
rect 164976 239974 165028 239980
rect 165540 146402 165568 279414
rect 166264 248532 166316 248538
rect 166264 248474 166316 248480
rect 165528 146396 165580 146402
rect 165528 146338 165580 146344
rect 165540 144226 165568 146338
rect 165528 144220 165580 144226
rect 165528 144162 165580 144168
rect 164884 68332 164936 68338
rect 164884 68274 164936 68280
rect 166276 29646 166304 248474
rect 166368 245002 166396 388855
rect 166446 290456 166502 290465
rect 166446 290391 166502 290400
rect 166460 289921 166488 290391
rect 166446 289912 166502 289921
rect 166446 289847 166502 289856
rect 166356 244996 166408 245002
rect 166356 244938 166408 244944
rect 166460 168366 166488 289847
rect 166920 288386 166948 460974
rect 168288 452736 168340 452742
rect 168288 452678 168340 452684
rect 167644 417444 167696 417450
rect 167644 417386 167696 417392
rect 167656 326398 167684 417386
rect 167644 326392 167696 326398
rect 167644 326334 167696 326340
rect 167656 325694 167684 326334
rect 167656 325666 167776 325694
rect 167642 322960 167698 322969
rect 167642 322895 167698 322904
rect 167656 298790 167684 322895
rect 167748 311982 167776 325666
rect 168300 322969 168328 452678
rect 169024 448588 169076 448594
rect 169024 448530 169076 448536
rect 169036 427106 169064 448530
rect 170404 447840 170456 447846
rect 170404 447782 170456 447788
rect 169666 443048 169722 443057
rect 169666 442983 169722 442992
rect 169024 427100 169076 427106
rect 169024 427042 169076 427048
rect 169024 405748 169076 405754
rect 169024 405690 169076 405696
rect 168378 381712 168434 381721
rect 168378 381647 168434 381656
rect 168392 375290 168420 381647
rect 169036 375329 169064 405690
rect 169022 375320 169078 375329
rect 168380 375284 168432 375290
rect 169022 375255 169078 375264
rect 168380 375226 168432 375232
rect 168286 322960 168342 322969
rect 168286 322895 168342 322904
rect 167736 311976 167788 311982
rect 167736 311918 167788 311924
rect 168288 311976 168340 311982
rect 168288 311918 168340 311924
rect 167644 298784 167696 298790
rect 167644 298726 167696 298732
rect 166540 288380 166592 288386
rect 166540 288322 166592 288328
rect 166908 288380 166960 288386
rect 166908 288322 166960 288328
rect 166552 287774 166580 288322
rect 166540 287768 166592 287774
rect 166540 287710 166592 287716
rect 168300 281518 168328 311918
rect 168288 281512 168340 281518
rect 168288 281454 168340 281460
rect 167736 280832 167788 280838
rect 167736 280774 167788 280780
rect 167644 258188 167696 258194
rect 167644 258130 167696 258136
rect 166538 238096 166594 238105
rect 166538 238031 166594 238040
rect 166552 237425 166580 238031
rect 166538 237416 166594 237425
rect 166538 237351 166594 237360
rect 166906 237416 166962 237425
rect 166906 237351 166962 237360
rect 166448 168360 166500 168366
rect 166448 168302 166500 168308
rect 166460 167686 166488 168302
rect 166448 167680 166500 167686
rect 166448 167622 166500 167628
rect 166920 107642 166948 237351
rect 166908 107636 166960 107642
rect 166908 107578 166960 107584
rect 167656 75177 167684 258130
rect 167748 111790 167776 280774
rect 168288 265668 168340 265674
rect 168288 265610 168340 265616
rect 168300 237318 168328 265610
rect 168392 251870 168420 375226
rect 169680 351218 169708 442983
rect 170416 422958 170444 447782
rect 172428 446412 172480 446418
rect 172428 446354 172480 446360
rect 171048 431248 171100 431254
rect 171048 431190 171100 431196
rect 170404 422952 170456 422958
rect 170404 422894 170456 422900
rect 170956 422952 171008 422958
rect 170956 422894 171008 422900
rect 170404 407176 170456 407182
rect 170404 407118 170456 407124
rect 170416 373998 170444 407118
rect 170404 373992 170456 373998
rect 170404 373934 170456 373940
rect 170494 364984 170550 364993
rect 170494 364919 170550 364928
rect 170508 364410 170536 364919
rect 170496 364404 170548 364410
rect 170496 364346 170548 364352
rect 169668 351212 169720 351218
rect 169668 351154 169720 351160
rect 169576 349852 169628 349858
rect 169576 349794 169628 349800
rect 169588 282878 169616 349794
rect 169668 336048 169720 336054
rect 169668 335990 169720 335996
rect 168472 282872 168524 282878
rect 168472 282814 168524 282820
rect 169576 282872 169628 282878
rect 169576 282814 169628 282820
rect 168484 282198 168512 282814
rect 168472 282192 168524 282198
rect 168472 282134 168524 282140
rect 168470 281616 168526 281625
rect 168470 281551 168526 281560
rect 168484 280158 168512 281551
rect 168472 280152 168524 280158
rect 168472 280094 168524 280100
rect 169024 262336 169076 262342
rect 169024 262278 169076 262284
rect 168380 251864 168432 251870
rect 168380 251806 168432 251812
rect 168288 237312 168340 237318
rect 168288 237254 168340 237260
rect 168300 152561 168328 237254
rect 168286 152552 168342 152561
rect 168286 152487 168342 152496
rect 167736 111784 167788 111790
rect 167736 111726 167788 111732
rect 167748 81326 167776 111726
rect 167736 81320 167788 81326
rect 167736 81262 167788 81268
rect 167642 75168 167698 75177
rect 167642 75103 167698 75112
rect 166264 29640 166316 29646
rect 166264 29582 166316 29588
rect 162124 25560 162176 25566
rect 162124 25502 162176 25508
rect 169036 19990 169064 262278
rect 169116 259684 169168 259690
rect 169116 259626 169168 259632
rect 169128 225622 169156 259626
rect 169116 225616 169168 225622
rect 169116 225558 169168 225564
rect 169128 203590 169156 225558
rect 169116 203584 169168 203590
rect 169116 203526 169168 203532
rect 169114 180024 169170 180033
rect 169114 179959 169170 179968
rect 169128 135930 169156 179959
rect 169208 137284 169260 137290
rect 169208 137226 169260 137232
rect 169116 135924 169168 135930
rect 169116 135866 169168 135872
rect 169220 124166 169248 137226
rect 169208 124160 169260 124166
rect 169208 124102 169260 124108
rect 169680 102134 169708 335990
rect 169760 289808 169812 289814
rect 169760 289750 169812 289756
rect 169772 289105 169800 289750
rect 169758 289096 169814 289105
rect 169758 289031 169814 289040
rect 169760 286340 169812 286346
rect 169760 286282 169812 286288
rect 169772 285734 169800 286282
rect 169760 285728 169812 285734
rect 169760 285670 169812 285676
rect 170404 259480 170456 259486
rect 170404 259422 170456 259428
rect 170128 115932 170180 115938
rect 170128 115874 170180 115880
rect 170140 115258 170168 115874
rect 170128 115252 170180 115258
rect 170128 115194 170180 115200
rect 169668 102128 169720 102134
rect 169668 102070 169720 102076
rect 169680 101454 169708 102070
rect 169668 101448 169720 101454
rect 169668 101390 169720 101396
rect 169024 19984 169076 19990
rect 169024 19926 169076 19932
rect 170416 8974 170444 259422
rect 170508 215286 170536 364346
rect 170968 314945 170996 422894
rect 170678 314936 170734 314945
rect 170678 314871 170734 314880
rect 170954 314936 171010 314945
rect 170954 314871 171010 314880
rect 170588 286340 170640 286346
rect 170588 286282 170640 286288
rect 170496 215280 170548 215286
rect 170496 215222 170548 215228
rect 170600 141438 170628 286282
rect 170692 259690 170720 314871
rect 171060 289814 171088 431190
rect 171968 313404 172020 313410
rect 171968 313346 172020 313352
rect 171140 307896 171192 307902
rect 171140 307838 171192 307844
rect 171152 304366 171180 307838
rect 171140 304360 171192 304366
rect 171140 304302 171192 304308
rect 171048 289808 171100 289814
rect 171048 289750 171100 289756
rect 171876 288312 171928 288318
rect 171876 288254 171928 288260
rect 171888 287706 171916 288254
rect 171876 287700 171928 287706
rect 171876 287642 171928 287648
rect 171876 281512 171928 281518
rect 171876 281454 171928 281460
rect 170770 260128 170826 260137
rect 170770 260063 170826 260072
rect 170680 259684 170732 259690
rect 170680 259626 170732 259632
rect 170784 224330 170812 260063
rect 171784 256760 171836 256766
rect 171784 256702 171836 256708
rect 171140 239420 171192 239426
rect 171140 239362 171192 239368
rect 170772 224324 170824 224330
rect 170772 224266 170824 224272
rect 171048 220856 171100 220862
rect 171048 220798 171100 220804
rect 170588 141432 170640 141438
rect 170588 141374 170640 141380
rect 171060 115258 171088 220798
rect 171048 115252 171100 115258
rect 171048 115194 171100 115200
rect 171152 99362 171180 239362
rect 171060 99334 171180 99362
rect 171060 98122 171088 99334
rect 171048 98116 171100 98122
rect 171048 98058 171100 98064
rect 171060 93226 171088 98058
rect 171048 93220 171100 93226
rect 171048 93162 171100 93168
rect 171796 76566 171824 256702
rect 171888 136610 171916 281454
rect 171980 257378 172008 313346
rect 172440 288318 172468 446354
rect 173164 419620 173216 419626
rect 173164 419562 173216 419568
rect 173176 309806 173204 419562
rect 173820 384985 173848 702714
rect 177948 702568 178000 702574
rect 177948 702510 178000 702516
rect 175186 457056 175242 457065
rect 175186 456991 175242 457000
rect 175200 456822 175228 456991
rect 175188 456816 175240 456822
rect 175188 456758 175240 456764
rect 174544 398880 174596 398886
rect 174544 398822 174596 398828
rect 174556 386374 174584 398822
rect 174544 386368 174596 386374
rect 174544 386310 174596 386316
rect 173254 384976 173310 384985
rect 173254 384911 173310 384920
rect 173806 384976 173862 384985
rect 173806 384911 173862 384920
rect 173268 368393 173296 384911
rect 173254 368384 173310 368393
rect 173254 368319 173310 368328
rect 172612 309800 172664 309806
rect 172612 309742 172664 309748
rect 173164 309800 173216 309806
rect 173164 309742 173216 309748
rect 172428 288312 172480 288318
rect 172428 288254 172480 288260
rect 172520 272604 172572 272610
rect 172520 272546 172572 272552
rect 171968 257372 172020 257378
rect 171968 257314 172020 257320
rect 171876 136604 171928 136610
rect 171876 136546 171928 136552
rect 172532 135289 172560 272546
rect 172624 269793 172652 309742
rect 172610 269784 172666 269793
rect 172610 269719 172666 269728
rect 173164 263696 173216 263702
rect 173164 263638 173216 263644
rect 172612 240168 172664 240174
rect 172612 240110 172664 240116
rect 172624 235657 172652 240110
rect 172610 235648 172666 235657
rect 172610 235583 172666 235592
rect 172518 135280 172574 135289
rect 172518 135215 172574 135224
rect 171784 76560 171836 76566
rect 171784 76502 171836 76508
rect 170404 8968 170456 8974
rect 170404 8910 170456 8916
rect 159364 7608 159416 7614
rect 159364 7550 159416 7556
rect 173176 4894 173204 263638
rect 173268 240961 173296 368319
rect 173348 340944 173400 340950
rect 173348 340886 173400 340892
rect 173254 240952 173310 240961
rect 173254 240887 173310 240896
rect 173360 220862 173388 340886
rect 174556 327214 174584 386310
rect 174726 329896 174782 329905
rect 174726 329831 174782 329840
rect 174544 327208 174596 327214
rect 174544 327150 174596 327156
rect 174556 313410 174584 327150
rect 174636 324352 174688 324358
rect 174636 324294 174688 324300
rect 174544 313404 174596 313410
rect 174544 313346 174596 313352
rect 174544 310548 174596 310554
rect 174544 310490 174596 310496
rect 173808 281580 173860 281586
rect 173808 281522 173860 281528
rect 173820 278730 173848 281522
rect 173808 278724 173860 278730
rect 173808 278666 173860 278672
rect 174556 278050 174584 310490
rect 174648 296002 174676 324294
rect 174636 295996 174688 296002
rect 174636 295938 174688 295944
rect 174636 278724 174688 278730
rect 174636 278666 174688 278672
rect 174544 278044 174596 278050
rect 174544 277986 174596 277992
rect 174648 277438 174676 278666
rect 174636 277432 174688 277438
rect 174636 277374 174688 277380
rect 173808 272604 173860 272610
rect 173808 272546 173860 272552
rect 173820 271930 173848 272546
rect 173808 271924 173860 271930
rect 173808 271866 173860 271872
rect 174544 255332 174596 255338
rect 174544 255274 174596 255280
rect 173348 220856 173400 220862
rect 173348 220798 173400 220804
rect 173254 220280 173310 220289
rect 173254 220215 173310 220224
rect 173268 191146 173296 220215
rect 173256 191140 173308 191146
rect 173256 191082 173308 191088
rect 173268 95305 173296 191082
rect 173346 144256 173402 144265
rect 173346 144191 173402 144200
rect 173360 123457 173388 144191
rect 173806 135280 173862 135289
rect 173806 135215 173862 135224
rect 173820 133890 173848 135215
rect 173808 133884 173860 133890
rect 173808 133826 173860 133832
rect 173346 123448 173402 123457
rect 173346 123383 173402 123392
rect 173254 95296 173310 95305
rect 173254 95231 173310 95240
rect 174556 15910 174584 255274
rect 174648 140078 174676 277374
rect 174740 253230 174768 329831
rect 175200 324358 175228 456758
rect 176568 448588 176620 448594
rect 176568 448530 176620 448536
rect 175188 324352 175240 324358
rect 175188 324294 175240 324300
rect 176580 305017 176608 448530
rect 176660 444440 176712 444446
rect 176660 444382 176712 444388
rect 176014 305008 176070 305017
rect 176014 304943 176070 304952
rect 176566 305008 176622 305017
rect 176566 304943 176622 304952
rect 175924 300960 175976 300966
rect 175924 300902 175976 300908
rect 175936 280838 175964 300902
rect 175924 280832 175976 280838
rect 175924 280774 175976 280780
rect 175924 270564 175976 270570
rect 175924 270506 175976 270512
rect 174820 255400 174872 255406
rect 174820 255342 174872 255348
rect 174728 253224 174780 253230
rect 174728 253166 174780 253172
rect 174832 238066 174860 255342
rect 174820 238060 174872 238066
rect 174820 238002 174872 238008
rect 175186 236736 175242 236745
rect 175186 236671 175242 236680
rect 175200 209681 175228 236671
rect 175186 209672 175242 209681
rect 175186 209607 175242 209616
rect 175200 208418 175228 209607
rect 175188 208412 175240 208418
rect 175188 208354 175240 208360
rect 174636 140072 174688 140078
rect 174636 140014 174688 140020
rect 174648 139466 174676 140014
rect 174636 139460 174688 139466
rect 174636 139402 174688 139408
rect 174636 134564 174688 134570
rect 174636 134506 174688 134512
rect 174648 106282 174676 134506
rect 174636 106276 174688 106282
rect 174636 106218 174688 106224
rect 174636 103556 174688 103562
rect 174636 103498 174688 103504
rect 174648 73098 174676 103498
rect 174636 73092 174688 73098
rect 174636 73034 174688 73040
rect 175936 28286 175964 270506
rect 176028 267034 176056 304943
rect 176672 294001 176700 444382
rect 176752 427100 176804 427106
rect 176752 427042 176804 427048
rect 176764 426494 176792 427042
rect 176752 426488 176804 426494
rect 176752 426430 176804 426436
rect 177856 426488 177908 426494
rect 177856 426430 177908 426436
rect 176752 397452 176804 397458
rect 176752 397394 176804 397400
rect 176764 396681 176792 397394
rect 176750 396672 176806 396681
rect 176750 396607 176806 396616
rect 177868 316062 177896 426430
rect 177960 397458 177988 702510
rect 187608 576904 187660 576910
rect 187608 576846 187660 576852
rect 186964 463752 187016 463758
rect 184202 463720 184258 463729
rect 186964 463694 187016 463700
rect 184202 463655 184258 463664
rect 180062 461136 180118 461145
rect 180062 461071 180118 461080
rect 178682 454064 178738 454073
rect 178682 453999 178738 454008
rect 178696 434722 178724 453999
rect 178960 447840 179012 447846
rect 178960 447782 179012 447788
rect 178972 447166 179000 447782
rect 178960 447160 179012 447166
rect 178960 447102 179012 447108
rect 179236 447160 179288 447166
rect 179236 447102 179288 447108
rect 178684 434716 178736 434722
rect 178684 434658 178736 434664
rect 177948 397452 178000 397458
rect 177948 397394 178000 397400
rect 178684 351212 178736 351218
rect 178684 351154 178736 351160
rect 177948 345704 178000 345710
rect 177948 345646 178000 345652
rect 177856 316056 177908 316062
rect 177856 315998 177908 316004
rect 177302 309360 177358 309369
rect 177302 309295 177358 309304
rect 176658 293992 176714 294001
rect 176658 293927 176714 293936
rect 177210 293992 177266 294001
rect 177210 293927 177266 293936
rect 177224 287054 177252 293927
rect 177316 293282 177344 309295
rect 177304 293276 177356 293282
rect 177304 293218 177356 293224
rect 177224 287026 177344 287054
rect 177316 284986 177344 287026
rect 177304 284980 177356 284986
rect 177304 284922 177356 284928
rect 176568 284368 176620 284374
rect 176568 284310 176620 284316
rect 176016 267028 176068 267034
rect 176016 266970 176068 266976
rect 176476 251932 176528 251938
rect 176476 251874 176528 251880
rect 176488 233238 176516 251874
rect 176476 233232 176528 233238
rect 176476 233174 176528 233180
rect 176488 233034 176516 233174
rect 176016 233028 176068 233034
rect 176016 232970 176068 232976
rect 176476 233028 176528 233034
rect 176476 232970 176528 232976
rect 176028 205698 176056 232970
rect 176016 205692 176068 205698
rect 176016 205634 176068 205640
rect 176028 126274 176056 205634
rect 176580 160206 176608 284310
rect 177316 272542 177344 284922
rect 177868 274650 177896 315998
rect 177856 274644 177908 274650
rect 177856 274586 177908 274592
rect 177304 272536 177356 272542
rect 177304 272478 177356 272484
rect 177396 271992 177448 271998
rect 177396 271934 177448 271940
rect 177304 255400 177356 255406
rect 177304 255342 177356 255348
rect 176568 160200 176620 160206
rect 176568 160142 176620 160148
rect 176580 159390 176608 160142
rect 176568 159384 176620 159390
rect 176568 159326 176620 159332
rect 176016 126268 176068 126274
rect 176016 126210 176068 126216
rect 175924 28280 175976 28286
rect 175924 28222 175976 28228
rect 174544 15904 174596 15910
rect 174544 15846 174596 15852
rect 177316 13122 177344 255342
rect 177408 238134 177436 271934
rect 177488 251864 177540 251870
rect 177488 251806 177540 251812
rect 177500 238754 177528 251806
rect 177960 240145 177988 345646
rect 178040 300824 178092 300830
rect 178040 300766 178092 300772
rect 178052 299606 178080 300766
rect 178040 299600 178092 299606
rect 178040 299542 178092 299548
rect 178052 284374 178080 299542
rect 178696 291961 178724 351154
rect 179248 318850 179276 447102
rect 180076 438938 180104 461071
rect 183466 456920 183522 456929
rect 183466 456855 183522 456864
rect 180154 455832 180210 455841
rect 180154 455767 180210 455776
rect 180064 438932 180116 438938
rect 180064 438874 180116 438880
rect 179328 416152 179380 416158
rect 179328 416094 179380 416100
rect 178776 318844 178828 318850
rect 178776 318786 178828 318792
rect 179236 318844 179288 318850
rect 179236 318786 179288 318792
rect 178788 300830 178816 318786
rect 178776 300824 178828 300830
rect 178776 300766 178828 300772
rect 178682 291952 178738 291961
rect 178682 291887 178738 291896
rect 178696 287054 178724 291887
rect 178696 287026 178816 287054
rect 178040 284368 178092 284374
rect 178040 284310 178092 284316
rect 178684 242956 178736 242962
rect 178684 242898 178736 242904
rect 177946 240136 178002 240145
rect 177946 240071 178002 240080
rect 177500 238726 177988 238754
rect 177396 238128 177448 238134
rect 177396 238070 177448 238076
rect 177960 235929 177988 238726
rect 177946 235920 178002 235929
rect 177946 235855 178002 235864
rect 177396 224256 177448 224262
rect 177396 224198 177448 224204
rect 177408 215966 177436 224198
rect 177396 215960 177448 215966
rect 177396 215902 177448 215908
rect 177394 144936 177450 144945
rect 177394 144871 177450 144880
rect 177408 111790 177436 144871
rect 177396 111784 177448 111790
rect 177396 111726 177448 111732
rect 177396 108316 177448 108322
rect 177396 108258 177448 108264
rect 177408 79966 177436 108258
rect 177960 92449 177988 235855
rect 178040 120760 178092 120766
rect 178040 120702 178092 120708
rect 178052 117978 178080 120702
rect 178040 117972 178092 117978
rect 178040 117914 178092 117920
rect 177946 92440 178002 92449
rect 177946 92375 178002 92384
rect 177396 79960 177448 79966
rect 177396 79902 177448 79908
rect 177304 13116 177356 13122
rect 177304 13058 177356 13064
rect 173164 4888 173216 4894
rect 173164 4830 173216 4836
rect 143540 3528 143592 3534
rect 143540 3470 143592 3476
rect 144828 3528 144880 3534
rect 144828 3470 144880 3476
rect 147128 3528 147180 3534
rect 147128 3470 147180 3476
rect 147588 3528 147640 3534
rect 147588 3470 147640 3476
rect 140044 2780 140096 2786
rect 140044 2722 140096 2728
rect 142988 2780 143040 2786
rect 142988 2722 143040 2728
rect 140056 480 140084 2722
rect 143552 480 143580 3470
rect 147140 480 147168 3470
rect 178696 2106 178724 242898
rect 178788 155242 178816 287026
rect 178866 284336 178922 284345
rect 178866 284271 178922 284280
rect 178880 239737 178908 284271
rect 178866 239728 178922 239737
rect 178866 239663 178922 239672
rect 179340 228993 179368 416094
rect 179510 388512 179566 388521
rect 179510 388447 179566 388456
rect 179524 387841 179552 388447
rect 179510 387832 179566 387841
rect 179510 387767 179566 387776
rect 179524 373994 179552 387767
rect 179432 373966 179552 373994
rect 179432 251938 179460 373966
rect 179420 251932 179472 251938
rect 179420 251874 179472 251880
rect 179326 228984 179382 228993
rect 179326 228919 179382 228928
rect 180076 228313 180104 438874
rect 180168 431254 180196 455767
rect 181534 447944 181590 447953
rect 181534 447879 181590 447888
rect 180156 431248 180208 431254
rect 180156 431190 180208 431196
rect 181444 425128 181496 425134
rect 181444 425070 181496 425076
rect 180156 419552 180208 419558
rect 180156 419494 180208 419500
rect 180168 387734 180196 419494
rect 180248 397588 180300 397594
rect 180248 397530 180300 397536
rect 180156 387728 180208 387734
rect 180156 387670 180208 387676
rect 180260 373994 180288 397530
rect 180168 373966 180288 373994
rect 180168 369753 180196 373966
rect 180154 369744 180210 369753
rect 180154 369679 180210 369688
rect 180168 329186 180196 369679
rect 180156 329180 180208 329186
rect 180156 329122 180208 329128
rect 180156 320204 180208 320210
rect 180156 320146 180208 320152
rect 180168 286346 180196 320146
rect 180248 302252 180300 302258
rect 180248 302194 180300 302200
rect 180156 286340 180208 286346
rect 180156 286282 180208 286288
rect 180260 273873 180288 302194
rect 181456 285569 181484 425070
rect 181548 424386 181576 447879
rect 181536 424380 181588 424386
rect 181536 424322 181588 424328
rect 182916 404388 182968 404394
rect 182916 404330 182968 404336
rect 181536 394732 181588 394738
rect 181536 394674 181588 394680
rect 181548 375290 181576 394674
rect 181536 375284 181588 375290
rect 181536 375226 181588 375232
rect 182086 317384 182142 317393
rect 182086 317319 182142 317328
rect 182100 316713 182128 317319
rect 182086 316704 182142 316713
rect 182086 316639 182142 316648
rect 181536 311908 181588 311914
rect 181536 311850 181588 311856
rect 181548 304298 181576 311850
rect 181536 304292 181588 304298
rect 181536 304234 181588 304240
rect 181534 300112 181590 300121
rect 181534 300047 181590 300056
rect 181548 291825 181576 300047
rect 181534 291816 181590 291825
rect 181534 291751 181590 291760
rect 181442 285560 181498 285569
rect 181442 285495 181498 285504
rect 180246 273864 180302 273873
rect 180246 273799 180302 273808
rect 180156 267776 180208 267782
rect 180156 267718 180208 267724
rect 180062 228304 180118 228313
rect 180062 228239 180118 228248
rect 180062 226264 180118 226273
rect 180062 226199 180118 226208
rect 180076 215937 180104 226199
rect 180168 217297 180196 267718
rect 181456 265033 181484 285495
rect 181442 265024 181498 265033
rect 181442 264959 181498 264968
rect 180616 257372 180668 257378
rect 180616 257314 180668 257320
rect 180248 240780 180300 240786
rect 180248 240722 180300 240728
rect 180260 237386 180288 240722
rect 180248 237380 180300 237386
rect 180248 237322 180300 237328
rect 180260 230489 180288 237322
rect 180246 230480 180302 230489
rect 180246 230415 180302 230424
rect 180260 219434 180288 230415
rect 180628 226273 180656 257314
rect 181444 252612 181496 252618
rect 181444 252554 181496 252560
rect 180614 226264 180670 226273
rect 180614 226199 180670 226208
rect 180260 219406 180748 219434
rect 180154 217288 180210 217297
rect 180154 217223 180210 217232
rect 180062 215928 180118 215937
rect 180062 215863 180118 215872
rect 180076 209774 180104 215863
rect 180076 209746 180196 209774
rect 180064 208412 180116 208418
rect 180064 208354 180116 208360
rect 178868 203584 178920 203590
rect 178868 203526 178920 203532
rect 178776 155236 178828 155242
rect 178776 155178 178828 155184
rect 178788 121446 178816 155178
rect 178776 121440 178828 121446
rect 178776 121382 178828 121388
rect 178880 114510 178908 203526
rect 179328 117972 179380 117978
rect 179328 117914 179380 117920
rect 178868 114504 178920 114510
rect 178868 114446 178920 114452
rect 178776 113212 178828 113218
rect 178776 113154 178828 113160
rect 178788 84017 178816 113154
rect 178774 84008 178830 84017
rect 178774 83943 178830 83952
rect 179340 39370 179368 117914
rect 179420 92404 179472 92410
rect 179420 92346 179472 92352
rect 179432 92313 179460 92346
rect 179418 92304 179474 92313
rect 179418 92239 179474 92248
rect 180076 86737 180104 208354
rect 180168 145586 180196 209746
rect 180248 150544 180300 150550
rect 180248 150486 180300 150492
rect 180156 145580 180208 145586
rect 180156 145522 180208 145528
rect 180156 135312 180208 135318
rect 180156 135254 180208 135260
rect 180062 86728 180118 86737
rect 180062 86663 180118 86672
rect 180168 62830 180196 135254
rect 180260 125594 180288 150486
rect 180248 125588 180300 125594
rect 180248 125530 180300 125536
rect 180616 123480 180668 123486
rect 180616 123422 180668 123428
rect 180156 62824 180208 62830
rect 180156 62766 180208 62772
rect 179328 39364 179380 39370
rect 179328 39306 179380 39312
rect 180628 37942 180656 123422
rect 180720 92410 180748 219406
rect 180708 92404 180760 92410
rect 180708 92346 180760 92352
rect 181456 58682 181484 252554
rect 181534 246256 181590 246265
rect 181534 246191 181590 246200
rect 181548 231849 181576 246191
rect 182100 238649 182128 316639
rect 182824 303816 182876 303822
rect 182824 303758 182876 303764
rect 182180 274644 182232 274650
rect 182180 274586 182232 274592
rect 182086 238640 182142 238649
rect 182086 238575 182142 238584
rect 181534 231840 181590 231849
rect 181534 231775 181590 231784
rect 181548 210361 181576 231775
rect 182192 230518 182220 274586
rect 182180 230512 182232 230518
rect 182180 230454 182232 230460
rect 181534 210352 181590 210361
rect 181534 210287 181590 210296
rect 181548 209774 181576 210287
rect 181548 209746 181668 209774
rect 181534 143576 181590 143585
rect 181534 143511 181590 143520
rect 181548 129742 181576 143511
rect 181536 129736 181588 129742
rect 181536 129678 181588 129684
rect 181536 127016 181588 127022
rect 181536 126958 181588 126964
rect 181548 122806 181576 126958
rect 181536 122800 181588 122806
rect 181536 122742 181588 122748
rect 181444 58676 181496 58682
rect 181444 58618 181496 58624
rect 180616 37936 180668 37942
rect 180616 37878 180668 37884
rect 181548 13122 181576 122742
rect 181640 121990 181668 209746
rect 182088 160132 182140 160138
rect 182088 160074 182140 160080
rect 182100 152590 182128 160074
rect 182088 152584 182140 152590
rect 182088 152526 182140 152532
rect 182364 122868 182416 122874
rect 182364 122810 182416 122816
rect 181628 121984 181680 121990
rect 181628 121926 181680 121932
rect 182376 120057 182404 122810
rect 182362 120048 182418 120057
rect 182362 119983 182418 119992
rect 182836 77897 182864 303758
rect 182928 291786 182956 404330
rect 183480 318753 183508 456855
rect 183560 367056 183612 367062
rect 183560 366998 183612 367004
rect 183572 366858 183600 366998
rect 183560 366852 183612 366858
rect 183560 366794 183612 366800
rect 183466 318744 183522 318753
rect 183466 318679 183522 318688
rect 183480 318073 183508 318679
rect 183466 318064 183522 318073
rect 183466 317999 183522 318008
rect 183008 317552 183060 317558
rect 183008 317494 183060 317500
rect 182916 291780 182968 291786
rect 182916 291722 182968 291728
rect 182928 251841 182956 291722
rect 183020 274582 183048 317494
rect 183466 291952 183522 291961
rect 183466 291887 183522 291896
rect 183480 291854 183508 291887
rect 183468 291848 183520 291854
rect 183468 291790 183520 291796
rect 183008 274576 183060 274582
rect 183008 274518 183060 274524
rect 183572 257378 183600 366794
rect 184216 317393 184244 463655
rect 184848 459672 184900 459678
rect 184848 459614 184900 459620
rect 184388 451308 184440 451314
rect 184388 451250 184440 451256
rect 184296 418192 184348 418198
rect 184296 418134 184348 418140
rect 184308 380866 184336 418134
rect 184400 417450 184428 451250
rect 184388 417444 184440 417450
rect 184388 417386 184440 417392
rect 184388 400240 184440 400246
rect 184388 400182 184440 400188
rect 184296 380860 184348 380866
rect 184296 380802 184348 380808
rect 184400 367062 184428 400182
rect 184388 367056 184440 367062
rect 184388 366998 184440 367004
rect 184202 317384 184258 317393
rect 184202 317319 184258 317328
rect 184202 308136 184258 308145
rect 184202 308071 184258 308080
rect 184216 280809 184244 308071
rect 184860 294166 184888 459614
rect 185674 458416 185730 458425
rect 185674 458351 185730 458360
rect 185584 449200 185636 449206
rect 185584 449142 185636 449148
rect 184938 320104 184994 320113
rect 184938 320039 184994 320048
rect 184848 294160 184900 294166
rect 184848 294102 184900 294108
rect 184860 290465 184888 294102
rect 184846 290456 184902 290465
rect 184846 290391 184902 290400
rect 184848 290352 184900 290358
rect 184848 290294 184900 290300
rect 184860 289882 184888 290294
rect 184848 289876 184900 289882
rect 184848 289818 184900 289824
rect 184296 281580 184348 281586
rect 184296 281522 184348 281528
rect 184202 280800 184258 280809
rect 184202 280735 184258 280744
rect 184308 271862 184336 281522
rect 184296 271856 184348 271862
rect 184296 271798 184348 271804
rect 184204 264988 184256 264994
rect 184204 264930 184256 264936
rect 183560 257372 183612 257378
rect 183560 257314 183612 257320
rect 182914 251832 182970 251841
rect 182914 251767 182970 251776
rect 183008 247104 183060 247110
rect 183008 247046 183060 247052
rect 182916 230512 182968 230518
rect 182916 230454 182968 230460
rect 182928 117230 182956 230454
rect 183020 214577 183048 247046
rect 184216 218822 184244 264930
rect 184296 263628 184348 263634
rect 184296 263570 184348 263576
rect 184308 236881 184336 263570
rect 184860 246362 184888 289818
rect 184952 265674 184980 320039
rect 185596 289134 185624 449142
rect 185688 320113 185716 458351
rect 186976 432041 187004 463694
rect 187054 450120 187110 450129
rect 187054 450055 187110 450064
rect 187068 437481 187096 450055
rect 187054 437472 187110 437481
rect 187054 437407 187110 437416
rect 186962 432032 187018 432041
rect 186962 431967 187018 431976
rect 187424 431996 187476 432002
rect 187424 431938 187476 431944
rect 186962 418296 187018 418305
rect 186962 418231 187018 418240
rect 185768 403028 185820 403034
rect 185768 402970 185820 402976
rect 185780 379370 185808 402970
rect 186976 386374 187004 418231
rect 187054 400888 187110 400897
rect 187054 400823 187110 400832
rect 186964 386368 187016 386374
rect 186964 386310 187016 386316
rect 187068 386209 187096 400823
rect 187054 386200 187110 386209
rect 187054 386135 187110 386144
rect 186320 384328 186372 384334
rect 186320 384270 186372 384276
rect 185768 379364 185820 379370
rect 185768 379306 185820 379312
rect 185674 320104 185730 320113
rect 185674 320039 185730 320048
rect 185674 309496 185730 309505
rect 185674 309431 185730 309440
rect 185584 289128 185636 289134
rect 185584 289070 185636 289076
rect 185596 287054 185624 289070
rect 185504 287026 185624 287054
rect 185504 277370 185532 287026
rect 185688 277394 185716 309431
rect 185492 277364 185544 277370
rect 185492 277306 185544 277312
rect 185596 277366 185716 277394
rect 185596 276010 185624 277366
rect 185584 276004 185636 276010
rect 185584 275946 185636 275952
rect 184940 265668 184992 265674
rect 184940 265610 184992 265616
rect 184848 246356 184900 246362
rect 184848 246298 184900 246304
rect 184480 244996 184532 245002
rect 184480 244938 184532 244944
rect 184388 243568 184440 243574
rect 184388 243510 184440 243516
rect 184294 236872 184350 236881
rect 184294 236807 184350 236816
rect 184294 232656 184350 232665
rect 184294 232591 184350 232600
rect 184308 228993 184336 232591
rect 184400 231810 184428 243510
rect 184492 234569 184520 244938
rect 184478 234560 184534 234569
rect 184478 234495 184534 234504
rect 184388 231804 184440 231810
rect 184388 231746 184440 231752
rect 184294 228984 184350 228993
rect 184294 228919 184350 228928
rect 184308 227769 184336 228919
rect 184294 227760 184350 227769
rect 184294 227695 184350 227704
rect 184204 218816 184256 218822
rect 184204 218758 184256 218764
rect 183006 214568 183062 214577
rect 183006 214503 183062 214512
rect 184296 186992 184348 186998
rect 184296 186934 184348 186940
rect 183008 155304 183060 155310
rect 183008 155246 183060 155252
rect 183020 148442 183048 155246
rect 184308 152522 184336 186934
rect 184296 152516 184348 152522
rect 184296 152458 184348 152464
rect 184204 151836 184256 151842
rect 184204 151778 184256 151784
rect 183008 148436 183060 148442
rect 183008 148378 183060 148384
rect 183006 147112 183062 147121
rect 183006 147047 183062 147056
rect 183020 133929 183048 147047
rect 183006 133920 183062 133929
rect 183006 133855 183062 133864
rect 183006 120048 183062 120057
rect 183006 119983 183062 119992
rect 182916 117224 182968 117230
rect 182916 117166 182968 117172
rect 182916 101448 182968 101454
rect 182916 101390 182968 101396
rect 182928 85377 182956 101390
rect 182914 85368 182970 85377
rect 182914 85303 182970 85312
rect 182822 77888 182878 77897
rect 182822 77823 182878 77832
rect 183020 47598 183048 119983
rect 184216 110430 184244 151778
rect 184308 121650 184336 152458
rect 184386 150512 184442 150521
rect 184386 150447 184442 150456
rect 184400 133210 184428 150447
rect 185596 145081 185624 275946
rect 185768 269136 185820 269142
rect 185768 269078 185820 269084
rect 185676 252680 185728 252686
rect 185676 252622 185728 252628
rect 185688 148345 185716 252622
rect 185780 216034 185808 269078
rect 186332 240786 186360 384270
rect 187436 370530 187464 431938
rect 187516 409896 187568 409902
rect 187516 409838 187568 409844
rect 187424 370524 187476 370530
rect 187424 370466 187476 370472
rect 187424 351212 187476 351218
rect 187424 351154 187476 351160
rect 186964 299940 187016 299946
rect 186964 299882 187016 299888
rect 186976 294642 187004 299882
rect 186964 294636 187016 294642
rect 186964 294578 187016 294584
rect 187436 292602 187464 351154
rect 187528 340202 187556 409838
rect 187620 400790 187648 576846
rect 188988 484424 189040 484430
rect 188988 484366 189040 484372
rect 188344 465180 188396 465186
rect 188344 465122 188396 465128
rect 188066 452976 188122 452985
rect 188066 452911 188122 452920
rect 188080 444961 188108 452911
rect 188066 444952 188122 444961
rect 188066 444887 188122 444896
rect 188356 418130 188384 465122
rect 188436 444372 188488 444378
rect 188436 444314 188488 444320
rect 188448 434722 188476 444314
rect 188436 434716 188488 434722
rect 188436 434658 188488 434664
rect 188896 434716 188948 434722
rect 188896 434658 188948 434664
rect 188908 433294 188936 434658
rect 188896 433288 188948 433294
rect 188896 433230 188948 433236
rect 188802 432576 188858 432585
rect 188802 432511 188858 432520
rect 188344 418124 188396 418130
rect 188344 418066 188396 418072
rect 187700 416832 187752 416838
rect 187700 416774 187752 416780
rect 187712 416090 187740 416774
rect 187700 416084 187752 416090
rect 187700 416026 187752 416032
rect 188344 408536 188396 408542
rect 188344 408478 188396 408484
rect 187608 400784 187660 400790
rect 187608 400726 187660 400732
rect 187620 400246 187648 400726
rect 187608 400240 187660 400246
rect 187608 400182 187660 400188
rect 187608 385688 187660 385694
rect 187608 385630 187660 385636
rect 187620 382226 187648 385630
rect 187608 382220 187660 382226
rect 187608 382162 187660 382168
rect 187516 340196 187568 340202
rect 187516 340138 187568 340144
rect 187620 299946 187648 382162
rect 188356 378146 188384 408478
rect 188528 397520 188580 397526
rect 188528 397462 188580 397468
rect 188436 393372 188488 393378
rect 188436 393314 188488 393320
rect 188448 381546 188476 393314
rect 188540 391950 188568 397462
rect 188528 391944 188580 391950
rect 188528 391886 188580 391892
rect 188526 382392 188582 382401
rect 188526 382327 188582 382336
rect 188436 381540 188488 381546
rect 188436 381482 188488 381488
rect 188344 378140 188396 378146
rect 188344 378082 188396 378088
rect 188540 373969 188568 382327
rect 188526 373960 188582 373969
rect 188526 373895 188582 373904
rect 188816 366382 188844 432511
rect 189000 416158 189028 484366
rect 191196 463752 191248 463758
rect 191196 463694 191248 463700
rect 190368 455524 190420 455530
rect 190368 455466 190420 455472
rect 189722 452840 189778 452849
rect 189722 452775 189778 452784
rect 189736 438841 189764 452775
rect 189722 438832 189778 438841
rect 189722 438767 189778 438776
rect 188988 416152 189040 416158
rect 188988 416094 189040 416100
rect 190274 412720 190330 412729
rect 190274 412655 190330 412664
rect 190182 394768 190238 394777
rect 190182 394703 190238 394712
rect 190090 393408 190146 393417
rect 190090 393343 190146 393352
rect 190104 382945 190132 393343
rect 190090 382936 190146 382945
rect 190090 382871 190146 382880
rect 190104 382401 190132 382871
rect 190090 382392 190146 382401
rect 190090 382327 190146 382336
rect 189078 381576 189134 381585
rect 189078 381511 189134 381520
rect 189092 380866 189120 381511
rect 189080 380860 189132 380866
rect 189080 380802 189132 380808
rect 189724 380860 189776 380866
rect 189724 380802 189776 380808
rect 188896 378140 188948 378146
rect 188896 378082 188948 378088
rect 188804 366376 188856 366382
rect 188804 366318 188856 366324
rect 187700 362228 187752 362234
rect 187700 362170 187752 362176
rect 187712 361593 187740 362170
rect 187698 361584 187754 361593
rect 187698 361519 187754 361528
rect 188618 319016 188674 319025
rect 188618 318951 188674 318960
rect 188632 312497 188660 318951
rect 188618 312488 188674 312497
rect 188618 312423 188674 312432
rect 188434 312080 188490 312089
rect 188434 312015 188490 312024
rect 187698 305144 187754 305153
rect 187698 305079 187754 305088
rect 187608 299940 187660 299946
rect 187608 299882 187660 299888
rect 187712 298897 187740 305079
rect 187698 298888 187754 298897
rect 187698 298823 187754 298832
rect 187608 295384 187660 295390
rect 187608 295326 187660 295332
rect 187424 292596 187476 292602
rect 187424 292538 187476 292544
rect 186964 266416 187016 266422
rect 186964 266358 187016 266364
rect 186320 240780 186372 240786
rect 186320 240722 186372 240728
rect 185768 216028 185820 216034
rect 185768 215970 185820 215976
rect 186228 158024 186280 158030
rect 186228 157966 186280 157972
rect 185766 151192 185822 151201
rect 185766 151127 185822 151136
rect 185674 148336 185730 148345
rect 185674 148271 185730 148280
rect 185582 145072 185638 145081
rect 185582 145007 185638 145016
rect 185596 138718 185624 145007
rect 185584 138712 185636 138718
rect 185584 138654 185636 138660
rect 184388 133204 184440 133210
rect 184388 133146 184440 133152
rect 185584 126268 185636 126274
rect 185584 126210 185636 126216
rect 184296 121644 184348 121650
rect 184296 121586 184348 121592
rect 184848 121644 184900 121650
rect 184848 121586 184900 121592
rect 184860 118658 184888 121586
rect 184848 118652 184900 118658
rect 184848 118594 184900 118600
rect 184848 115252 184900 115258
rect 184848 115194 184900 115200
rect 184480 114164 184532 114170
rect 184480 114106 184532 114112
rect 184296 111852 184348 111858
rect 184296 111794 184348 111800
rect 184204 110424 184256 110430
rect 184204 110366 184256 110372
rect 184308 81433 184336 111794
rect 184388 93152 184440 93158
rect 184388 93094 184440 93100
rect 184294 81424 184350 81433
rect 184294 81359 184350 81368
rect 184204 80028 184256 80034
rect 184204 79970 184256 79976
rect 183008 47592 183060 47598
rect 183008 47534 183060 47540
rect 184216 44878 184244 79970
rect 184400 79937 184428 93094
rect 184492 80034 184520 114106
rect 184480 80028 184532 80034
rect 184480 79970 184532 79976
rect 184386 79928 184442 79937
rect 184386 79863 184442 79872
rect 184204 44872 184256 44878
rect 184204 44814 184256 44820
rect 184860 15910 184888 115194
rect 185596 89593 185624 126210
rect 185780 122913 185808 151127
rect 185766 122904 185822 122913
rect 185766 122839 185822 122848
rect 186240 114170 186268 157966
rect 186976 144129 187004 266358
rect 187620 265577 187648 295326
rect 188342 282976 188398 282985
rect 188342 282911 188398 282920
rect 187606 265568 187662 265577
rect 187606 265503 187662 265512
rect 187054 265024 187110 265033
rect 187054 264959 187110 264968
rect 187068 241505 187096 264959
rect 187148 244316 187200 244322
rect 187148 244258 187200 244264
rect 187054 241496 187110 241505
rect 187054 241431 187110 241440
rect 187160 233889 187188 244258
rect 187606 241496 187662 241505
rect 187606 241431 187662 241440
rect 187620 240825 187648 241431
rect 187698 240952 187754 240961
rect 187698 240887 187754 240896
rect 187606 240816 187662 240825
rect 187606 240751 187662 240760
rect 187146 233880 187202 233889
rect 187146 233815 187202 233824
rect 187056 216028 187108 216034
rect 187056 215970 187108 215976
rect 187068 153882 187096 215970
rect 187056 153876 187108 153882
rect 187056 153818 187108 153824
rect 186962 144120 187018 144129
rect 186962 144055 187018 144064
rect 186872 143676 186924 143682
rect 186872 143618 186924 143624
rect 186884 135969 186912 143618
rect 186870 135960 186926 135969
rect 186870 135895 186926 135904
rect 187068 120086 187096 153818
rect 187148 153332 187200 153338
rect 187148 153274 187200 153280
rect 187160 137290 187188 153274
rect 187148 137284 187200 137290
rect 187148 137226 187200 137232
rect 187148 121984 187200 121990
rect 187148 121926 187200 121932
rect 187056 120080 187108 120086
rect 187056 120022 187108 120028
rect 186964 118652 187016 118658
rect 186964 118594 187016 118600
rect 186320 117360 186372 117366
rect 186320 117302 186372 117308
rect 186332 115258 186360 117302
rect 186320 115252 186372 115258
rect 186320 115194 186372 115200
rect 186228 114164 186280 114170
rect 186228 114106 186280 114112
rect 186240 113218 186268 114106
rect 186228 113212 186280 113218
rect 186228 113154 186280 113160
rect 185768 106344 185820 106350
rect 185768 106286 185820 106292
rect 185676 99612 185728 99618
rect 185676 99554 185728 99560
rect 185582 89584 185638 89593
rect 185582 89519 185638 89528
rect 185688 66162 185716 99554
rect 185780 86902 185808 106286
rect 185860 99408 185912 99414
rect 185860 99350 185912 99356
rect 185872 93158 185900 99350
rect 185860 93152 185912 93158
rect 185860 93094 185912 93100
rect 185768 86896 185820 86902
rect 185768 86838 185820 86844
rect 185676 66156 185728 66162
rect 185676 66098 185728 66104
rect 185688 64874 185716 66098
rect 185596 64846 185716 64874
rect 185596 50386 185624 64846
rect 185584 50380 185636 50386
rect 185584 50322 185636 50328
rect 186976 40730 187004 118594
rect 187056 103556 187108 103562
rect 187056 103498 187108 103504
rect 187068 81161 187096 103498
rect 187160 97986 187188 121926
rect 187620 115462 187648 240751
rect 187712 216073 187740 240887
rect 188356 239873 188384 282911
rect 188448 269822 188476 312015
rect 188908 290358 188936 378082
rect 189078 367160 189134 367169
rect 189078 367095 189134 367104
rect 189092 366994 189120 367095
rect 189080 366988 189132 366994
rect 189080 366930 189132 366936
rect 188986 361584 189042 361593
rect 188986 361519 189042 361528
rect 188896 290352 188948 290358
rect 188896 290294 188948 290300
rect 188436 269816 188488 269822
rect 188436 269758 188488 269764
rect 188436 267844 188488 267850
rect 188436 267786 188488 267792
rect 188342 239864 188398 239873
rect 188342 239799 188398 239808
rect 188448 237969 188476 267786
rect 188526 248432 188582 248441
rect 188526 248367 188582 248376
rect 188434 237960 188490 237969
rect 188434 237895 188490 237904
rect 188540 235249 188568 248367
rect 189000 241097 189028 361519
rect 189736 272513 189764 380802
rect 190196 367169 190224 394703
rect 190288 385014 190316 412655
rect 190276 385008 190328 385014
rect 190276 384950 190328 384956
rect 190182 367160 190238 367169
rect 190182 367095 190238 367104
rect 190380 332722 190408 455466
rect 191104 451920 191156 451926
rect 191104 451862 191156 451868
rect 190458 447264 190514 447273
rect 190458 447199 190514 447208
rect 190472 444378 190500 447199
rect 190460 444372 190512 444378
rect 190460 444314 190512 444320
rect 191116 432002 191144 451862
rect 191208 446457 191236 463694
rect 191286 454336 191342 454345
rect 191286 454271 191342 454280
rect 191194 446448 191250 446457
rect 191194 446383 191250 446392
rect 191300 440910 191328 454271
rect 191472 449880 191524 449886
rect 191472 449822 191524 449828
rect 191484 449177 191512 449822
rect 191470 449168 191526 449177
rect 191470 449103 191526 449112
rect 191654 449168 191710 449177
rect 191654 449103 191710 449112
rect 191668 448594 191696 449103
rect 191656 448588 191708 448594
rect 191656 448530 191708 448536
rect 191760 447250 191788 703326
rect 202800 702642 202828 703520
rect 215208 703248 215260 703254
rect 215208 703190 215260 703196
rect 213184 702840 213236 702846
rect 213184 702782 213236 702788
rect 202788 702636 202840 702642
rect 202788 702578 202840 702584
rect 208398 470656 208454 470665
rect 208398 470591 208454 470600
rect 194598 465216 194654 465225
rect 194598 465151 194654 465160
rect 194612 460934 194640 465151
rect 195980 460964 196032 460970
rect 194612 460906 195192 460934
rect 202144 460964 202196 460970
rect 196032 460912 196112 460934
rect 195980 460906 196112 460912
rect 202144 460906 202196 460912
rect 192484 456952 192536 456958
rect 192484 456894 192536 456900
rect 191760 447222 191880 447250
rect 191746 446448 191802 446457
rect 191746 446383 191802 446392
rect 191760 445806 191788 446383
rect 191748 445800 191800 445806
rect 191748 445742 191800 445748
rect 191746 445088 191802 445097
rect 191746 445023 191802 445032
rect 191760 444446 191788 445023
rect 191748 444440 191800 444446
rect 191748 444382 191800 444388
rect 191288 440904 191340 440910
rect 191288 440846 191340 440852
rect 191196 440292 191248 440298
rect 191196 440234 191248 440240
rect 191104 431996 191156 432002
rect 191104 431938 191156 431944
rect 191208 429593 191236 440234
rect 191746 438016 191802 438025
rect 191746 437951 191802 437960
rect 191760 437510 191788 437951
rect 191748 437504 191800 437510
rect 191748 437446 191800 437452
rect 191748 435396 191800 435402
rect 191748 435338 191800 435344
rect 191760 435305 191788 435338
rect 191746 435296 191802 435305
rect 191746 435231 191802 435240
rect 191748 434716 191800 434722
rect 191748 434658 191800 434664
rect 191654 433664 191710 433673
rect 191654 433599 191710 433608
rect 191668 433362 191696 433599
rect 191656 433356 191708 433362
rect 191656 433298 191708 433304
rect 191194 429584 191250 429593
rect 191194 429519 191250 429528
rect 191470 429584 191526 429593
rect 191470 429519 191526 429528
rect 191010 425504 191066 425513
rect 191010 425439 191066 425448
rect 191024 425134 191052 425439
rect 191012 425128 191064 425134
rect 191012 425070 191064 425076
rect 190828 422952 190880 422958
rect 190828 422894 190880 422900
rect 190840 422521 190868 422894
rect 190826 422512 190882 422521
rect 190826 422447 190882 422456
rect 191012 416152 191064 416158
rect 191012 416094 191064 416100
rect 191024 415449 191052 416094
rect 191010 415440 191066 415449
rect 191010 415375 191066 415384
rect 191484 412634 191512 429519
rect 191564 429140 191616 429146
rect 191564 429082 191616 429088
rect 191576 428233 191604 429082
rect 191562 428224 191618 428233
rect 191562 428159 191618 428168
rect 191562 426864 191618 426873
rect 191562 426799 191618 426808
rect 191576 426494 191604 426799
rect 191564 426488 191616 426494
rect 191564 426430 191616 426436
rect 191562 419792 191618 419801
rect 191562 419727 191618 419736
rect 191576 419626 191604 419727
rect 191564 419620 191616 419626
rect 191564 419562 191616 419568
rect 191562 418432 191618 418441
rect 191562 418367 191618 418376
rect 191576 418198 191604 418367
rect 191564 418192 191616 418198
rect 191564 418134 191616 418140
rect 191562 417072 191618 417081
rect 191562 417007 191618 417016
rect 191576 416838 191604 417007
rect 191564 416832 191616 416838
rect 191564 416774 191616 416780
rect 191564 414724 191616 414730
rect 191564 414666 191616 414672
rect 191576 414089 191604 414666
rect 191562 414080 191618 414089
rect 191562 414015 191618 414024
rect 191484 412606 191604 412634
rect 191472 411936 191524 411942
rect 191472 411878 191524 411884
rect 191484 411369 191512 411878
rect 191470 411360 191526 411369
rect 191470 411295 191526 411304
rect 190826 410000 190882 410009
rect 190826 409935 190882 409944
rect 190840 409902 190868 409935
rect 190828 409896 190880 409902
rect 190828 409838 190880 409844
rect 191470 407008 191526 407017
rect 191470 406943 191526 406952
rect 191484 405822 191512 406943
rect 191472 405816 191524 405822
rect 191472 405758 191524 405764
rect 191378 405648 191434 405657
rect 191378 405583 191434 405592
rect 191392 404394 191420 405583
rect 191380 404388 191432 404394
rect 191380 404330 191432 404336
rect 191470 404288 191526 404297
rect 191470 404223 191526 404232
rect 191484 403102 191512 404223
rect 191472 403096 191524 403102
rect 191472 403038 191524 403044
rect 191378 402928 191434 402937
rect 191378 402863 191434 402872
rect 190826 400208 190882 400217
rect 190826 400143 190882 400152
rect 190840 398886 190868 400143
rect 190828 398880 190880 398886
rect 190828 398822 190880 398828
rect 191102 398576 191158 398585
rect 191102 398511 191158 398520
rect 191116 397594 191144 398511
rect 191104 397588 191156 397594
rect 191104 397530 191156 397536
rect 191392 396098 191420 402863
rect 191470 401568 191526 401577
rect 191470 401503 191526 401512
rect 191484 400790 191512 401503
rect 191472 400784 191524 400790
rect 191472 400726 191524 400732
rect 191472 397452 191524 397458
rect 191472 397394 191524 397400
rect 191484 397225 191512 397394
rect 191470 397216 191526 397225
rect 191470 397151 191526 397160
rect 191196 396092 191248 396098
rect 191196 396034 191248 396040
rect 191380 396092 191432 396098
rect 191380 396034 191432 396040
rect 191010 390960 191066 390969
rect 191010 390895 191066 390904
rect 191024 390658 191052 390895
rect 191012 390652 191064 390658
rect 191012 390594 191064 390600
rect 189908 332716 189960 332722
rect 189908 332658 189960 332664
rect 190368 332716 190420 332722
rect 190368 332658 190420 332664
rect 189816 303748 189868 303754
rect 189816 303690 189868 303696
rect 189722 272504 189778 272513
rect 189722 272439 189778 272448
rect 189722 245848 189778 245857
rect 189722 245783 189778 245792
rect 188986 241088 189042 241097
rect 188986 241023 189042 241032
rect 188986 240136 189042 240145
rect 188986 240071 189042 240080
rect 188526 235240 188582 235249
rect 188526 235175 188582 235184
rect 187698 216064 187754 216073
rect 187698 215999 187754 216008
rect 187712 215393 187740 215999
rect 187698 215384 187754 215393
rect 187698 215319 187754 215328
rect 188342 215384 188398 215393
rect 188342 215319 188398 215328
rect 188356 201482 188384 215319
rect 188344 201476 188396 201482
rect 188344 201418 188396 201424
rect 188896 201476 188948 201482
rect 188896 201418 188948 201424
rect 188908 201385 188936 201418
rect 188894 201376 188950 201385
rect 188894 201311 188950 201320
rect 189000 193866 189028 240071
rect 188988 193860 189040 193866
rect 188988 193802 189040 193808
rect 189736 184210 189764 245783
rect 189828 232529 189856 303690
rect 189920 279478 189948 332658
rect 189998 306504 190054 306513
rect 189998 306439 190054 306448
rect 190012 294545 190040 306439
rect 191102 301608 191158 301617
rect 191102 301543 191158 301552
rect 191116 301073 191144 301543
rect 191102 301064 191158 301073
rect 191102 300999 191104 301008
rect 191156 300999 191158 301008
rect 191104 300970 191156 300976
rect 191116 300939 191144 300970
rect 190644 299464 190696 299470
rect 190644 299406 190696 299412
rect 190656 299033 190684 299406
rect 190642 299024 190698 299033
rect 190642 298959 190698 298968
rect 189998 294536 190054 294545
rect 189998 294471 190054 294480
rect 190644 288312 190696 288318
rect 190644 288254 190696 288260
rect 190656 287473 190684 288254
rect 190642 287464 190698 287473
rect 190642 287399 190698 287408
rect 191010 286512 191066 286521
rect 191010 286447 191066 286456
rect 191024 285802 191052 286447
rect 191012 285796 191064 285802
rect 191012 285738 191064 285744
rect 191102 284336 191158 284345
rect 191102 284271 191158 284280
rect 189908 279472 189960 279478
rect 189908 279414 189960 279420
rect 190460 277296 190512 277302
rect 190460 277238 190512 277244
rect 189908 247716 189960 247722
rect 189908 247658 189960 247664
rect 189814 232520 189870 232529
rect 189814 232455 189870 232464
rect 189920 224777 189948 247658
rect 189998 242992 190054 243001
rect 189998 242927 190054 242936
rect 190012 236609 190040 242927
rect 189998 236600 190054 236609
rect 189998 236535 190054 236544
rect 189906 224768 189962 224777
rect 189906 224703 189962 224712
rect 190368 191140 190420 191146
rect 190368 191082 190420 191088
rect 189724 184204 189776 184210
rect 189724 184146 189776 184152
rect 189724 170400 189776 170406
rect 189724 170342 189776 170348
rect 189736 162897 189764 170342
rect 189722 162888 189778 162897
rect 189722 162823 189778 162832
rect 188894 158808 188950 158817
rect 188894 158743 188950 158752
rect 187698 147928 187754 147937
rect 187698 147863 187754 147872
rect 187712 145625 187740 147863
rect 188434 146432 188490 146441
rect 188434 146367 188490 146376
rect 187698 145616 187754 145625
rect 187698 145551 187754 145560
rect 188344 145580 188396 145586
rect 188344 145522 188396 145528
rect 187700 120148 187752 120154
rect 187700 120090 187752 120096
rect 187712 117298 187740 120090
rect 187700 117292 187752 117298
rect 187700 117234 187752 117240
rect 187608 115456 187660 115462
rect 187608 115398 187660 115404
rect 187240 102808 187292 102814
rect 187240 102750 187292 102756
rect 187148 97980 187200 97986
rect 187148 97922 187200 97928
rect 187252 82822 187280 102750
rect 188356 100706 188384 145522
rect 188448 130422 188476 146367
rect 188436 130416 188488 130422
rect 188436 130358 188488 130364
rect 188908 128489 188936 158743
rect 189078 142216 189134 142225
rect 189078 142151 189134 142160
rect 188988 140480 189040 140486
rect 188988 140422 189040 140428
rect 188894 128480 188950 128489
rect 188894 128415 188950 128424
rect 188436 116068 188488 116074
rect 188436 116010 188488 116016
rect 188448 111110 188476 116010
rect 188436 111104 188488 111110
rect 188436 111046 188488 111052
rect 188896 104916 188948 104922
rect 188896 104858 188948 104864
rect 188528 102196 188580 102202
rect 188528 102138 188580 102144
rect 188344 100700 188396 100706
rect 188344 100642 188396 100648
rect 188436 98184 188488 98190
rect 188436 98126 188488 98132
rect 187700 98048 187752 98054
rect 187700 97990 187752 97996
rect 187712 97306 187740 97990
rect 187700 97300 187752 97306
rect 187700 97242 187752 97248
rect 187608 95328 187660 95334
rect 187608 95270 187660 95276
rect 187620 87961 187648 95270
rect 187606 87952 187662 87961
rect 187606 87887 187662 87896
rect 188342 85504 188398 85513
rect 188342 85439 188398 85448
rect 187240 82816 187292 82822
rect 187240 82758 187292 82764
rect 187054 81152 187110 81161
rect 187054 81087 187110 81096
rect 187068 58682 187096 81087
rect 187698 71768 187754 71777
rect 187698 71703 187700 71712
rect 187752 71703 187754 71712
rect 187700 71674 187752 71680
rect 187056 58676 187108 58682
rect 187056 58618 187108 58624
rect 188356 46918 188384 85439
rect 188448 68950 188476 98126
rect 188540 93129 188568 102138
rect 188526 93120 188582 93129
rect 188526 93055 188582 93064
rect 188908 71777 188936 104858
rect 189000 102270 189028 140422
rect 189092 139369 189120 142151
rect 189078 139360 189134 139369
rect 189078 139295 189134 139304
rect 189736 132569 189764 162823
rect 189908 157412 189960 157418
rect 189908 157354 189960 157360
rect 189814 135144 189870 135153
rect 189814 135079 189870 135088
rect 189722 132560 189778 132569
rect 189722 132495 189778 132504
rect 189080 128716 189132 128722
rect 189080 128658 189132 128664
rect 189092 123486 189120 128658
rect 189722 124264 189778 124273
rect 189722 124199 189778 124208
rect 189080 123480 189132 123486
rect 189080 123422 189132 123428
rect 189736 120018 189764 124199
rect 189724 120012 189776 120018
rect 189724 119954 189776 119960
rect 188988 102264 189040 102270
rect 188988 102206 189040 102212
rect 188894 71768 188950 71777
rect 188894 71703 188950 71712
rect 188436 68944 188488 68950
rect 188436 68886 188488 68892
rect 189736 53106 189764 119954
rect 189828 92313 189856 135079
rect 189920 133929 189948 157354
rect 190380 138553 190408 191082
rect 190472 165646 190500 277238
rect 190826 270056 190882 270065
rect 190826 269991 190882 270000
rect 190840 269142 190868 269991
rect 190828 269136 190880 269142
rect 190828 269078 190880 269084
rect 190826 266112 190882 266121
rect 190826 266047 190882 266056
rect 190840 264994 190868 266047
rect 190828 264988 190880 264994
rect 190828 264930 190880 264936
rect 191010 263256 191066 263265
rect 191010 263191 191066 263200
rect 191024 262342 191052 263191
rect 191012 262336 191064 262342
rect 191012 262278 191064 262284
rect 190644 258120 190696 258126
rect 190696 258068 190776 258074
rect 190644 258062 190776 258068
rect 190656 258058 190776 258062
rect 190656 258052 190788 258058
rect 190656 258046 190736 258052
rect 190736 257994 190788 258000
rect 190826 256456 190882 256465
rect 190826 256391 190882 256400
rect 190840 255338 190868 256391
rect 191010 255504 191066 255513
rect 191010 255439 191066 255448
rect 191024 255406 191052 255439
rect 191012 255400 191064 255406
rect 191012 255342 191064 255348
rect 190828 255332 190880 255338
rect 190828 255274 190880 255280
rect 190642 250744 190698 250753
rect 190642 250679 190698 250688
rect 190656 249830 190684 250679
rect 190644 249824 190696 249830
rect 190644 249766 190696 249772
rect 190826 249656 190882 249665
rect 190826 249591 190882 249600
rect 190840 248538 190868 249591
rect 190828 248532 190880 248538
rect 190828 248474 190880 248480
rect 190460 165640 190512 165646
rect 190460 165582 190512 165588
rect 190366 138544 190422 138553
rect 190366 138479 190422 138488
rect 190092 137828 190144 137834
rect 190092 137770 190144 137776
rect 189906 133920 189962 133929
rect 189906 133855 189962 133864
rect 190104 125798 190132 137770
rect 191116 132462 191144 284271
rect 191208 274825 191236 396034
rect 191472 391944 191524 391950
rect 191472 391886 191524 391892
rect 191484 391785 191512 391886
rect 191470 391776 191526 391785
rect 191470 391711 191526 391720
rect 191472 301504 191524 301510
rect 191472 301446 191524 301452
rect 191484 298081 191512 301446
rect 191470 298072 191526 298081
rect 191470 298007 191526 298016
rect 191576 291281 191604 412606
rect 191562 291272 191618 291281
rect 191562 291207 191618 291216
rect 191564 289808 191616 289814
rect 191564 289750 191616 289756
rect 191576 289377 191604 289750
rect 191562 289368 191618 289377
rect 191562 289303 191618 289312
rect 191668 285569 191696 433298
rect 191760 301510 191788 434658
rect 191852 425513 191880 447222
rect 192496 446418 192524 456894
rect 192576 455456 192628 455462
rect 192576 455398 192628 455404
rect 192588 447846 192616 455398
rect 193404 454164 193456 454170
rect 193404 454106 193456 454112
rect 193310 451480 193366 451489
rect 193310 451415 193366 451424
rect 193324 447953 193352 451415
rect 193416 449206 193444 454106
rect 194598 450256 194654 450265
rect 195164 450242 195192 460906
rect 196084 450242 196112 460906
rect 197084 458312 197136 458318
rect 197082 458280 197084 458289
rect 197136 458280 197138 458289
rect 197082 458215 197138 458224
rect 197360 456884 197412 456890
rect 197360 456826 197412 456832
rect 197372 450242 197400 456826
rect 197910 454200 197966 454209
rect 197910 454135 197966 454144
rect 197924 450242 197952 454135
rect 202156 452985 202184 460906
rect 207478 457056 207534 457065
rect 207478 456991 207534 457000
rect 204444 456816 204496 456822
rect 204444 456758 204496 456764
rect 202878 455696 202934 455705
rect 202878 455631 202934 455640
rect 202142 452976 202198 452985
rect 202142 452911 202198 452920
rect 200396 452736 200448 452742
rect 200396 452678 200448 452684
rect 201592 452736 201644 452742
rect 201592 452678 201644 452684
rect 199292 451308 199344 451314
rect 199292 451250 199344 451256
rect 194654 450214 194718 450242
rect 195164 450214 195638 450242
rect 196084 450214 196558 450242
rect 197372 450214 197478 450242
rect 197924 450214 198398 450242
rect 199304 450228 199332 451250
rect 200408 450228 200436 452678
rect 201316 452668 201368 452674
rect 201316 452610 201368 452616
rect 201328 450228 201356 452610
rect 201604 450401 201632 452678
rect 201590 450392 201646 450401
rect 201590 450327 201646 450336
rect 202156 450242 202184 452911
rect 202788 452668 202840 452674
rect 202788 452610 202840 452616
rect 202800 451926 202828 452610
rect 202788 451920 202840 451926
rect 202788 451862 202840 451868
rect 202892 450242 202920 455631
rect 204456 451897 204484 456758
rect 204536 455524 204588 455530
rect 204536 455466 204588 455472
rect 204442 451888 204498 451897
rect 204442 451823 204498 451832
rect 204076 451308 204128 451314
rect 204076 451250 204128 451256
rect 202156 450214 202262 450242
rect 202892 450214 203182 450242
rect 204088 450228 204116 451250
rect 204548 450242 204576 455466
rect 205916 452736 205968 452742
rect 205916 452678 205968 452684
rect 204548 450214 205022 450242
rect 205928 450228 205956 452678
rect 207018 451480 207074 451489
rect 207018 451415 207074 451424
rect 207032 450228 207060 451415
rect 207492 450242 207520 456991
rect 208412 450242 208440 470591
rect 211160 466540 211212 466546
rect 211160 466482 211212 466488
rect 210698 452840 210754 452849
rect 210698 452775 210754 452784
rect 209780 452668 209832 452674
rect 209780 452610 209832 452616
rect 207492 450214 207966 450242
rect 208412 450214 208886 450242
rect 209792 450228 209820 452610
rect 210712 451489 210740 452775
rect 210698 451480 210754 451489
rect 210698 451415 210754 451424
rect 210712 450228 210740 451415
rect 211172 450242 211200 466482
rect 213196 462233 213224 702782
rect 215220 465225 215248 703190
rect 215944 702636 215996 702642
rect 215944 702578 215996 702584
rect 213918 465216 213974 465225
rect 213918 465151 213974 465160
rect 215206 465216 215262 465225
rect 215206 465151 215262 465160
rect 212538 462224 212594 462233
rect 212538 462159 212594 462168
rect 213182 462224 213238 462233
rect 213182 462159 213238 462168
rect 212552 461145 212580 462159
rect 212538 461136 212594 461145
rect 212538 461071 212594 461080
rect 212552 450242 212580 461071
rect 213932 460934 213960 465151
rect 215956 465089 215984 702578
rect 218992 700330 219020 703520
rect 220084 703044 220136 703050
rect 220084 702986 220136 702992
rect 218980 700324 219032 700330
rect 218980 700266 219032 700272
rect 218060 478916 218112 478922
rect 218060 478858 218112 478864
rect 215298 465080 215354 465089
rect 215298 465015 215354 465024
rect 215942 465080 215998 465089
rect 215942 465015 215998 465024
rect 215312 463729 215340 465015
rect 215298 463720 215354 463729
rect 215298 463655 215354 463664
rect 215312 460934 215340 463655
rect 213932 460906 214236 460934
rect 215312 460906 216076 460934
rect 213184 455456 213236 455462
rect 213184 455398 213236 455404
rect 213196 450242 213224 455398
rect 211172 450214 211646 450242
rect 212552 450214 212750 450242
rect 213196 450214 213670 450242
rect 194598 450191 194654 450200
rect 214208 450022 214236 460906
rect 215390 456920 215446 456929
rect 215390 456855 215446 456864
rect 215404 450242 215432 456855
rect 216048 450242 216076 460906
rect 216678 458688 216734 458697
rect 216678 458623 216734 458632
rect 216692 458425 216720 458623
rect 216678 458416 216734 458425
rect 216678 458351 216734 458360
rect 216692 451274 216720 458351
rect 216692 451246 216904 451274
rect 216876 450242 216904 451246
rect 218072 450242 218100 478858
rect 220096 458697 220124 702986
rect 235184 702914 235212 703520
rect 240784 703180 240836 703186
rect 240784 703122 240836 703128
rect 235172 702908 235224 702914
rect 235172 702850 235224 702856
rect 240796 487830 240824 703122
rect 249708 703112 249760 703118
rect 249708 703054 249760 703060
rect 241520 700324 241572 700330
rect 241520 700266 241572 700272
rect 240784 487824 240836 487830
rect 240784 487766 240836 487772
rect 227812 473408 227864 473414
rect 227812 473350 227864 473356
rect 225604 462460 225656 462466
rect 225604 462402 225656 462408
rect 223580 462392 223632 462398
rect 223580 462334 223632 462340
rect 223592 460934 223620 462334
rect 223592 460906 223712 460934
rect 220082 458688 220138 458697
rect 220082 458623 220138 458632
rect 220818 458416 220874 458425
rect 220818 458351 220874 458360
rect 218888 456952 218940 456958
rect 218888 456894 218940 456900
rect 218900 450242 218928 456894
rect 219806 455832 219862 455841
rect 219806 455767 219862 455776
rect 219820 450242 219848 455767
rect 215404 450214 215510 450242
rect 216048 450214 216430 450242
rect 216876 450214 217350 450242
rect 218072 450214 218652 450242
rect 218900 450214 219374 450242
rect 219820 450214 220294 450242
rect 218624 450022 218652 450214
rect 214196 450016 214248 450022
rect 218612 450016 218664 450022
rect 214248 449964 214590 449970
rect 214196 449958 214590 449964
rect 220832 449993 220860 458351
rect 222566 454336 222622 454345
rect 222566 454271 222622 454280
rect 222106 452976 222162 452985
rect 222106 452911 222162 452920
rect 222120 450228 222148 452911
rect 222580 450242 222608 454271
rect 223684 450242 223712 460906
rect 224958 455696 225014 455705
rect 224958 455631 225014 455640
rect 224972 450242 225000 455631
rect 225616 452849 225644 462402
rect 227720 458312 227772 458318
rect 227720 458254 227772 458260
rect 226432 456884 226484 456890
rect 226432 456826 226484 456832
rect 225970 453112 226026 453121
rect 225970 453047 226026 453056
rect 225602 452840 225658 452849
rect 225602 452775 225658 452784
rect 222580 450214 223054 450242
rect 223684 450214 224158 450242
rect 224972 450214 225078 450242
rect 225984 450228 226012 453047
rect 226444 450242 226472 456826
rect 227732 452674 227760 458254
rect 227720 452668 227772 452674
rect 227720 452610 227772 452616
rect 227824 450242 227852 473350
rect 240140 465112 240192 465118
rect 240140 465054 240192 465060
rect 231124 463752 231176 463758
rect 231124 463694 231176 463700
rect 231136 456929 231164 463694
rect 233240 461032 233292 461038
rect 233240 460974 233292 460980
rect 233252 460934 233280 460974
rect 240152 460934 240180 465054
rect 233252 460906 234108 460934
rect 240152 460906 240640 460934
rect 233332 459672 233384 459678
rect 233332 459614 233384 459620
rect 230478 456920 230534 456929
rect 230478 456855 230534 456864
rect 231122 456920 231178 456929
rect 231122 456855 231178 456864
rect 228730 452840 228786 452849
rect 228730 452775 228786 452784
rect 228086 450256 228142 450265
rect 226444 450214 226918 450242
rect 227824 450228 228086 450242
rect 227838 450214 228086 450228
rect 228744 450228 228772 452775
rect 229652 452668 229704 452674
rect 229652 452610 229704 452616
rect 229664 450228 229692 452610
rect 230492 450242 230520 456855
rect 231676 453416 231728 453422
rect 231676 453358 231728 453364
rect 230492 450214 230782 450242
rect 231688 450228 231716 453358
rect 232596 452804 232648 452810
rect 232596 452746 232648 452752
rect 228086 450191 228142 450200
rect 218612 449958 218664 449964
rect 220818 449984 220874 449993
rect 214208 449942 214590 449958
rect 232608 449970 232636 452746
rect 233344 450242 233372 459614
rect 234080 450242 234108 460906
rect 236000 455524 236052 455530
rect 236000 455466 236052 455472
rect 235354 451616 235410 451625
rect 235354 451551 235410 451560
rect 233344 450214 233542 450242
rect 234080 450214 234462 450242
rect 235368 450228 235396 451551
rect 236012 450242 236040 455466
rect 237380 455456 237432 455462
rect 237380 455398 237432 455404
rect 237392 453422 237420 455398
rect 237840 454164 237892 454170
rect 237840 454106 237892 454112
rect 237380 453416 237432 453422
rect 237380 453358 237432 453364
rect 237852 450242 237880 454106
rect 239220 454028 239272 454034
rect 239220 453970 239272 453976
rect 236012 450214 236486 450242
rect 237852 450214 238326 450242
rect 239232 450228 239260 453970
rect 240140 453484 240192 453490
rect 240140 453426 240192 453432
rect 240152 452742 240180 453426
rect 240140 452736 240192 452742
rect 240140 452678 240192 452684
rect 240152 450228 240180 452678
rect 240612 450242 240640 460906
rect 240796 454170 240824 487766
rect 241532 481642 241560 700266
rect 241520 481636 241572 481642
rect 241520 481578 241572 481584
rect 242164 481636 242216 481642
rect 242164 481578 242216 481584
rect 242176 480962 242204 481578
rect 242164 480956 242216 480962
rect 242164 480898 242216 480904
rect 241520 476128 241572 476134
rect 241520 476070 241572 476076
rect 240876 466472 240928 466478
rect 240876 466414 240928 466420
rect 240784 454164 240836 454170
rect 240784 454106 240836 454112
rect 240796 454034 240824 454106
rect 240784 454028 240836 454034
rect 240784 453970 240836 453976
rect 240888 453490 240916 466414
rect 240876 453484 240928 453490
rect 240876 453426 240928 453432
rect 240612 450214 241086 450242
rect 233146 450120 233202 450129
rect 241532 450106 241560 476070
rect 242176 455433 242204 480898
rect 245660 467900 245712 467906
rect 245660 467842 245712 467848
rect 245672 460934 245700 467842
rect 245672 460906 246436 460934
rect 242162 455424 242218 455433
rect 242162 455359 242218 455368
rect 243542 455424 243598 455433
rect 243542 455359 243598 455368
rect 243556 454209 243584 455359
rect 243542 454200 243598 454209
rect 243542 454135 243598 454144
rect 243556 450242 243584 454135
rect 245752 454096 245804 454102
rect 245752 454038 245804 454044
rect 245764 450242 245792 454038
rect 246026 452976 246082 452985
rect 246026 452911 246082 452920
rect 243556 450214 244030 450242
rect 245764 450214 245870 450242
rect 242438 450120 242494 450129
rect 241532 450078 242438 450106
rect 233146 450055 233202 450064
rect 242438 450055 242494 450064
rect 220874 449942 221214 449970
rect 232240 449956 232636 449970
rect 232240 449954 232622 449956
rect 233160 449954 233188 450055
rect 237654 449984 237710 449993
rect 232228 449948 232622 449954
rect 220818 449919 220874 449928
rect 232280 449942 232622 449948
rect 233148 449948 233200 449954
rect 232228 449890 232280 449896
rect 237406 449942 237654 449970
rect 244568 449954 244950 449970
rect 237654 449919 237710 449928
rect 244556 449948 244950 449954
rect 233148 449890 233200 449896
rect 244608 449942 244950 449948
rect 244556 449890 244608 449896
rect 246040 449886 246068 452911
rect 246408 450242 246436 460906
rect 247408 456816 247460 456822
rect 247408 456758 247460 456764
rect 247420 450242 247448 456758
rect 248788 451376 248840 451382
rect 249720 451353 249748 703054
rect 267660 703050 267688 703520
rect 283852 703390 283880 703520
rect 283840 703384 283892 703390
rect 283840 703326 283892 703332
rect 273904 703316 273956 703322
rect 273904 703258 273956 703264
rect 267648 703044 267700 703050
rect 267648 702986 267700 702992
rect 271144 702908 271196 702914
rect 271144 702850 271196 702856
rect 255412 474768 255464 474774
rect 255412 474710 255464 474716
rect 253940 469328 253992 469334
rect 253940 469270 253992 469276
rect 252560 469260 252612 469266
rect 252560 469202 252612 469208
rect 252572 460934 252600 469202
rect 252572 460906 252968 460934
rect 251546 452976 251602 452985
rect 251546 452911 251602 452920
rect 248788 451318 248840 451324
rect 249706 451344 249762 451353
rect 246408 450214 246790 450242
rect 247420 450214 247894 450242
rect 248800 450228 248828 451318
rect 249706 451279 249762 451288
rect 249720 450228 249748 451279
rect 250258 449984 250314 449993
rect 250314 449942 250654 449970
rect 250258 449919 250314 449928
rect 246028 449880 246080 449886
rect 246028 449822 246080 449828
rect 193494 449712 193550 449721
rect 242990 449712 243046 449721
rect 193550 449670 193614 449698
rect 193494 449647 193550 449656
rect 251560 449698 251588 452911
rect 252466 452704 252522 452713
rect 252466 452639 252522 452648
rect 252480 450228 252508 452639
rect 252940 450242 252968 460906
rect 253846 452840 253902 452849
rect 253846 452775 253902 452784
rect 252940 450214 253414 450242
rect 251824 449744 251876 449750
rect 243046 449670 243110 449698
rect 251560 449692 251824 449698
rect 251560 449686 251876 449692
rect 251560 449684 251864 449686
rect 251574 449670 251864 449684
rect 242990 449647 243046 449656
rect 193404 449200 193456 449206
rect 193404 449142 193456 449148
rect 193310 447944 193366 447953
rect 193310 447879 193366 447888
rect 192576 447840 192628 447846
rect 192576 447782 192628 447788
rect 253860 446418 253888 452775
rect 192484 446412 192536 446418
rect 192484 446354 192536 446360
rect 253848 446412 253900 446418
rect 253848 446354 253900 446360
rect 193126 442096 193182 442105
rect 193126 442031 193182 442040
rect 192942 436656 192998 436665
rect 192942 436591 192998 436600
rect 191838 425504 191894 425513
rect 191838 425439 191894 425448
rect 192850 423872 192906 423881
rect 192850 423807 192906 423816
rect 192864 385665 192892 423807
rect 192956 387025 192984 436591
rect 193034 408640 193090 408649
rect 193034 408575 193090 408584
rect 192942 387016 192998 387025
rect 192942 386951 192998 386960
rect 192850 385656 192906 385665
rect 192850 385591 192906 385600
rect 193048 351286 193076 408575
rect 193140 363633 193168 442031
rect 253952 440473 253980 469270
rect 254122 459640 254178 459649
rect 254122 459575 254178 459584
rect 254032 451376 254084 451382
rect 254032 451318 254084 451324
rect 253938 440464 253994 440473
rect 253938 440399 253994 440408
rect 253938 432032 253994 432041
rect 253938 431967 253994 431976
rect 193404 393440 193456 393446
rect 193404 393382 193456 393388
rect 193310 391232 193366 391241
rect 193310 391167 193366 391176
rect 193324 383654 193352 391167
rect 193416 391082 193444 393382
rect 253662 392864 253718 392873
rect 253662 392799 253718 392808
rect 253572 391604 253624 391610
rect 253572 391546 253624 391552
rect 193416 391054 193614 391082
rect 250536 390992 250588 390998
rect 250536 390934 250588 390940
rect 195978 390824 196034 390833
rect 196034 390782 196374 390810
rect 195978 390759 196034 390768
rect 203536 390658 203918 390674
rect 203524 390652 203918 390658
rect 203576 390646 203918 390652
rect 203524 390594 203576 390600
rect 194140 390584 194192 390590
rect 194192 390532 194534 390538
rect 194140 390526 194534 390532
rect 194152 390510 194534 390526
rect 194612 390374 195454 390402
rect 196544 390374 197294 390402
rect 197372 390374 198214 390402
rect 198752 390374 199134 390402
rect 200132 390374 200238 390402
rect 193324 383626 193536 383654
rect 193126 363624 193182 363633
rect 193126 363559 193182 363568
rect 193508 353977 193536 383626
rect 194612 361554 194640 390374
rect 196544 373994 196572 390374
rect 197372 383897 197400 390374
rect 197358 383888 197414 383897
rect 197358 383823 197414 383832
rect 197372 381721 197400 383823
rect 197358 381712 197414 381721
rect 197358 381647 197414 381656
rect 195992 373966 196572 373994
rect 195888 363656 195940 363662
rect 195888 363598 195940 363604
rect 195900 362846 195928 363598
rect 195888 362840 195940 362846
rect 195888 362782 195940 362788
rect 194600 361548 194652 361554
rect 194600 361490 194652 361496
rect 195992 356017 196020 373966
rect 198004 370524 198056 370530
rect 198004 370466 198056 370472
rect 195978 356008 196034 356017
rect 195978 355943 196034 355952
rect 196622 356008 196678 356017
rect 196622 355943 196678 355952
rect 196636 355337 196664 355943
rect 196622 355328 196678 355337
rect 196622 355263 196678 355272
rect 193494 353968 193550 353977
rect 193494 353903 193550 353912
rect 193036 351280 193088 351286
rect 193036 351222 193088 351228
rect 192852 347064 192904 347070
rect 192852 347006 192904 347012
rect 192484 313404 192536 313410
rect 192484 313346 192536 313352
rect 192496 302938 192524 313346
rect 192574 306640 192630 306649
rect 192574 306575 192630 306584
rect 192484 302932 192536 302938
rect 192484 302874 192536 302880
rect 191748 301504 191800 301510
rect 191748 301446 191800 301452
rect 191748 301368 191800 301374
rect 191748 301310 191800 301316
rect 191760 300937 191788 301310
rect 191746 300928 191802 300937
rect 191746 300863 191802 300872
rect 192208 300824 192260 300830
rect 192208 300766 192260 300772
rect 191746 299976 191802 299985
rect 191746 299911 191748 299920
rect 191800 299911 191802 299920
rect 191748 299882 191800 299888
rect 192220 299577 192248 300766
rect 192206 299568 192262 299577
rect 192206 299503 192262 299512
rect 192588 298217 192616 306575
rect 192760 302320 192812 302326
rect 192758 302288 192760 302297
rect 192812 302288 192814 302297
rect 192758 302223 192814 302232
rect 192574 298208 192630 298217
rect 192574 298143 192630 298152
rect 191746 297120 191802 297129
rect 191746 297055 191802 297064
rect 191760 296750 191788 297055
rect 191748 296744 191800 296750
rect 191748 296686 191800 296692
rect 192482 295216 192538 295225
rect 192482 295151 192538 295160
rect 191746 294264 191802 294273
rect 191746 294199 191802 294208
rect 191760 294166 191788 294199
rect 191748 294160 191800 294166
rect 191748 294102 191800 294108
rect 191746 292632 191802 292641
rect 191746 292567 191748 292576
rect 191800 292567 191802 292576
rect 191748 292538 191800 292544
rect 191746 292224 191802 292233
rect 191746 292159 191802 292168
rect 191760 291854 191788 292159
rect 191748 291848 191800 291854
rect 191748 291790 191800 291796
rect 191748 290352 191800 290358
rect 191746 290320 191748 290329
rect 191800 290320 191802 290329
rect 191746 290255 191802 290264
rect 191746 288416 191802 288425
rect 191746 288351 191748 288360
rect 191800 288351 191802 288360
rect 191748 288322 191800 288328
rect 191654 285560 191710 285569
rect 191654 285495 191710 285504
rect 191668 284345 191696 285495
rect 191748 284980 191800 284986
rect 191748 284922 191800 284928
rect 191760 284481 191788 284922
rect 191746 284472 191802 284481
rect 191746 284407 191802 284416
rect 191654 284336 191710 284345
rect 191654 284271 191710 284280
rect 191564 282872 191616 282878
rect 191564 282814 191616 282820
rect 191576 282577 191604 282814
rect 191562 282568 191618 282577
rect 191562 282503 191618 282512
rect 191746 281616 191802 281625
rect 191746 281551 191748 281560
rect 191800 281551 191802 281560
rect 191748 281522 191800 281528
rect 191286 280664 191342 280673
rect 191286 280599 191342 280608
rect 191300 277302 191328 280599
rect 191564 280152 191616 280158
rect 191564 280094 191616 280100
rect 191576 279721 191604 280094
rect 191562 279712 191618 279721
rect 191562 279647 191618 279656
rect 191288 277296 191340 277302
rect 191288 277238 191340 277244
rect 191194 274816 191250 274825
rect 191194 274751 191250 274760
rect 191562 274816 191618 274825
rect 191562 274751 191618 274760
rect 191470 269104 191526 269113
rect 191470 269039 191526 269048
rect 191484 267782 191512 269039
rect 191472 267776 191524 267782
rect 191472 267718 191524 267724
rect 191576 267734 191604 274751
rect 191654 272912 191710 272921
rect 191654 272847 191710 272856
rect 191668 271930 191696 272847
rect 191748 271992 191800 271998
rect 191746 271960 191748 271969
rect 191800 271960 191802 271969
rect 191656 271924 191708 271930
rect 191746 271895 191802 271904
rect 191656 271866 191708 271872
rect 191746 271008 191802 271017
rect 191746 270943 191802 270952
rect 191760 270570 191788 270943
rect 191748 270564 191800 270570
rect 191748 270506 191800 270512
rect 191746 268152 191802 268161
rect 191746 268087 191802 268096
rect 191760 267850 191788 268087
rect 191748 267844 191800 267850
rect 191748 267786 191800 267792
rect 191576 267706 191696 267734
rect 191562 261352 191618 261361
rect 191562 261287 191618 261296
rect 191576 260914 191604 261287
rect 191564 260908 191616 260914
rect 191564 260850 191616 260856
rect 191668 258074 191696 267706
rect 191746 267064 191802 267073
rect 191746 266999 191802 267008
rect 191760 266422 191788 266999
rect 191748 266416 191800 266422
rect 191748 266358 191800 266364
rect 191746 264208 191802 264217
rect 191746 264143 191802 264152
rect 191760 263702 191788 264143
rect 191748 263696 191800 263702
rect 191748 263638 191800 263644
rect 191746 262304 191802 262313
rect 191746 262239 191748 262248
rect 191800 262239 191802 262248
rect 191748 262210 191800 262216
rect 191746 260400 191802 260409
rect 191746 260335 191802 260344
rect 191760 259486 191788 260335
rect 191748 259480 191800 259486
rect 191748 259422 191800 259428
rect 191746 258360 191802 258369
rect 191746 258295 191802 258304
rect 191760 258194 191788 258295
rect 191748 258188 191800 258194
rect 191748 258130 191800 258136
rect 191668 258046 191788 258074
rect 191654 257408 191710 257417
rect 191654 257343 191710 257352
rect 191668 256766 191696 257343
rect 191656 256760 191708 256766
rect 191656 256702 191708 256708
rect 191654 254552 191710 254561
rect 191654 254487 191710 254496
rect 191668 253978 191696 254487
rect 191656 253972 191708 253978
rect 191656 253914 191708 253920
rect 191562 253600 191618 253609
rect 191562 253535 191618 253544
rect 191576 252618 191604 253535
rect 191656 252680 191708 252686
rect 191654 252648 191656 252657
rect 191708 252648 191710 252657
rect 191564 252612 191616 252618
rect 191654 252583 191710 252592
rect 191564 252554 191616 252560
rect 191654 247752 191710 247761
rect 191654 247687 191710 247696
rect 191668 247110 191696 247687
rect 191656 247104 191708 247110
rect 191656 247046 191708 247052
rect 191654 244896 191710 244905
rect 191654 244831 191710 244840
rect 191668 244322 191696 244831
rect 191656 244316 191708 244322
rect 191656 244258 191708 244264
rect 191654 243944 191710 243953
rect 191654 243879 191710 243888
rect 191668 242962 191696 243879
rect 191656 242956 191708 242962
rect 191656 242898 191708 242904
rect 191196 165640 191248 165646
rect 191196 165582 191248 165588
rect 190460 132456 190512 132462
rect 190460 132398 190512 132404
rect 191104 132456 191156 132462
rect 191104 132398 191156 132404
rect 190092 125792 190144 125798
rect 190092 125734 190144 125740
rect 190092 125656 190144 125662
rect 190092 125598 190144 125604
rect 190104 121446 190132 125598
rect 190092 121440 190144 121446
rect 190092 121382 190144 121388
rect 190472 120329 190500 132398
rect 191208 132025 191236 165582
rect 191656 145920 191708 145926
rect 191656 145862 191708 145868
rect 191668 139913 191696 145862
rect 191654 139904 191710 139913
rect 191654 139839 191710 139848
rect 191656 136604 191708 136610
rect 191656 136546 191708 136552
rect 191668 136377 191696 136546
rect 191654 136368 191710 136377
rect 191654 136303 191710 136312
rect 191654 135552 191710 135561
rect 191654 135487 191710 135496
rect 191668 135318 191696 135487
rect 191656 135312 191708 135318
rect 191656 135254 191708 135260
rect 191194 132016 191250 132025
rect 191194 131951 191250 131960
rect 190828 131096 190880 131102
rect 190828 131038 190880 131044
rect 190840 130121 190868 131038
rect 190826 130112 190882 130121
rect 190826 130047 190882 130056
rect 191012 125792 191064 125798
rect 191010 125760 191012 125769
rect 191064 125760 191066 125769
rect 191010 125695 191066 125704
rect 191208 122834 191236 131951
rect 191654 129296 191710 129305
rect 191654 129231 191710 129240
rect 191668 128722 191696 129231
rect 191656 128716 191708 128722
rect 191656 128658 191708 128664
rect 191654 127664 191710 127673
rect 191654 127599 191710 127608
rect 191668 127022 191696 127599
rect 191656 127016 191708 127022
rect 191656 126958 191708 126964
rect 191208 122806 191696 122834
rect 191562 122224 191618 122233
rect 191562 122159 191618 122168
rect 191576 121650 191604 122159
rect 191564 121644 191616 121650
rect 191564 121586 191616 121592
rect 190826 121408 190882 121417
rect 190826 121343 190882 121352
rect 190458 120320 190514 120329
rect 190380 120278 190458 120306
rect 190274 110800 190330 110809
rect 190274 110735 190330 110744
rect 190288 108934 190316 110735
rect 190276 108928 190328 108934
rect 190276 108870 190328 108876
rect 189906 98288 189962 98297
rect 189906 98223 189962 98232
rect 189814 92304 189870 92313
rect 189814 92239 189870 92248
rect 189920 81394 189948 98223
rect 189908 81388 189960 81394
rect 189908 81330 189960 81336
rect 190380 79354 190408 120278
rect 190458 120255 190514 120264
rect 190840 120154 190868 121343
rect 190828 120148 190880 120154
rect 190828 120090 190880 120096
rect 191564 120080 191616 120086
rect 191564 120022 191616 120028
rect 191576 119513 191604 120022
rect 191562 119504 191618 119513
rect 191562 119439 191618 119448
rect 191562 118688 191618 118697
rect 191562 118623 191618 118632
rect 190826 118008 190882 118017
rect 190826 117943 190828 117952
rect 190880 117943 190882 117952
rect 190828 117914 190880 117920
rect 191576 117366 191604 118623
rect 191564 117360 191616 117366
rect 191564 117302 191616 117308
rect 191380 117224 191432 117230
rect 191380 117166 191432 117172
rect 191392 115977 191420 117166
rect 191562 116784 191618 116793
rect 191562 116719 191618 116728
rect 191576 116074 191604 116719
rect 191564 116068 191616 116074
rect 191564 116010 191616 116016
rect 191378 115968 191434 115977
rect 191378 115903 191434 115912
rect 191012 115456 191064 115462
rect 191012 115398 191064 115404
rect 191024 115161 191052 115398
rect 191010 115152 191066 115161
rect 191010 115087 191066 115096
rect 191564 114504 191616 114510
rect 191564 114446 191616 114452
rect 190826 114064 190882 114073
rect 190826 113999 190882 114008
rect 190840 113218 190868 113999
rect 191576 113257 191604 114446
rect 191562 113248 191618 113257
rect 190828 113212 190880 113218
rect 191562 113183 191618 113192
rect 190828 113154 190880 113160
rect 191564 113144 191616 113150
rect 191564 113086 191616 113092
rect 191576 112441 191604 113086
rect 191562 112432 191618 112441
rect 191562 112367 191618 112376
rect 191196 111784 191248 111790
rect 191196 111726 191248 111732
rect 191208 110537 191236 111726
rect 191194 110528 191250 110537
rect 191194 110463 191250 110472
rect 191012 110356 191064 110362
rect 191012 110298 191064 110304
rect 191024 109721 191052 110298
rect 191010 109712 191066 109721
rect 191010 109647 191066 109656
rect 190644 107636 190696 107642
rect 190644 107578 190696 107584
rect 190656 107001 190684 107578
rect 190642 106992 190698 107001
rect 190642 106927 190698 106936
rect 191012 106276 191064 106282
rect 191012 106218 191064 106224
rect 191024 106185 191052 106218
rect 191010 106176 191066 106185
rect 191010 106111 191066 106120
rect 191562 105088 191618 105097
rect 191562 105023 191618 105032
rect 191576 104922 191604 105023
rect 191564 104916 191616 104922
rect 191564 104858 191616 104864
rect 191562 103456 191618 103465
rect 191562 103391 191618 103400
rect 191470 102640 191526 102649
rect 191470 102575 191526 102584
rect 191484 102270 191512 102575
rect 191472 102264 191524 102270
rect 191472 102206 191524 102212
rect 190642 101552 190698 101561
rect 190642 101487 190698 101496
rect 190656 100774 190684 101487
rect 190644 100768 190696 100774
rect 190644 100710 190696 100716
rect 190644 97980 190696 97986
rect 190644 97922 190696 97928
rect 190656 97209 190684 97922
rect 190642 97200 190698 97209
rect 190642 97135 190698 97144
rect 190460 95260 190512 95266
rect 190460 95202 190512 95208
rect 190472 92478 190500 95202
rect 190460 92472 190512 92478
rect 190460 92414 190512 92420
rect 191484 84289 191512 102206
rect 191576 102202 191604 103391
rect 191564 102196 191616 102202
rect 191564 102138 191616 102144
rect 191562 100736 191618 100745
rect 191562 100671 191618 100680
rect 191576 99618 191604 100671
rect 191564 99612 191616 99618
rect 191564 99554 191616 99560
rect 191102 84280 191158 84289
rect 191102 84215 191158 84224
rect 191470 84280 191526 84289
rect 191470 84215 191526 84224
rect 190368 79348 190420 79354
rect 190368 79290 190420 79296
rect 191116 67590 191144 84215
rect 191668 83570 191696 122806
rect 191760 100881 191788 258046
rect 192496 248470 192524 295151
rect 192864 277817 192892 347006
rect 196636 341562 196664 355263
rect 196624 341556 196676 341562
rect 196624 341498 196676 341504
rect 193404 334620 193456 334626
rect 193404 334562 193456 334568
rect 193036 331900 193088 331906
rect 193036 331842 193088 331848
rect 192942 302288 192998 302297
rect 192942 302223 192998 302232
rect 192956 280673 192984 302223
rect 193048 296177 193076 331842
rect 193312 311160 193364 311166
rect 193312 311102 193364 311108
rect 193034 296168 193090 296177
rect 193034 296103 193090 296112
rect 193048 295390 193076 296103
rect 193036 295384 193088 295390
rect 193036 295326 193088 295332
rect 193324 295225 193352 311102
rect 193310 295216 193366 295225
rect 193310 295151 193366 295160
rect 193036 284300 193088 284306
rect 193036 284242 193088 284248
rect 193048 283529 193076 284242
rect 193034 283520 193090 283529
rect 193034 283455 193090 283464
rect 192942 280664 192998 280673
rect 192942 280599 192998 280608
rect 192850 277808 192906 277817
rect 192850 277743 192906 277752
rect 192864 277438 192892 277743
rect 192852 277432 192904 277438
rect 192852 277374 192904 277380
rect 192484 248464 192536 248470
rect 192484 248406 192536 248412
rect 192022 246256 192078 246265
rect 192022 246191 192078 246200
rect 192036 245721 192064 246191
rect 192022 245712 192078 245721
rect 192022 245647 192078 245656
rect 192496 237969 192524 248406
rect 192944 244928 192996 244934
rect 192944 244870 192996 244876
rect 192956 241398 192984 244870
rect 192944 241392 192996 241398
rect 192944 241334 192996 241340
rect 192482 237960 192538 237969
rect 192482 237895 192538 237904
rect 193048 232529 193076 283455
rect 193416 278769 193444 334562
rect 197360 332648 197412 332654
rect 197360 332590 197412 332596
rect 195702 303784 195758 303793
rect 195702 303719 195758 303728
rect 196348 303748 196400 303754
rect 194138 301608 194194 301617
rect 194194 301566 194442 301594
rect 195716 301580 195744 303719
rect 196348 303690 196400 303696
rect 196360 301580 196388 303690
rect 197372 303686 197400 332590
rect 198016 325694 198044 370466
rect 198094 367160 198150 367169
rect 198094 367095 198150 367104
rect 198108 344350 198136 367095
rect 198752 362846 198780 390374
rect 198740 362840 198792 362846
rect 198740 362782 198792 362788
rect 198752 362234 198780 362782
rect 198740 362228 198792 362234
rect 198740 362170 198792 362176
rect 200132 356697 200160 390374
rect 201144 388385 201172 390388
rect 202064 389298 202092 390388
rect 202892 390374 202998 390402
rect 204272 390374 204838 390402
rect 205652 390374 205942 390402
rect 206020 390374 206862 390402
rect 202052 389292 202104 389298
rect 202052 389234 202104 389240
rect 201130 388376 201186 388385
rect 201130 388311 201186 388320
rect 200118 356688 200174 356697
rect 200118 356623 200174 356632
rect 198096 344344 198148 344350
rect 198096 344286 198148 344292
rect 198016 325666 198136 325694
rect 197450 312080 197506 312089
rect 197450 312015 197506 312024
rect 197360 303680 197412 303686
rect 197360 303622 197412 303628
rect 197464 301594 197492 312015
rect 198004 303680 198056 303686
rect 198004 303622 198056 303628
rect 198016 301594 198044 303622
rect 198108 303521 198136 325666
rect 198740 323604 198792 323610
rect 198740 323546 198792 323552
rect 198752 323105 198780 323546
rect 198738 323096 198794 323105
rect 198738 323031 198740 323040
rect 198792 323031 198794 323040
rect 198740 323002 198792 323008
rect 198752 322971 198780 323002
rect 200132 313410 200160 356623
rect 202892 348430 202920 390374
rect 204272 379438 204300 390374
rect 204260 379432 204312 379438
rect 204260 379374 204312 379380
rect 204272 376689 204300 379374
rect 204258 376680 204314 376689
rect 204258 376615 204314 376624
rect 205546 376680 205602 376689
rect 205546 376615 205602 376624
rect 202880 348424 202932 348430
rect 202880 348366 202932 348372
rect 204260 327140 204312 327146
rect 204260 327082 204312 327088
rect 204272 325694 204300 327082
rect 204272 325666 204760 325694
rect 202326 324456 202382 324465
rect 202326 324391 202382 324400
rect 200302 316160 200358 316169
rect 200302 316095 200358 316104
rect 200120 313404 200172 313410
rect 200120 313346 200172 313352
rect 200210 309224 200266 309233
rect 200210 309159 200266 309168
rect 199474 306504 199530 306513
rect 199474 306439 199530 306448
rect 198094 303512 198150 303521
rect 198094 303447 198150 303456
rect 198832 302320 198884 302326
rect 198832 302262 198884 302268
rect 197464 301566 197662 301594
rect 198016 301566 198306 301594
rect 198844 301580 198872 302262
rect 199488 301580 199516 306439
rect 200224 303686 200252 309159
rect 200212 303680 200264 303686
rect 200212 303622 200264 303628
rect 200118 302560 200174 302569
rect 200118 302495 200174 302504
rect 200132 301580 200160 302495
rect 200316 301594 200344 316095
rect 201408 313404 201460 313410
rect 201408 313346 201460 313352
rect 201420 309874 201448 313346
rect 201408 309868 201460 309874
rect 201408 309810 201460 309816
rect 202050 307864 202106 307873
rect 202050 307799 202106 307808
rect 201132 303680 201184 303686
rect 201132 303622 201184 303628
rect 201144 301594 201172 303622
rect 201408 303612 201460 303618
rect 201408 303554 201460 303560
rect 201420 303521 201448 303554
rect 201406 303512 201462 303521
rect 201406 303447 201462 303456
rect 200316 301566 200790 301594
rect 201144 301566 201434 301594
rect 202064 301580 202092 307799
rect 202340 301594 202368 324391
rect 203430 311944 203486 311953
rect 203430 311879 203486 311888
rect 203444 301594 203472 311879
rect 204732 301594 204760 325666
rect 205560 313993 205588 376615
rect 205652 336054 205680 390374
rect 206020 373994 206048 390374
rect 207768 384985 207796 390388
rect 208412 390374 208702 390402
rect 208872 390374 209622 390402
rect 209792 390374 210542 390402
rect 211172 390374 211646 390402
rect 207754 384976 207810 384985
rect 207754 384911 207810 384920
rect 205744 373966 206048 373994
rect 205744 362914 205772 373966
rect 207112 366376 207164 366382
rect 207112 366318 207164 366324
rect 205732 362908 205784 362914
rect 205732 362850 205784 362856
rect 205640 336048 205692 336054
rect 205640 335990 205692 335996
rect 205546 313984 205602 313993
rect 205546 313919 205602 313928
rect 205744 311166 205772 362850
rect 207018 317520 207074 317529
rect 207018 317455 207074 317464
rect 205732 311160 205784 311166
rect 205732 311102 205784 311108
rect 205638 310584 205694 310593
rect 205638 310519 205694 310528
rect 205652 301594 205680 310519
rect 207032 306374 207060 317455
rect 207124 307737 207152 366318
rect 208412 337385 208440 390374
rect 208492 386368 208544 386374
rect 208492 386310 208544 386316
rect 208504 385665 208532 386310
rect 208490 385656 208546 385665
rect 208490 385591 208546 385600
rect 208872 373994 208900 390374
rect 208504 373966 208900 373994
rect 208504 367713 208532 373966
rect 208490 367704 208546 367713
rect 208490 367639 208546 367648
rect 209792 342922 209820 390374
rect 211172 356046 211200 390374
rect 212552 371929 212580 390388
rect 213472 388521 213500 390388
rect 213932 390374 214406 390402
rect 215326 390374 215432 390402
rect 213458 388512 213514 388521
rect 213458 388447 213514 388456
rect 212538 371920 212594 371929
rect 212538 371855 212594 371864
rect 213828 364404 213880 364410
rect 213828 364346 213880 364352
rect 213840 362914 213868 364346
rect 213828 362908 213880 362914
rect 213828 362850 213880 362856
rect 211160 356040 211212 356046
rect 211160 355982 211212 355988
rect 211804 356040 211856 356046
rect 211804 355982 211856 355988
rect 209780 342916 209832 342922
rect 209780 342858 209832 342864
rect 208398 337376 208454 337385
rect 208398 337311 208454 337320
rect 211816 331809 211844 355982
rect 213932 334665 213960 390374
rect 214564 387864 214616 387870
rect 214564 387806 214616 387812
rect 214576 354006 214604 387806
rect 215404 360126 215432 390374
rect 216232 387870 216260 390388
rect 216692 390374 217350 390402
rect 216220 387864 216272 387870
rect 216220 387806 216272 387812
rect 216404 385008 216456 385014
rect 216404 384950 216456 384956
rect 216416 384033 216444 384950
rect 216402 384024 216458 384033
rect 216402 383959 216458 383968
rect 216416 383722 216444 383959
rect 216404 383716 216456 383722
rect 216404 383658 216456 383664
rect 215392 360120 215444 360126
rect 215392 360062 215444 360068
rect 215404 359718 215432 360062
rect 215392 359712 215444 359718
rect 215392 359654 215444 359660
rect 215944 359712 215996 359718
rect 215944 359654 215996 359660
rect 214564 354000 214616 354006
rect 214564 353942 214616 353948
rect 213918 334656 213974 334665
rect 213918 334591 213974 334600
rect 211802 331800 211858 331809
rect 211802 331735 211858 331744
rect 211252 331288 211304 331294
rect 211252 331230 211304 331236
rect 209044 329928 209096 329934
rect 209044 329870 209096 329876
rect 208398 328536 208454 328545
rect 208398 328471 208454 328480
rect 208412 325694 208440 328471
rect 208412 325666 208624 325694
rect 207110 307728 207166 307737
rect 207110 307663 207166 307672
rect 207124 307057 207152 307663
rect 207110 307048 207166 307057
rect 207110 306983 207166 306992
rect 207032 306346 207888 306374
rect 207662 302424 207718 302433
rect 207662 302359 207718 302368
rect 202340 301566 202722 301594
rect 203444 301566 203918 301594
rect 204732 301566 205206 301594
rect 205652 301566 205850 301594
rect 207676 301580 207704 302359
rect 207860 301594 207888 306346
rect 208596 301594 208624 325666
rect 209056 304570 209084 329870
rect 210424 310616 210476 310622
rect 210424 310558 210476 310564
rect 210238 306640 210294 306649
rect 210238 306575 210294 306584
rect 209594 305280 209650 305289
rect 209594 305215 209650 305224
rect 209044 304564 209096 304570
rect 209044 304506 209096 304512
rect 207860 301566 208334 301594
rect 208596 301566 208978 301594
rect 209608 301580 209636 305215
rect 210252 301580 210280 306575
rect 210436 303618 210464 310558
rect 210424 303612 210476 303618
rect 210424 303554 210476 303560
rect 211264 301594 211292 331230
rect 215956 325825 215984 359654
rect 216692 354074 216720 390374
rect 218256 387802 218284 390388
rect 218532 390374 219190 390402
rect 219452 390374 220110 390402
rect 218244 387796 218296 387802
rect 218244 387738 218296 387744
rect 218532 373994 218560 390374
rect 219256 387796 219308 387802
rect 219256 387738 219308 387744
rect 219268 387122 219296 387738
rect 219256 387116 219308 387122
rect 219256 387058 219308 387064
rect 218072 373966 218560 373994
rect 216680 354068 216732 354074
rect 216680 354010 216732 354016
rect 218072 352578 218100 373966
rect 219452 361593 219480 390374
rect 221016 384334 221044 390388
rect 221292 390374 221950 390402
rect 222212 390374 222870 390402
rect 223684 390374 223974 390402
rect 224512 390374 224894 390402
rect 224972 390374 225814 390402
rect 226352 390374 226734 390402
rect 226904 390374 227654 390402
rect 221004 384328 221056 384334
rect 221004 384270 221056 384276
rect 221292 380866 221320 390374
rect 221280 380860 221332 380866
rect 221280 380802 221332 380808
rect 219438 361584 219494 361593
rect 219438 361519 219494 361528
rect 218060 352572 218112 352578
rect 218060 352514 218112 352520
rect 220084 334008 220136 334014
rect 220084 333950 220136 333956
rect 215942 325816 215998 325825
rect 215942 325751 215998 325760
rect 215956 324970 215984 325751
rect 215944 324964 215996 324970
rect 215944 324906 215996 324912
rect 211804 319456 211856 319462
rect 211804 319398 211856 319404
rect 211816 312497 211844 319398
rect 216218 318064 216274 318073
rect 216218 317999 216274 318008
rect 214288 314764 214340 314770
rect 214288 314706 214340 314712
rect 211802 312488 211858 312497
rect 211802 312423 211858 312432
rect 212722 308136 212778 308145
rect 212722 308071 212778 308080
rect 212172 304564 212224 304570
rect 212172 304506 212224 304512
rect 211264 301566 211554 301594
rect 212184 301580 212212 304506
rect 212736 301580 212764 308071
rect 214010 305144 214066 305153
rect 214010 305079 214066 305088
rect 213366 303920 213422 303929
rect 213366 303855 213422 303864
rect 213380 301580 213408 303855
rect 214024 301580 214052 305079
rect 214300 301594 214328 314706
rect 216232 311273 216260 317999
rect 216218 311264 216274 311273
rect 216218 311199 216274 311208
rect 219990 310720 220046 310729
rect 219990 310655 220046 310664
rect 217416 309188 217468 309194
rect 217416 309130 217468 309136
rect 215300 307896 215352 307902
rect 215300 307838 215352 307844
rect 214300 301566 214682 301594
rect 215312 301580 215340 307838
rect 215944 306468 215996 306474
rect 215944 306410 215996 306416
rect 215956 301580 215984 306410
rect 216588 305108 216640 305114
rect 216588 305050 216640 305056
rect 216600 301580 216628 305050
rect 217428 301594 217456 309130
rect 218058 308408 218114 308417
rect 218058 308343 218114 308352
rect 218072 303657 218100 308343
rect 219716 307828 219768 307834
rect 219716 307770 219768 307776
rect 219072 305040 219124 305046
rect 219072 304982 219124 304988
rect 218058 303648 218114 303657
rect 218058 303583 218114 303592
rect 218428 302252 218480 302258
rect 218428 302194 218480 302200
rect 217428 301566 217810 301594
rect 218440 301580 218468 302194
rect 219084 301580 219112 304982
rect 219728 301580 219756 307770
rect 220004 301594 220032 310655
rect 220096 307766 220124 333950
rect 220818 313304 220874 313313
rect 220818 313239 220874 313248
rect 220084 307760 220136 307766
rect 220084 307702 220136 307708
rect 220832 301594 220860 313239
rect 222212 307737 222240 390374
rect 223580 387048 223632 387054
rect 223580 386990 223632 386996
rect 223488 381540 223540 381546
rect 223488 381482 223540 381488
rect 223500 380866 223528 381482
rect 223488 380860 223540 380866
rect 223488 380802 223540 380808
rect 223500 329934 223528 380802
rect 223488 329928 223540 329934
rect 223488 329870 223540 329876
rect 223500 326369 223528 329870
rect 223486 326360 223542 326369
rect 223486 326295 223542 326304
rect 223118 314800 223174 314809
rect 223118 314735 223174 314744
rect 222198 307728 222254 307737
rect 222198 307663 222254 307672
rect 221554 306776 221610 306785
rect 221554 306711 221610 306720
rect 220004 301566 220386 301594
rect 220832 301566 221030 301594
rect 221568 301580 221596 306711
rect 222566 301608 222622 301617
rect 194138 301543 194194 301552
rect 223132 301594 223160 314735
rect 223592 309806 223620 386990
rect 223684 333266 223712 390374
rect 224512 387054 224540 390374
rect 224500 387048 224552 387054
rect 224500 386990 224552 386996
rect 224972 375358 225000 390374
rect 224960 375352 225012 375358
rect 224960 375294 225012 375300
rect 226352 368490 226380 390374
rect 226904 383654 226932 390374
rect 228560 389230 228588 390388
rect 229112 390374 229678 390402
rect 230492 390374 230598 390402
rect 230768 390374 231518 390402
rect 231872 390374 232438 390402
rect 227720 389224 227772 389230
rect 227720 389166 227772 389172
rect 228548 389224 228600 389230
rect 228548 389166 228600 389172
rect 226904 383626 227024 383654
rect 226996 382294 227024 383626
rect 226984 382288 227036 382294
rect 226984 382230 227036 382236
rect 226996 373318 227024 382230
rect 226984 373312 227036 373318
rect 226984 373254 227036 373260
rect 226340 368484 226392 368490
rect 226340 368426 226392 368432
rect 226984 368484 227036 368490
rect 226984 368426 227036 368432
rect 223672 333260 223724 333266
rect 223672 333202 223724 333208
rect 226996 327758 227024 368426
rect 226984 327752 227036 327758
rect 226984 327694 227036 327700
rect 226984 311976 227036 311982
rect 226984 311918 227036 311924
rect 223580 309800 223632 309806
rect 223580 309742 223632 309748
rect 224776 307760 224828 307766
rect 224776 307702 224828 307708
rect 222622 301566 222870 301594
rect 223132 301566 223514 301594
rect 224788 301580 224816 307702
rect 226996 305658 227024 311918
rect 226984 305652 227036 305658
rect 226984 305594 227036 305600
rect 227732 305153 227760 389166
rect 228362 338736 228418 338745
rect 228362 338671 228418 338680
rect 227810 331256 227866 331265
rect 227810 331191 227866 331200
rect 227718 305144 227774 305153
rect 227718 305079 227774 305088
rect 225050 301880 225106 301889
rect 225050 301815 225106 301824
rect 225064 301594 225092 301815
rect 226982 301608 227038 301617
rect 225064 301566 225446 301594
rect 222566 301543 222622 301552
rect 227824 301594 227852 331191
rect 228376 324970 228404 338671
rect 229112 334626 229140 390374
rect 229100 334620 229152 334626
rect 229100 334562 229152 334568
rect 228364 324964 228416 324970
rect 228364 324906 228416 324912
rect 229744 318844 229796 318850
rect 229744 318786 229796 318792
rect 229756 315314 229784 318786
rect 229744 315308 229796 315314
rect 229744 315250 229796 315256
rect 230492 308446 230520 390374
rect 230768 380934 230796 390374
rect 231124 386368 231176 386374
rect 231124 386310 231176 386316
rect 230756 380928 230808 380934
rect 230756 380870 230808 380876
rect 230768 377466 230796 380870
rect 230756 377460 230808 377466
rect 230756 377402 230808 377408
rect 231136 362914 231164 386310
rect 231872 385082 231900 390374
rect 233344 387870 233372 390388
rect 234066 389464 234122 389473
rect 234066 389399 234122 389408
rect 234080 388754 234108 389399
rect 234068 388748 234120 388754
rect 234068 388690 234120 388696
rect 232504 387864 232556 387870
rect 232504 387806 232556 387812
rect 233332 387864 233384 387870
rect 233332 387806 233384 387812
rect 231860 385076 231912 385082
rect 231860 385018 231912 385024
rect 231872 382974 231900 385018
rect 231860 382968 231912 382974
rect 231860 382910 231912 382916
rect 231124 362908 231176 362914
rect 231124 362850 231176 362856
rect 231122 355464 231178 355473
rect 231122 355399 231178 355408
rect 231136 319462 231164 355399
rect 231124 319456 231176 319462
rect 231124 319398 231176 319404
rect 232516 316713 232544 387806
rect 232596 387116 232648 387122
rect 232596 387058 232648 387064
rect 232608 358057 232636 387058
rect 234264 386374 234292 390388
rect 234908 390374 235382 390402
rect 234908 389230 234936 390374
rect 234896 389224 234948 389230
rect 234896 389166 234948 389172
rect 234528 388748 234580 388754
rect 234528 388690 234580 388696
rect 234252 386368 234304 386374
rect 234252 386310 234304 386316
rect 233882 384296 233938 384305
rect 233882 384231 233938 384240
rect 232594 358048 232650 358057
rect 232594 357983 232650 357992
rect 233896 331906 233924 384231
rect 233884 331900 233936 331906
rect 233884 331842 233936 331848
rect 234540 326398 234568 388690
rect 234908 373994 234936 389166
rect 236288 386481 236316 390388
rect 236656 390374 237222 390402
rect 237392 390374 238142 390402
rect 236274 386472 236330 386481
rect 236274 386407 236330 386416
rect 236656 373994 236684 390374
rect 234632 373966 234936 373994
rect 236012 373966 236684 373994
rect 234632 358766 234660 373966
rect 236012 371210 236040 373966
rect 236000 371204 236052 371210
rect 236000 371146 236052 371152
rect 236012 369918 236040 371146
rect 237392 370569 237420 390374
rect 239048 388754 239076 390388
rect 239140 390374 239982 390402
rect 239036 388748 239088 388754
rect 239036 388690 239088 388696
rect 238114 384432 238170 384441
rect 238114 384367 238170 384376
rect 237378 370560 237434 370569
rect 237378 370495 237434 370504
rect 236000 369912 236052 369918
rect 236000 369854 236052 369860
rect 236644 369912 236696 369918
rect 237392 369889 237420 370495
rect 236644 369854 236696 369860
rect 237378 369880 237434 369889
rect 234620 358760 234672 358766
rect 234620 358702 234672 358708
rect 235264 358760 235316 358766
rect 235264 358702 235316 358708
rect 234528 326392 234580 326398
rect 234528 326334 234580 326340
rect 233884 317484 233936 317490
rect 233884 317426 233936 317432
rect 232502 316704 232558 316713
rect 232502 316639 232558 316648
rect 232504 309868 232556 309874
rect 232504 309810 232556 309816
rect 230480 308440 230532 308446
rect 230480 308382 230532 308388
rect 232516 304366 232544 309810
rect 233896 305697 233924 317426
rect 235276 314129 235304 358702
rect 236656 337414 236684 369854
rect 237378 369815 237434 369824
rect 238022 369880 238078 369889
rect 238022 369815 238078 369824
rect 236644 337408 236696 337414
rect 236644 337350 236696 337356
rect 236644 336048 236696 336054
rect 236644 335990 236696 335996
rect 235262 314120 235318 314129
rect 235262 314055 235318 314064
rect 236656 307086 236684 335990
rect 238036 331906 238064 369815
rect 238128 347070 238156 384367
rect 239140 382226 239168 390374
rect 241072 389337 241100 390388
rect 240138 389328 240194 389337
rect 240138 389263 240194 389272
rect 241058 389328 241114 389337
rect 241058 389263 241114 389272
rect 239404 382356 239456 382362
rect 239404 382298 239456 382304
rect 239128 382220 239180 382226
rect 239128 382162 239180 382168
rect 238116 347064 238168 347070
rect 238116 347006 238168 347012
rect 239416 345710 239444 382298
rect 239404 345704 239456 345710
rect 239404 345646 239456 345652
rect 238116 333260 238168 333266
rect 238116 333202 238168 333208
rect 238024 331900 238076 331906
rect 238024 331842 238076 331848
rect 238128 307193 238156 333202
rect 240152 308514 240180 389263
rect 241992 389094 242020 390388
rect 242164 389836 242216 389842
rect 242164 389778 242216 389784
rect 241980 389088 242032 389094
rect 241980 389030 242032 389036
rect 241992 387870 242020 389030
rect 241980 387864 242032 387870
rect 241980 387806 242032 387812
rect 240232 383716 240284 383722
rect 240232 383658 240284 383664
rect 240244 379506 240272 383658
rect 240232 379500 240284 379506
rect 240232 379442 240284 379448
rect 242176 373998 242204 389778
rect 242808 387864 242860 387870
rect 242808 387806 242860 387812
rect 242164 373992 242216 373998
rect 242164 373934 242216 373940
rect 240784 373312 240836 373318
rect 240784 373254 240836 373260
rect 240796 329866 240824 373254
rect 240876 340196 240928 340202
rect 240876 340138 240928 340144
rect 240232 329860 240284 329866
rect 240232 329802 240284 329808
rect 240784 329860 240836 329866
rect 240784 329802 240836 329808
rect 240140 308508 240192 308514
rect 240140 308450 240192 308456
rect 238114 307184 238170 307193
rect 238114 307119 238170 307128
rect 236644 307080 236696 307086
rect 236644 307022 236696 307028
rect 239312 306400 239364 306406
rect 239312 306342 239364 306348
rect 233882 305688 233938 305697
rect 233882 305623 233938 305632
rect 232504 304360 232556 304366
rect 232504 304302 232556 304308
rect 231032 303816 231084 303822
rect 229190 303784 229246 303793
rect 231032 303758 231084 303764
rect 229190 303719 229246 303728
rect 227038 301566 227286 301594
rect 227824 301566 227930 301594
rect 229204 301580 229232 303719
rect 230112 303680 230164 303686
rect 230112 303622 230164 303628
rect 229834 302288 229890 302297
rect 229834 302223 229890 302232
rect 229848 301580 229876 302223
rect 226982 301543 227038 301552
rect 230124 301481 230152 303622
rect 231044 301580 231072 303758
rect 238668 303680 238720 303686
rect 238668 303622 238720 303628
rect 236090 302288 236146 302297
rect 236090 302223 236146 302232
rect 231306 301608 231362 301617
rect 235262 301608 235318 301617
rect 231362 301566 231702 301594
rect 231306 301543 231362 301552
rect 235318 301566 235474 301594
rect 236104 301580 236132 302223
rect 237746 301608 237802 301617
rect 235262 301543 235318 301552
rect 237802 301566 238050 301594
rect 238680 301580 238708 303622
rect 239324 301580 239352 306342
rect 240244 301753 240272 329802
rect 240888 303657 240916 340138
rect 241796 307080 241848 307086
rect 241796 307022 241848 307028
rect 240874 303648 240930 303657
rect 240874 303583 240930 303592
rect 241150 302288 241206 302297
rect 241150 302223 241206 302232
rect 241060 302184 241112 302190
rect 241060 302126 241112 302132
rect 241072 301753 241100 302126
rect 240230 301744 240286 301753
rect 240230 301679 240286 301688
rect 241058 301744 241114 301753
rect 241058 301679 241114 301688
rect 241164 301580 241192 302223
rect 241808 301580 241836 307022
rect 242176 306406 242204 373934
rect 242820 357406 242848 387806
rect 242912 372570 242940 390388
rect 243832 383722 243860 390388
rect 244292 390374 244766 390402
rect 242992 383716 243044 383722
rect 242992 383658 243044 383664
rect 243820 383716 243872 383722
rect 243820 383658 243872 383664
rect 244004 383716 244056 383722
rect 244004 383658 244056 383664
rect 243004 383625 243032 383658
rect 244016 383625 244044 383658
rect 242990 383616 243046 383625
rect 242990 383551 243046 383560
rect 244002 383616 244058 383625
rect 244002 383551 244058 383560
rect 244292 382362 244320 390374
rect 244924 384328 244976 384334
rect 244924 384270 244976 384276
rect 244280 382356 244332 382362
rect 244280 382298 244332 382304
rect 244370 380216 244426 380225
rect 244370 380151 244426 380160
rect 242900 372564 242952 372570
rect 242900 372506 242952 372512
rect 242912 371278 242940 372506
rect 242900 371272 242952 371278
rect 242900 371214 242952 371220
rect 243544 371272 243596 371278
rect 243544 371214 243596 371220
rect 243556 359514 243584 371214
rect 243544 359508 243596 359514
rect 243544 359450 243596 359456
rect 242808 357400 242860 357406
rect 242808 357342 242860 357348
rect 242820 356726 242848 357342
rect 242808 356720 242860 356726
rect 242808 356662 242860 356668
rect 244278 353968 244334 353977
rect 244278 353903 244334 353912
rect 242992 351280 243044 351286
rect 242992 351222 243044 351228
rect 243004 325694 243032 351222
rect 244292 340950 244320 353903
rect 244280 340944 244332 340950
rect 244280 340886 244332 340892
rect 243004 325666 243400 325694
rect 242164 306400 242216 306406
rect 242164 306342 242216 306348
rect 242176 301594 242204 306342
rect 242806 304192 242862 304201
rect 242862 304150 242940 304178
rect 242806 304127 242862 304136
rect 242912 301594 242940 304150
rect 242176 301566 242466 301594
rect 242912 301566 243110 301594
rect 237746 301543 237802 301552
rect 203062 301472 203118 301481
rect 204350 301472 204406 301481
rect 203118 301430 203274 301458
rect 203062 301407 203118 301416
rect 207018 301472 207074 301481
rect 204406 301430 204562 301458
rect 204350 301407 204406 301416
rect 210606 301472 210662 301481
rect 207074 301430 207138 301458
rect 207018 301407 207074 301416
rect 216770 301472 216826 301481
rect 210662 301430 210910 301458
rect 210606 301407 210662 301416
rect 222566 301472 222622 301481
rect 216826 301430 217166 301458
rect 222226 301430 222566 301458
rect 216770 301407 216826 301416
rect 222566 301407 222622 301416
rect 223854 301472 223910 301481
rect 225786 301472 225842 301481
rect 223910 301430 224158 301458
rect 223854 301407 223910 301416
rect 226706 301472 226762 301481
rect 225842 301430 226090 301458
rect 226642 301430 226706 301458
rect 225786 301407 225842 301416
rect 226706 301407 226762 301416
rect 228270 301472 228326 301481
rect 230110 301472 230166 301481
rect 228326 301430 228574 301458
rect 228270 301407 228326 301416
rect 230570 301472 230626 301481
rect 230506 301430 230570 301458
rect 230110 301407 230166 301416
rect 230570 301407 230626 301416
rect 232134 301472 232190 301481
rect 232686 301472 232742 301481
rect 232190 301430 232346 301458
rect 232134 301407 232190 301416
rect 233330 301472 233386 301481
rect 232742 301430 232990 301458
rect 232686 301407 232742 301416
rect 233974 301472 234030 301481
rect 233386 301430 233634 301458
rect 233330 301407 233386 301416
rect 234802 301472 234858 301481
rect 234030 301430 234278 301458
rect 233974 301407 234030 301416
rect 236642 301472 236698 301481
rect 234858 301430 234922 301458
rect 234802 301407 234858 301416
rect 237654 301472 237710 301481
rect 236698 301430 236762 301458
rect 237406 301430 237654 301458
rect 236642 301407 236698 301416
rect 237654 301407 237710 301416
rect 239678 301472 239734 301481
rect 243372 301458 243400 325666
rect 244292 303686 244320 340886
rect 244384 329905 244412 380151
rect 244936 379370 244964 384270
rect 244924 379364 244976 379370
rect 244924 379306 244976 379312
rect 244370 329896 244426 329905
rect 244370 329831 244426 329840
rect 244280 303680 244332 303686
rect 244280 303622 244332 303628
rect 244384 301580 244412 329831
rect 244462 314936 244518 314945
rect 244462 314871 244518 314880
rect 244476 307086 244504 314871
rect 244936 311982 244964 379306
rect 245672 360194 245700 390388
rect 245764 390374 246606 390402
rect 245764 378214 245792 390374
rect 247696 388385 247724 390388
rect 248432 390374 248630 390402
rect 248708 390374 249550 390402
rect 249996 390374 250470 390402
rect 247038 388376 247094 388385
rect 247038 388311 247094 388320
rect 247682 388376 247738 388385
rect 247682 388311 247738 388320
rect 247052 387705 247080 388311
rect 247038 387696 247094 387705
rect 247038 387631 247094 387640
rect 247684 383716 247736 383722
rect 247684 383658 247736 383664
rect 246396 380180 246448 380186
rect 246396 380122 246448 380128
rect 245752 378208 245804 378214
rect 245752 378150 245804 378156
rect 246304 378208 246356 378214
rect 246304 378150 246356 378156
rect 245844 369776 245896 369782
rect 245844 369718 245896 369724
rect 245856 369374 245884 369718
rect 245844 369368 245896 369374
rect 245844 369310 245896 369316
rect 245750 363624 245806 363633
rect 245750 363559 245806 363568
rect 245660 360188 245712 360194
rect 245660 360130 245712 360136
rect 245672 359718 245700 360130
rect 245660 359712 245712 359718
rect 245660 359654 245712 359660
rect 244556 311976 244608 311982
rect 244556 311918 244608 311924
rect 244924 311976 244976 311982
rect 244924 311918 244976 311924
rect 244568 308417 244596 311918
rect 244554 308408 244610 308417
rect 244554 308343 244610 308352
rect 244464 307080 244516 307086
rect 244464 307022 244516 307028
rect 244556 303680 244608 303686
rect 244556 303622 244608 303628
rect 245566 303648 245622 303657
rect 244568 301594 244596 303622
rect 245566 303583 245622 303592
rect 244568 301566 244950 301594
rect 245580 301580 245608 303583
rect 245764 301753 245792 363559
rect 245856 306513 245884 369310
rect 246316 365702 246344 378150
rect 246408 369374 246436 380122
rect 246396 369368 246448 369374
rect 246396 369310 246448 369316
rect 246304 365696 246356 365702
rect 246304 365638 246356 365644
rect 246304 359712 246356 359718
rect 246304 359654 246356 359660
rect 246316 308553 246344 359654
rect 247696 341630 247724 383658
rect 248432 372502 248460 390374
rect 248708 379409 248736 390374
rect 249706 390280 249762 390289
rect 249706 390215 249762 390224
rect 249248 389292 249300 389298
rect 249248 389234 249300 389240
rect 248694 379400 248750 379409
rect 248694 379335 248750 379344
rect 249062 379400 249118 379409
rect 249062 379335 249118 379344
rect 248420 372496 248472 372502
rect 248420 372438 248472 372444
rect 247684 341624 247736 341630
rect 247684 341566 247736 341572
rect 249076 316713 249104 379335
rect 249260 353258 249288 389234
rect 249720 389230 249748 390215
rect 249708 389224 249760 389230
rect 249996 389201 250024 390374
rect 249708 389166 249760 389172
rect 249982 389192 250038 389201
rect 249982 389127 250038 389136
rect 249996 378049 250024 389127
rect 249982 378040 250038 378049
rect 249982 377975 250038 377984
rect 250444 372496 250496 372502
rect 250444 372438 250496 372444
rect 249248 353252 249300 353258
rect 249248 353194 249300 353200
rect 249156 352572 249208 352578
rect 249156 352514 249208 352520
rect 249062 316704 249118 316713
rect 249062 316639 249118 316648
rect 246302 308544 246358 308553
rect 246302 308479 246358 308488
rect 245842 306504 245898 306513
rect 245842 306439 245898 306448
rect 245750 301744 245806 301753
rect 245750 301679 245806 301688
rect 245856 301594 245884 306439
rect 247500 304292 247552 304298
rect 247500 304234 247552 304240
rect 246486 301608 246542 301617
rect 245856 301566 246238 301594
rect 247512 301580 247540 304234
rect 248786 302424 248842 302433
rect 248786 302359 248842 302368
rect 248800 301580 248828 302359
rect 246486 301543 246542 301552
rect 243450 301472 243506 301481
rect 239734 301430 239982 301458
rect 243372 301430 243450 301458
rect 239678 301407 239734 301416
rect 243506 301430 243754 301458
rect 243450 301407 243506 301416
rect 246500 301374 246528 301543
rect 246578 301472 246634 301481
rect 247866 301472 247922 301481
rect 246634 301430 246882 301458
rect 246578 301407 246634 301416
rect 247922 301430 248170 301458
rect 247866 301407 247922 301416
rect 249168 301374 249196 352514
rect 249706 336696 249762 336705
rect 249706 336631 249762 336640
rect 249614 321736 249670 321745
rect 249614 321671 249670 321680
rect 249338 307728 249394 307737
rect 249338 307663 249394 307672
rect 249352 306513 249380 307663
rect 249338 306504 249394 306513
rect 249338 306439 249394 306448
rect 249352 301580 249380 306439
rect 249628 302433 249656 321671
rect 249720 307737 249748 336631
rect 249706 307728 249762 307737
rect 249706 307663 249762 307672
rect 250456 303226 250484 372438
rect 250548 349110 250576 390934
rect 251284 390374 251390 390402
rect 251836 390374 252310 390402
rect 251284 360913 251312 390374
rect 251836 389162 251864 390374
rect 251914 389192 251970 389201
rect 251824 389156 251876 389162
rect 251914 389127 251970 389136
rect 251824 389098 251876 389104
rect 251270 360904 251326 360913
rect 251270 360839 251326 360848
rect 250536 349104 250588 349110
rect 250536 349046 250588 349052
rect 250536 344344 250588 344350
rect 250536 344286 250588 344292
rect 250548 314090 250576 344286
rect 251836 326466 251864 389098
rect 251928 380866 251956 389127
rect 253400 387122 253428 390388
rect 253388 387116 253440 387122
rect 253388 387058 253440 387064
rect 251916 380860 251968 380866
rect 251916 380802 251968 380808
rect 253584 373994 253612 391546
rect 253676 389298 253704 392799
rect 253664 389292 253716 389298
rect 253664 389234 253716 389240
rect 253492 373966 253612 373994
rect 252560 368416 252612 368422
rect 252558 368384 252560 368393
rect 252612 368384 252614 368393
rect 252558 368319 252614 368328
rect 253492 349858 253520 373966
rect 253952 364993 253980 431967
rect 254044 391610 254072 451318
rect 254136 447545 254164 459575
rect 255318 455560 255374 455569
rect 255318 455495 255374 455504
rect 254674 451344 254730 451353
rect 254674 451279 254730 451288
rect 254122 447536 254178 447545
rect 254122 447471 254178 447480
rect 254582 447536 254638 447545
rect 254582 447471 254638 447480
rect 254596 432614 254624 447471
rect 254688 442270 254716 451279
rect 255332 444825 255360 455495
rect 255318 444816 255374 444825
rect 255318 444751 255374 444760
rect 254676 442264 254728 442270
rect 254676 442206 254728 442212
rect 255134 442096 255190 442105
rect 255134 442031 255190 442040
rect 254584 432608 254636 432614
rect 254584 432550 254636 432556
rect 255148 429894 255176 442031
rect 255226 436792 255282 436801
rect 255226 436727 255282 436736
rect 255136 429888 255188 429894
rect 255136 429830 255188 429836
rect 255240 424289 255268 436727
rect 255226 424280 255282 424289
rect 255226 424215 255282 424224
rect 254122 413808 254178 413817
rect 254122 413743 254178 413752
rect 254032 391604 254084 391610
rect 254032 391546 254084 391552
rect 254030 391504 254086 391513
rect 254030 391439 254086 391448
rect 253938 364984 253994 364993
rect 253938 364919 253994 364928
rect 254044 364342 254072 391439
rect 254136 389842 254164 413743
rect 254214 402656 254270 402665
rect 254214 402591 254270 402600
rect 254124 389836 254176 389842
rect 254124 389778 254176 389784
rect 254228 380186 254256 402591
rect 254216 380180 254268 380186
rect 254216 380122 254268 380128
rect 254032 364336 254084 364342
rect 254032 364278 254084 364284
rect 254044 362982 254072 364278
rect 254032 362976 254084 362982
rect 254032 362918 254084 362924
rect 254584 356720 254636 356726
rect 254584 356662 254636 356668
rect 253480 349852 253532 349858
rect 253480 349794 253532 349800
rect 252744 348424 252796 348430
rect 252744 348366 252796 348372
rect 251916 341556 251968 341562
rect 251916 341498 251968 341504
rect 251824 326460 251876 326466
rect 251824 326402 251876 326408
rect 250628 325712 250680 325718
rect 250628 325654 250680 325660
rect 250536 314084 250588 314090
rect 250536 314026 250588 314032
rect 250640 305046 250668 325654
rect 250718 313440 250774 313449
rect 250718 313375 250774 313384
rect 250628 305040 250680 305046
rect 250628 304982 250680 304988
rect 250456 303198 250668 303226
rect 249614 302424 249670 302433
rect 249614 302359 249670 302368
rect 250640 302326 250668 303198
rect 250732 302841 250760 313375
rect 251928 308417 251956 341498
rect 252558 338056 252614 338065
rect 252558 337991 252614 338000
rect 252572 336802 252600 337991
rect 252560 336796 252612 336802
rect 252560 336738 252612 336744
rect 252468 334620 252520 334626
rect 252468 334562 252520 334568
rect 252008 326392 252060 326398
rect 252008 326334 252060 326340
rect 251914 308408 251970 308417
rect 251914 308343 251970 308352
rect 251270 307184 251326 307193
rect 251270 307119 251326 307128
rect 251284 303657 251312 307119
rect 251914 303920 251970 303929
rect 251914 303855 251970 303864
rect 251270 303648 251326 303657
rect 251270 303583 251326 303592
rect 250718 302832 250774 302841
rect 250718 302767 250774 302776
rect 250628 302320 250680 302326
rect 250628 302262 250680 302268
rect 250640 301580 250668 302262
rect 251284 301580 251312 303583
rect 251928 301580 251956 303855
rect 252020 302258 252048 326334
rect 252480 304298 252508 334562
rect 252572 321745 252600 336738
rect 252558 321736 252614 321745
rect 252558 321671 252614 321680
rect 252652 304360 252704 304366
rect 252652 304302 252704 304308
rect 252468 304292 252520 304298
rect 252468 304234 252520 304240
rect 252008 302252 252060 302258
rect 252008 302194 252060 302200
rect 252664 301594 252692 304302
rect 252586 301566 252692 301594
rect 250258 301472 250314 301481
rect 250010 301430 250258 301458
rect 250258 301407 250314 301416
rect 196716 301368 196768 301374
rect 240140 301368 240192 301374
rect 196768 301316 197018 301322
rect 196716 301310 197018 301316
rect 246488 301368 246540 301374
rect 240192 301316 240534 301322
rect 240140 301310 240534 301316
rect 246488 301310 246540 301316
rect 249156 301368 249208 301374
rect 249156 301310 249208 301316
rect 196728 301294 197018 301310
rect 240152 301294 240534 301310
rect 193600 300886 193890 300914
rect 193600 298761 193628 300886
rect 195072 300830 195100 300900
rect 206480 300830 206508 300900
rect 195060 300824 195112 300830
rect 195060 300766 195112 300772
rect 206468 300824 206520 300830
rect 206468 300766 206520 300772
rect 252756 299474 252784 348366
rect 253296 335368 253348 335374
rect 253296 335310 253348 335316
rect 252928 305040 252980 305046
rect 252928 304982 252980 304988
rect 252836 300824 252888 300830
rect 252836 300766 252888 300772
rect 252848 300257 252876 300766
rect 252834 300248 252890 300257
rect 252834 300183 252890 300192
rect 252756 299446 252876 299474
rect 193586 298752 193642 298761
rect 193586 298687 193642 298696
rect 252848 296993 252876 299446
rect 252834 296984 252890 296993
rect 252834 296919 252890 296928
rect 252834 296576 252890 296585
rect 252834 296511 252890 296520
rect 252848 296426 252876 296511
rect 252664 296398 252876 296426
rect 193126 278760 193182 278769
rect 193126 278695 193182 278704
rect 193402 278760 193458 278769
rect 193402 278695 193458 278704
rect 193034 232520 193090 232529
rect 193034 232455 193090 232464
rect 193140 210361 193168 278695
rect 193220 277364 193272 277370
rect 193220 277306 193272 277312
rect 193232 276865 193260 277306
rect 193218 276856 193274 276865
rect 193218 276791 193274 276800
rect 193232 237454 193260 276791
rect 193402 258904 193458 258913
rect 193402 258839 193458 258848
rect 193416 258058 193444 258839
rect 193404 258052 193456 258058
rect 193404 257994 193456 258000
rect 193680 246356 193732 246362
rect 193680 246298 193732 246304
rect 193692 246242 193720 246298
rect 193692 246214 193812 246242
rect 193678 242856 193734 242865
rect 193678 242791 193734 242800
rect 193220 237448 193272 237454
rect 193220 237390 193272 237396
rect 193692 235822 193720 242791
rect 193680 235816 193732 235822
rect 193680 235758 193732 235764
rect 193126 210352 193182 210361
rect 193126 210287 193182 210296
rect 192944 199436 192996 199442
rect 192944 199378 192996 199384
rect 192482 153096 192538 153105
rect 192482 153031 192538 153040
rect 192496 137329 192524 153031
rect 192574 144936 192630 144945
rect 192574 144871 192630 144880
rect 192588 137834 192616 144871
rect 192956 138281 192984 199378
rect 193784 188358 193812 246214
rect 195256 240106 195284 241604
rect 198016 241590 198582 241618
rect 201604 241604 201894 241618
rect 201604 241590 201908 241604
rect 195244 240100 195296 240106
rect 195244 240042 195296 240048
rect 194784 235816 194836 235822
rect 194784 235758 194836 235764
rect 193772 188352 193824 188358
rect 193772 188294 193824 188300
rect 193218 178664 193274 178673
rect 193218 178599 193274 178608
rect 193036 160812 193088 160818
rect 193036 160754 193088 160760
rect 192666 138272 192722 138281
rect 192666 138207 192722 138216
rect 192942 138272 192998 138281
rect 192942 138207 192998 138216
rect 192576 137828 192628 137834
rect 192576 137770 192628 137776
rect 192482 137320 192538 137329
rect 192482 137255 192538 137264
rect 192482 134736 192538 134745
rect 192482 134671 192538 134680
rect 192496 133890 192524 134671
rect 192484 133884 192536 133890
rect 192484 133826 192536 133832
rect 191746 100872 191802 100881
rect 191746 100807 191802 100816
rect 191748 100700 191800 100706
rect 191748 100642 191800 100648
rect 191760 99929 191788 100642
rect 191746 99920 191802 99929
rect 191746 99855 191802 99864
rect 191748 98048 191800 98054
rect 191746 98016 191748 98025
rect 191800 98016 191802 98025
rect 191746 97951 191802 97960
rect 191748 93220 191800 93226
rect 191748 93162 191800 93168
rect 191656 83564 191708 83570
rect 191656 83506 191708 83512
rect 191104 67584 191156 67590
rect 191104 67526 191156 67532
rect 189724 53100 189776 53106
rect 189724 53042 189776 53048
rect 188344 46912 188396 46918
rect 188344 46854 188396 46860
rect 186964 40724 187016 40730
rect 186964 40666 187016 40672
rect 191760 21418 191788 93162
rect 192496 62830 192524 133826
rect 192680 132494 192708 138207
rect 192588 132466 192708 132494
rect 192588 132161 192616 132466
rect 192574 132152 192630 132161
rect 192574 132087 192630 132096
rect 192588 86193 192616 132087
rect 193048 123865 193076 160754
rect 193126 126576 193182 126585
rect 193126 126511 193182 126520
rect 193140 125662 193168 126511
rect 193128 125656 193180 125662
rect 193128 125598 193180 125604
rect 193034 123856 193090 123865
rect 193034 123791 193090 123800
rect 193048 122874 193076 123791
rect 193036 122868 193088 122874
rect 193036 122810 193088 122816
rect 193034 96384 193090 96393
rect 193034 96319 193090 96328
rect 192574 86184 192630 86193
rect 192574 86119 192630 86128
rect 193048 78441 193076 96319
rect 193034 78432 193090 78441
rect 193034 78367 193090 78376
rect 193048 69018 193076 78367
rect 192576 69012 192628 69018
rect 192576 68954 192628 68960
rect 193036 69012 193088 69018
rect 193036 68954 193088 68960
rect 192484 62824 192536 62830
rect 192484 62766 192536 62772
rect 192588 28286 192616 68954
rect 193140 68338 193168 125598
rect 193232 104281 193260 178599
rect 194508 169788 194560 169794
rect 194508 169730 194560 169736
rect 194520 168434 194548 169730
rect 193864 168428 193916 168434
rect 193864 168370 193916 168376
rect 194508 168428 194560 168434
rect 194508 168370 194560 168376
rect 193772 146396 193824 146402
rect 193772 146338 193824 146344
rect 193402 145752 193458 145761
rect 193402 145687 193458 145696
rect 193416 140978 193444 145687
rect 193784 140978 193812 146338
rect 193876 145926 193904 168370
rect 194600 158840 194652 158846
rect 194600 158782 194652 158788
rect 194612 147014 194640 158782
rect 194600 147008 194652 147014
rect 194600 146950 194652 146956
rect 193864 145920 193916 145926
rect 193864 145862 193916 145868
rect 193416 140950 193614 140978
rect 193784 140950 194166 140978
rect 194598 140584 194654 140593
rect 194654 140542 194718 140570
rect 194598 140519 194654 140528
rect 194796 140486 194824 235758
rect 195152 235272 195204 235278
rect 195152 235214 195204 235220
rect 195164 234530 195192 235214
rect 195152 234524 195204 234530
rect 195152 234466 195204 234472
rect 195256 214713 195284 240042
rect 198016 240009 198044 241590
rect 201604 241505 201632 241590
rect 201590 241496 201646 241505
rect 201590 241431 201646 241440
rect 198002 240000 198058 240009
rect 198002 239935 198058 239944
rect 197360 239488 197412 239494
rect 197360 239430 197412 239436
rect 195980 237448 196032 237454
rect 195980 237390 196032 237396
rect 195242 214704 195298 214713
rect 195242 214639 195298 214648
rect 195992 174554 196020 237390
rect 197372 235822 197400 239430
rect 197360 235816 197412 235822
rect 196622 235784 196678 235793
rect 197360 235758 197412 235764
rect 196622 235719 196678 235728
rect 195980 174548 196032 174554
rect 195980 174490 196032 174496
rect 195244 173188 195296 173194
rect 195244 173130 195296 173136
rect 195256 158846 195284 173130
rect 195978 163432 196034 163441
rect 195978 163367 196034 163376
rect 195244 158840 195296 158846
rect 195244 158782 195296 158788
rect 195060 147008 195112 147014
rect 195060 146950 195112 146956
rect 195072 140978 195100 146950
rect 195072 140950 195454 140978
rect 195992 140964 196020 163367
rect 196072 148436 196124 148442
rect 196072 148378 196124 148384
rect 196084 140978 196112 148378
rect 196636 142225 196664 235719
rect 197358 181384 197414 181393
rect 197358 181319 197414 181328
rect 196716 160200 196768 160206
rect 196716 160142 196768 160148
rect 196728 146266 196756 160142
rect 196716 146260 196768 146266
rect 196716 146202 196768 146208
rect 196622 142216 196678 142225
rect 196622 142151 196678 142160
rect 196084 140950 196558 140978
rect 194784 140480 194836 140486
rect 194784 140422 194836 140428
rect 196636 140434 196664 142151
rect 197372 140978 197400 181319
rect 198016 177410 198044 239935
rect 201880 236026 201908 241590
rect 205192 241398 205220 241604
rect 208412 241590 208518 241618
rect 208412 241505 208440 241590
rect 208398 241496 208454 241505
rect 208398 241431 208454 241440
rect 205180 241392 205232 241398
rect 205180 241334 205232 241340
rect 204258 240136 204314 240145
rect 204258 240071 204314 240080
rect 204272 239465 204300 240071
rect 204258 239456 204314 239465
rect 204258 239391 204314 239400
rect 202234 236872 202290 236881
rect 202234 236807 202290 236816
rect 200764 236020 200816 236026
rect 200764 235962 200816 235968
rect 201868 236020 201920 236026
rect 201868 235962 201920 235968
rect 198646 228440 198702 228449
rect 198646 228375 198702 228384
rect 198094 214568 198150 214577
rect 198094 214503 198150 214512
rect 198004 177404 198056 177410
rect 198004 177346 198056 177352
rect 198108 161673 198136 214503
rect 198094 161664 198150 161673
rect 198094 161599 198150 161608
rect 197452 155984 197504 155990
rect 197452 155926 197504 155932
rect 197464 151814 197492 155926
rect 197464 151786 197952 151814
rect 197924 140978 197952 151786
rect 198660 143177 198688 228375
rect 198738 228304 198794 228313
rect 198738 228239 198794 228248
rect 198646 143168 198702 143177
rect 198646 143103 198702 143112
rect 198752 140978 198780 228239
rect 200776 186998 200804 235962
rect 202248 235793 202276 236807
rect 202234 235784 202290 235793
rect 202234 235719 202290 235728
rect 202786 235784 202842 235793
rect 202786 235719 202842 235728
rect 200854 211984 200910 211993
rect 200854 211919 200910 211928
rect 200764 186992 200816 186998
rect 200764 186934 200816 186940
rect 200120 166388 200172 166394
rect 200120 166330 200172 166336
rect 199382 161664 199438 161673
rect 199382 161599 199438 161608
rect 199396 161566 199424 161599
rect 199384 161560 199436 161566
rect 199384 161502 199436 161508
rect 199200 146260 199252 146266
rect 199200 146202 199252 146208
rect 199212 140978 199240 146202
rect 200132 140978 200160 166330
rect 200868 164257 200896 211919
rect 200210 164248 200266 164257
rect 200210 164183 200266 164192
rect 200854 164248 200910 164257
rect 200854 164183 200910 164192
rect 200224 147014 200252 164183
rect 200302 157448 200358 157457
rect 202800 157418 202828 235719
rect 203522 184240 203578 184249
rect 203522 184175 203578 184184
rect 202880 171828 202932 171834
rect 202880 171770 202932 171776
rect 202892 164354 202920 171770
rect 202880 164348 202932 164354
rect 202880 164290 202932 164296
rect 200302 157383 200358 157392
rect 202144 157412 202196 157418
rect 200316 153105 200344 157383
rect 202144 157354 202196 157360
rect 202788 157412 202840 157418
rect 202788 157354 202840 157360
rect 200302 153096 200358 153105
rect 200302 153031 200358 153040
rect 200212 147008 200264 147014
rect 200212 146950 200264 146956
rect 200316 140978 200344 153031
rect 201590 152552 201646 152561
rect 201590 152487 201646 152496
rect 200948 147008 201000 147014
rect 200948 146950 201000 146956
rect 200960 140978 200988 146950
rect 201604 140978 201632 152487
rect 202050 152416 202106 152425
rect 202050 152351 202106 152360
rect 202064 151842 202092 152351
rect 202052 151836 202104 151842
rect 202052 151778 202104 151784
rect 202156 144265 202184 157354
rect 202892 151814 202920 164290
rect 203536 159361 203564 184175
rect 204272 175370 204300 239391
rect 205192 235278 205220 241334
rect 206284 236700 206336 236706
rect 206284 236642 206336 236648
rect 205180 235272 205232 235278
rect 205180 235214 205232 235220
rect 206296 181490 206324 236642
rect 206374 229120 206430 229129
rect 206374 229055 206430 229064
rect 206388 213246 206416 229055
rect 206376 213240 206428 213246
rect 206376 213182 206428 213188
rect 206284 181484 206336 181490
rect 206284 181426 206336 181432
rect 204260 175364 204312 175370
rect 204260 175306 204312 175312
rect 204904 175364 204956 175370
rect 204904 175306 204956 175312
rect 203522 159352 203578 159361
rect 203522 159287 203578 159296
rect 202892 151786 203472 151814
rect 202142 144256 202198 144265
rect 202142 144191 202198 144200
rect 203156 141500 203208 141506
rect 203156 141442 203208 141448
rect 202604 141432 202656 141438
rect 202604 141374 202656 141380
rect 197372 140950 197846 140978
rect 197924 140950 198398 140978
rect 198752 140950 198950 140978
rect 199212 140950 199686 140978
rect 200132 140950 200238 140978
rect 200316 140950 200790 140978
rect 200960 140950 201342 140978
rect 201604 140950 202078 140978
rect 202616 140964 202644 141374
rect 203168 140842 203196 141442
rect 203444 140978 203472 151786
rect 204258 151056 204314 151065
rect 204258 150991 204314 151000
rect 204272 140978 204300 150991
rect 204916 142186 204944 175306
rect 206388 173194 206416 213182
rect 207662 206272 207718 206281
rect 207662 206207 207718 206216
rect 207676 175273 207704 206207
rect 207018 175264 207074 175273
rect 207018 175199 207074 175208
rect 207662 175264 207718 175273
rect 207662 175199 207718 175208
rect 207032 174049 207060 175199
rect 207018 174040 207074 174049
rect 207018 173975 207074 173984
rect 206376 173188 206428 173194
rect 206376 173130 206428 173136
rect 204996 169040 205048 169046
rect 204996 168982 205048 168988
rect 205008 151814 205036 168982
rect 206284 156732 206336 156738
rect 206284 156674 206336 156680
rect 205008 151786 205220 151814
rect 205192 147694 205220 151786
rect 205180 147688 205232 147694
rect 205180 147630 205232 147636
rect 204994 142216 205050 142225
rect 204904 142180 204956 142186
rect 204994 142151 205050 142160
rect 204904 142122 204956 142128
rect 203444 140950 203918 140978
rect 204272 140950 204470 140978
rect 205008 140964 205036 142151
rect 205192 140978 205220 147630
rect 206296 143449 206324 156674
rect 206468 145036 206520 145042
rect 206468 144978 206520 144984
rect 206282 143440 206338 143449
rect 206282 143375 206338 143384
rect 206480 143313 206508 144978
rect 206834 143440 206890 143449
rect 206834 143375 206890 143384
rect 206466 143304 206522 143313
rect 206466 143239 206522 143248
rect 206480 140978 206508 143239
rect 205192 140950 205574 140978
rect 206310 140950 206508 140978
rect 206848 140964 206876 143375
rect 207032 140978 207060 173975
rect 208412 158030 208440 241431
rect 209044 240168 209096 240174
rect 209044 240110 209096 240116
rect 209778 240136 209834 240145
rect 209056 234530 209084 240110
rect 209778 240071 209834 240080
rect 209792 236706 209820 240071
rect 211908 239426 211936 241604
rect 215220 241534 215248 241604
rect 218546 241590 218744 241618
rect 214012 241528 214064 241534
rect 215208 241528 215260 241534
rect 214012 241470 214064 241476
rect 215206 241496 215208 241505
rect 218624 241505 218652 241590
rect 215260 241496 215262 241505
rect 211896 239420 211948 239426
rect 211896 239362 211948 239368
rect 209780 236700 209832 236706
rect 209780 236642 209832 236648
rect 209044 234524 209096 234530
rect 209044 234466 209096 234472
rect 208400 158024 208452 158030
rect 208400 157966 208452 157972
rect 208492 150408 208544 150414
rect 208492 150350 208544 150356
rect 208122 144120 208178 144129
rect 208122 144055 208178 144064
rect 208136 141409 208164 144055
rect 208122 141400 208178 141409
rect 208122 141335 208178 141344
rect 207032 140950 207414 140978
rect 208136 140964 208164 141335
rect 208504 140978 208532 150350
rect 209056 143857 209084 234466
rect 213184 225616 213236 225622
rect 213184 225558 213236 225564
rect 211158 221640 211214 221649
rect 211158 221575 211214 221584
rect 211172 219337 211200 221575
rect 211158 219328 211214 219337
rect 211158 219263 211214 219272
rect 212446 219328 212502 219337
rect 212446 219263 212502 219272
rect 210424 171148 210476 171154
rect 210424 171090 210476 171096
rect 211160 171148 211212 171154
rect 211160 171090 211212 171096
rect 210436 158710 210464 171090
rect 211172 168366 211200 171090
rect 211160 168360 211212 168366
rect 211160 168302 211212 168308
rect 210424 158704 210476 158710
rect 210424 158646 210476 158652
rect 210436 157486 210464 158646
rect 209780 157480 209832 157486
rect 209780 157422 209832 157428
rect 210424 157480 210476 157486
rect 210424 157422 210476 157428
rect 209134 156088 209190 156097
rect 209134 156023 209190 156032
rect 209148 150414 209176 156023
rect 209226 154592 209282 154601
rect 209226 154527 209282 154536
rect 209240 151745 209268 154527
rect 209792 151814 209820 157422
rect 211172 151814 211200 168302
rect 212460 155961 212488 219263
rect 213196 219201 213224 225558
rect 213920 224256 213972 224262
rect 213920 224198 213972 224204
rect 213182 219192 213238 219201
rect 213182 219127 213238 219136
rect 213196 218113 213224 219127
rect 213182 218104 213238 218113
rect 213182 218039 213238 218048
rect 213184 185632 213236 185638
rect 213184 185574 213236 185580
rect 213196 175953 213224 185574
rect 212630 175944 212686 175953
rect 212630 175879 212686 175888
rect 213182 175944 213238 175953
rect 213182 175879 213238 175888
rect 211802 155952 211858 155961
rect 211802 155887 211858 155896
rect 212446 155952 212502 155961
rect 212446 155887 212502 155896
rect 211816 154601 211844 155887
rect 211802 154592 211858 154601
rect 211802 154527 211858 154536
rect 209792 151786 210740 151814
rect 211172 151786 211752 151814
rect 209226 151736 209282 151745
rect 209226 151671 209282 151680
rect 209136 150408 209188 150414
rect 209136 150350 209188 150356
rect 209042 143848 209098 143857
rect 209042 143783 209098 143792
rect 209240 142154 209268 151671
rect 210054 146976 210110 146985
rect 210054 146911 210110 146920
rect 208872 142126 209268 142154
rect 209780 142180 209832 142186
rect 208872 140978 208900 142126
rect 209780 142122 209832 142128
rect 209792 140978 209820 142122
rect 209962 140992 210018 141001
rect 208504 140950 208702 140978
rect 208872 140950 209254 140978
rect 209792 140964 209962 140978
rect 209806 140950 209962 140964
rect 210068 140978 210096 146911
rect 210712 140978 210740 151786
rect 211158 149152 211214 149161
rect 211158 149087 211214 149096
rect 211172 142154 211200 149087
rect 211250 143712 211306 143721
rect 211250 143647 211306 143656
rect 211264 143614 211292 143647
rect 211252 143608 211304 143614
rect 211252 143550 211304 143556
rect 211724 142154 211752 151786
rect 211816 148374 211844 154527
rect 212446 149152 212502 149161
rect 212446 149087 212502 149096
rect 212460 149054 212488 149087
rect 212448 149048 212500 149054
rect 212448 148990 212500 148996
rect 211804 148368 211856 148374
rect 211804 148310 211856 148316
rect 212644 143449 212672 175879
rect 213932 172553 213960 224198
rect 213918 172544 213974 172553
rect 213918 172479 213974 172488
rect 213184 166320 213236 166326
rect 213184 166262 213236 166268
rect 213196 154562 213224 166262
rect 213276 160744 213328 160750
rect 213276 160686 213328 160692
rect 212724 154556 212776 154562
rect 212724 154498 212776 154504
rect 213184 154556 213236 154562
rect 213184 154498 213236 154504
rect 212736 153270 212764 154498
rect 212724 153264 212776 153270
rect 212724 153206 212776 153212
rect 212630 143440 212686 143449
rect 212630 143375 212686 143384
rect 211172 142126 211292 142154
rect 211724 142126 212028 142154
rect 211264 140978 211292 142126
rect 212000 140978 212028 142126
rect 212736 140978 212764 153206
rect 213288 151065 213316 160686
rect 213274 151056 213330 151065
rect 213274 150991 213330 151000
rect 213458 143440 213514 143449
rect 213458 143375 213514 143384
rect 210068 140950 210542 140978
rect 210712 140950 211094 140978
rect 211264 140950 211646 140978
rect 212000 140950 212382 140978
rect 212736 140950 212934 140978
rect 209962 140927 210018 140936
rect 203168 140828 203472 140842
rect 203182 140826 203472 140828
rect 203182 140820 203484 140826
rect 203182 140814 203432 140820
rect 203432 140762 203484 140768
rect 213472 140570 213500 143375
rect 213932 140842 213960 172479
rect 214024 150550 214052 241470
rect 215206 241431 215262 241440
rect 218610 241496 218666 241505
rect 218610 241431 218666 241440
rect 215220 241405 215248 241431
rect 218716 239737 218744 241590
rect 221568 241590 221858 241618
rect 224972 241590 225552 241618
rect 220084 241528 220136 241534
rect 221568 241505 221596 241590
rect 220084 241470 220136 241476
rect 220910 241496 220966 241505
rect 218702 239728 218758 239737
rect 218702 239663 218758 239672
rect 215944 236700 215996 236706
rect 215944 236642 215996 236648
rect 215300 229084 215352 229090
rect 215300 229026 215352 229032
rect 215312 228750 215340 229026
rect 215956 228750 215984 236642
rect 218716 229770 218744 239663
rect 219440 235272 219492 235278
rect 219440 235214 219492 235220
rect 218704 229764 218756 229770
rect 218704 229706 218756 229712
rect 215300 228744 215352 228750
rect 215300 228686 215352 228692
rect 215944 228744 215996 228750
rect 215944 228686 215996 228692
rect 215312 165753 215340 228686
rect 219452 175302 219480 235214
rect 220096 228993 220124 241470
rect 220910 241431 220966 241440
rect 221554 241496 221610 241505
rect 221554 241431 221610 241440
rect 220082 228984 220138 228993
rect 220082 228919 220138 228928
rect 220096 227769 220124 228919
rect 220082 227760 220138 227769
rect 220082 227695 220138 227704
rect 220820 222964 220872 222970
rect 220820 222906 220872 222912
rect 219714 177440 219770 177449
rect 219714 177375 219770 177384
rect 219728 177342 219756 177375
rect 219532 177336 219584 177342
rect 219532 177278 219584 177284
rect 219716 177336 219768 177342
rect 219716 177278 219768 177284
rect 219440 175296 219492 175302
rect 219440 175238 219492 175244
rect 215944 174548 215996 174554
rect 215944 174490 215996 174496
rect 215298 165744 215354 165753
rect 215298 165679 215354 165688
rect 215312 150906 215340 165679
rect 215390 160168 215446 160177
rect 215390 160103 215446 160112
rect 215404 153202 215432 160103
rect 215392 153196 215444 153202
rect 215392 153138 215444 153144
rect 215404 151814 215432 153138
rect 215404 151786 215892 151814
rect 215312 150878 215616 150906
rect 214012 150544 214064 150550
rect 214012 150486 214064 150492
rect 215484 150544 215536 150550
rect 215484 150486 215536 150492
rect 214024 146946 214052 150486
rect 214012 146940 214064 146946
rect 214012 146882 214064 146888
rect 215496 140978 215524 150486
rect 215326 140950 215524 140978
rect 215588 140978 215616 150878
rect 215864 142154 215892 151786
rect 215956 150550 215984 174490
rect 218060 166320 218112 166326
rect 218060 166262 218112 166268
rect 218072 162926 218100 166262
rect 218060 162920 218112 162926
rect 218060 162862 218112 162868
rect 216680 152584 216732 152590
rect 216680 152526 216732 152532
rect 215944 150544 215996 150550
rect 215944 150486 215996 150492
rect 215864 142126 216260 142154
rect 216232 140978 216260 142126
rect 216692 140978 216720 152526
rect 218072 151814 218100 162862
rect 218702 152688 218758 152697
rect 218702 152623 218758 152632
rect 218072 151786 218560 151814
rect 217230 145072 217286 145081
rect 217230 145007 217286 145016
rect 217244 140978 217272 145007
rect 218244 142996 218296 143002
rect 218244 142938 218296 142944
rect 218256 142186 218284 142938
rect 218244 142180 218296 142186
rect 218244 142122 218296 142128
rect 215588 140950 215878 140978
rect 216232 140950 216614 140978
rect 216692 140950 217166 140978
rect 217244 140950 217718 140978
rect 218256 140964 218284 142122
rect 218532 140978 218560 151786
rect 218716 143002 218744 152623
rect 219544 151814 219572 177278
rect 220084 175296 220136 175302
rect 220084 175238 220136 175244
rect 219452 151786 219572 151814
rect 218704 142996 218756 143002
rect 218704 142938 218756 142944
rect 219452 142225 219480 151786
rect 220096 143614 220124 175238
rect 220832 168473 220860 222906
rect 220924 195974 220952 241431
rect 222290 230344 222346 230353
rect 222290 230279 222346 230288
rect 222200 229764 222252 229770
rect 222200 229706 222252 229712
rect 222106 223000 222162 223009
rect 222106 222935 222108 222944
rect 222160 222935 222162 222944
rect 222108 222906 222160 222912
rect 220912 195968 220964 195974
rect 220912 195910 220964 195916
rect 221832 195968 221884 195974
rect 221832 195910 221884 195916
rect 221844 191826 221872 195910
rect 221832 191820 221884 191826
rect 221832 191762 221884 191768
rect 222212 173942 222240 229706
rect 222304 221513 222332 230279
rect 222290 221504 222346 221513
rect 222290 221439 222346 221448
rect 222844 221468 222896 221474
rect 222844 221410 222896 221416
rect 222200 173936 222252 173942
rect 222200 173878 222252 173884
rect 222856 169833 222884 221410
rect 223762 217288 223818 217297
rect 223762 217223 223818 217232
rect 223580 197328 223632 197334
rect 223580 197270 223632 197276
rect 223592 196722 223620 197270
rect 223580 196716 223632 196722
rect 223580 196658 223632 196664
rect 222936 173936 222988 173942
rect 222936 173878 222988 173884
rect 222198 169824 222254 169833
rect 222198 169759 222254 169768
rect 222842 169824 222898 169833
rect 222842 169759 222898 169768
rect 220818 168464 220874 168473
rect 220818 168399 220874 168408
rect 220832 156670 220860 168399
rect 221004 163532 221056 163538
rect 221004 163474 221056 163480
rect 220820 156664 220872 156670
rect 220740 156612 220820 156618
rect 220740 156606 220872 156612
rect 220740 156590 220860 156606
rect 220084 143608 220136 143614
rect 220084 143550 220136 143556
rect 219532 143132 219584 143138
rect 219532 143074 219584 143080
rect 219438 142216 219494 142225
rect 219438 142151 219494 142160
rect 219452 141438 219480 142151
rect 219440 141432 219492 141438
rect 219440 141374 219492 141380
rect 218532 140950 219006 140978
rect 219544 140964 219572 143074
rect 220096 140964 220124 143550
rect 220740 143138 220768 156590
rect 220832 156541 220860 156590
rect 220912 150476 220964 150482
rect 220912 150418 220964 150424
rect 220728 143132 220780 143138
rect 220728 143074 220780 143080
rect 220924 140978 220952 150418
rect 220846 140950 220952 140978
rect 221016 140978 221044 163474
rect 221924 142860 221976 142866
rect 221924 142802 221976 142808
rect 221936 142225 221964 142802
rect 221922 142216 221978 142225
rect 221922 142151 221978 142160
rect 221016 140950 221398 140978
rect 221936 140964 221964 142151
rect 222212 140978 222240 169759
rect 222948 142154 222976 173878
rect 223592 167074 223620 196658
rect 223776 171134 223804 217223
rect 224972 211138 225000 241590
rect 225524 241505 225552 241590
rect 225510 241496 225566 241505
rect 225510 241431 225566 241440
rect 228560 239465 228588 241604
rect 229098 240136 229154 240145
rect 229098 240071 229154 240080
rect 228546 239456 228602 239465
rect 228546 239391 228602 239400
rect 228454 236600 228510 236609
rect 228454 236535 228510 236544
rect 228364 233912 228416 233918
rect 228364 233854 228416 233860
rect 227720 215280 227772 215286
rect 227720 215222 227772 215228
rect 227732 214810 227760 215222
rect 227720 214804 227772 214810
rect 227720 214746 227772 214752
rect 224960 211132 225012 211138
rect 224960 211074 225012 211080
rect 224224 209092 224276 209098
rect 224224 209034 224276 209040
rect 224236 196722 224264 209034
rect 224224 196716 224276 196722
rect 224224 196658 224276 196664
rect 223776 171106 224264 171134
rect 223580 167068 223632 167074
rect 223580 167010 223632 167016
rect 223394 143576 223450 143585
rect 223394 143511 223450 143520
rect 223212 142248 223264 142254
rect 223212 142190 223264 142196
rect 223224 142154 223252 142190
rect 222948 142126 223252 142154
rect 222212 140950 222502 140978
rect 223224 140964 223252 142126
rect 214286 140856 214342 140865
rect 213932 140814 214286 140842
rect 214286 140791 214342 140800
rect 214656 140616 214708 140622
rect 213472 140556 213776 140570
rect 214708 140564 214880 140570
rect 214656 140558 214880 140564
rect 213486 140554 213776 140556
rect 213486 140548 213788 140554
rect 213486 140542 213736 140548
rect 214668 140542 214880 140558
rect 213736 140490 213788 140496
rect 214852 140486 214880 140542
rect 214840 140480 214892 140486
rect 196806 140448 196862 140457
rect 196636 140406 196806 140434
rect 196862 140406 197110 140434
rect 223408 140457 223436 143511
rect 223592 140978 223620 167010
rect 223672 158772 223724 158778
rect 223672 158714 223724 158720
rect 223684 147014 223712 158714
rect 224236 157593 224264 171106
rect 224222 157584 224278 157593
rect 224222 157519 224278 157528
rect 223672 147008 223724 147014
rect 223672 146950 223724 146956
rect 224236 142361 224264 157519
rect 224408 153332 224460 153338
rect 224408 153274 224460 153280
rect 224420 151814 224448 153274
rect 224420 151786 224540 151814
rect 224222 142352 224278 142361
rect 224222 142287 224278 142296
rect 224236 142154 224264 142287
rect 224236 142126 224356 142154
rect 223592 140950 223790 140978
rect 224328 140964 224356 142126
rect 224512 140486 224540 151786
rect 224592 147008 224644 147014
rect 224592 146950 224644 146956
rect 224604 140978 224632 146950
rect 224604 140950 224894 140978
rect 224500 140480 224552 140486
rect 214840 140422 214892 140428
rect 223394 140448 223450 140457
rect 196806 140383 196862 140392
rect 224500 140422 224552 140428
rect 223394 140383 223450 140392
rect 193218 104272 193274 104281
rect 193218 104207 193274 104216
rect 193232 103562 193260 104207
rect 193220 103556 193272 103562
rect 193220 103498 193272 103504
rect 193404 94512 193456 94518
rect 193404 94454 193456 94460
rect 193416 93854 193444 94454
rect 193232 93826 193444 93854
rect 193232 85474 193260 93826
rect 211710 93392 211766 93401
rect 211646 93350 211710 93378
rect 211710 93327 211766 93336
rect 224774 93392 224830 93401
rect 224830 93350 224894 93378
rect 224774 93327 224830 93336
rect 193784 93226 194166 93242
rect 193772 93220 194166 93226
rect 193824 93214 194166 93220
rect 193772 93162 193824 93168
rect 205088 93152 205140 93158
rect 205088 93094 205140 93100
rect 201590 92848 201646 92857
rect 193324 92806 193614 92834
rect 193220 85468 193272 85474
rect 193220 85410 193272 85416
rect 193324 75857 193352 92806
rect 194704 88602 194732 92820
rect 194796 92806 195270 92834
rect 194692 88596 194744 88602
rect 194692 88538 194744 88544
rect 194796 88482 194824 92806
rect 194612 88454 194824 88482
rect 193310 75848 193366 75857
rect 193310 75783 193366 75792
rect 193862 75848 193918 75857
rect 193862 75783 193918 75792
rect 193128 68332 193180 68338
rect 193128 68274 193180 68280
rect 193876 64802 193904 75783
rect 194612 66201 194640 88454
rect 194692 88392 194744 88398
rect 194692 88334 194744 88340
rect 194704 70378 194732 88334
rect 195992 71398 196020 92820
rect 196162 92712 196218 92721
rect 196162 92647 196218 92656
rect 196176 73166 196204 92647
rect 196544 92449 196572 92820
rect 196530 92440 196586 92449
rect 196530 92375 196586 92384
rect 197096 86601 197124 92820
rect 197372 92806 197662 92834
rect 197832 92806 198398 92834
rect 198950 92806 199332 92834
rect 197372 92585 197400 92806
rect 197358 92576 197414 92585
rect 197358 92511 197414 92520
rect 197082 86592 197138 86601
rect 197082 86527 197138 86536
rect 196164 73160 196216 73166
rect 196164 73102 196216 73108
rect 195980 71392 196032 71398
rect 195980 71334 196032 71340
rect 194692 70372 194744 70378
rect 194692 70314 194744 70320
rect 194704 69970 194732 70314
rect 194692 69964 194744 69970
rect 194692 69906 194744 69912
rect 195336 69964 195388 69970
rect 195336 69906 195388 69912
rect 194598 66192 194654 66201
rect 194598 66127 194654 66136
rect 195242 66192 195298 66201
rect 195242 66127 195298 66136
rect 193864 64796 193916 64802
rect 193864 64738 193916 64744
rect 193876 36582 193904 64738
rect 195256 57934 195284 66127
rect 195348 64802 195376 69906
rect 196176 67590 196204 73102
rect 196624 71732 196676 71738
rect 196624 71674 196676 71680
rect 196636 71398 196664 71674
rect 196624 71392 196676 71398
rect 196624 71334 196676 71340
rect 196164 67584 196216 67590
rect 196164 67526 196216 67532
rect 195336 64796 195388 64802
rect 195336 64738 195388 64744
rect 195244 57928 195296 57934
rect 195244 57870 195296 57876
rect 193864 36576 193916 36582
rect 193864 36518 193916 36524
rect 192576 28280 192628 28286
rect 192576 28222 192628 28228
rect 191748 21412 191800 21418
rect 191748 21354 191800 21360
rect 184848 15904 184900 15910
rect 184848 15846 184900 15852
rect 181536 13116 181588 13122
rect 181536 13058 181588 13064
rect 195256 11762 195284 57870
rect 196636 56574 196664 71334
rect 196624 56568 196676 56574
rect 196624 56510 196676 56516
rect 195244 11756 195296 11762
rect 195244 11698 195296 11704
rect 196636 8974 196664 56510
rect 197372 31074 197400 92511
rect 197832 84194 197860 92806
rect 198738 92576 198794 92585
rect 198738 92511 198794 92520
rect 197464 84166 197860 84194
rect 197464 78577 197492 84166
rect 198752 80102 198780 92511
rect 199304 92449 199332 92806
rect 199488 92585 199516 92820
rect 200132 92806 200238 92834
rect 199474 92576 199530 92585
rect 199474 92511 199530 92520
rect 199290 92440 199346 92449
rect 199290 92375 199346 92384
rect 199304 84194 199332 92375
rect 199304 84166 199424 84194
rect 198740 80096 198792 80102
rect 198740 80038 198792 80044
rect 197450 78568 197506 78577
rect 197450 78503 197506 78512
rect 198752 75886 198780 80038
rect 198740 75880 198792 75886
rect 198740 75822 198792 75828
rect 199396 60722 199424 84166
rect 199384 60716 199436 60722
rect 199384 60658 199436 60664
rect 199396 42090 199424 60658
rect 200132 59362 200160 92806
rect 200776 86737 200804 92820
rect 200762 86728 200818 86737
rect 200762 86663 200818 86672
rect 201328 85377 201356 92820
rect 201646 92820 201894 92834
rect 201646 92806 201908 92820
rect 201590 92783 201646 92792
rect 201880 90273 201908 92806
rect 202616 92313 202644 92820
rect 203182 92806 203564 92834
rect 202602 92304 202658 92313
rect 202602 92239 202658 92248
rect 203536 90545 203564 92806
rect 203522 90536 203578 90545
rect 203522 90471 203578 90480
rect 201866 90264 201922 90273
rect 201866 90199 201922 90208
rect 202786 90264 202842 90273
rect 202786 90199 202842 90208
rect 200394 85368 200450 85377
rect 200394 85303 200450 85312
rect 201314 85368 201370 85377
rect 201314 85303 201370 85312
rect 200408 82142 200436 85303
rect 200396 82136 200448 82142
rect 200396 82078 200448 82084
rect 200120 59356 200172 59362
rect 200120 59298 200172 59304
rect 201408 59356 201460 59362
rect 201408 59298 201460 59304
rect 201420 56574 201448 59298
rect 201408 56568 201460 56574
rect 201408 56510 201460 56516
rect 199384 42084 199436 42090
rect 199384 42026 199436 42032
rect 197360 31068 197412 31074
rect 197360 31010 197412 31016
rect 202800 17270 202828 90199
rect 203536 79665 203564 90471
rect 203720 90409 203748 92820
rect 204456 90681 204484 92820
rect 204442 90672 204498 90681
rect 204442 90607 204498 90616
rect 203706 90400 203762 90409
rect 203706 90335 203762 90344
rect 203720 88262 203748 90335
rect 204350 90264 204406 90273
rect 204350 90199 204406 90208
rect 203708 88256 203760 88262
rect 203708 88198 203760 88204
rect 204166 80064 204222 80073
rect 204166 79999 204222 80008
rect 204180 79665 204208 79999
rect 204364 79801 204392 90199
rect 204456 86873 204484 90607
rect 205008 89622 205036 92820
rect 205100 89622 205128 93094
rect 222658 92984 222714 92993
rect 222502 92956 222658 92970
rect 222488 92942 222658 92956
rect 205454 92848 205510 92857
rect 208398 92848 208454 92857
rect 205510 92820 205574 92834
rect 205510 92806 205588 92820
rect 205454 92783 205510 92792
rect 205560 90273 205588 92806
rect 205546 90264 205602 90273
rect 205546 90199 205602 90208
rect 204996 89616 205048 89622
rect 204996 89558 205048 89564
rect 205088 89616 205140 89622
rect 206112 89593 206140 92820
rect 206204 92806 206862 92834
rect 205088 89558 205140 89564
rect 206098 89584 206154 89593
rect 206098 89519 206154 89528
rect 204996 88256 205048 88262
rect 204996 88198 205048 88204
rect 205008 88097 205036 88198
rect 204994 88088 205050 88097
rect 204994 88023 205050 88032
rect 204442 86864 204498 86873
rect 204442 86799 204498 86808
rect 206204 84194 206232 92806
rect 207400 88262 207428 92820
rect 207492 92806 207966 92834
rect 206284 88256 206336 88262
rect 206284 88198 206336 88204
rect 207388 88256 207440 88262
rect 207388 88198 207440 88204
rect 205652 84182 206232 84194
rect 205640 84176 206232 84182
rect 205692 84166 206232 84176
rect 205640 84118 205692 84124
rect 204350 79792 204406 79801
rect 204350 79727 204406 79736
rect 203522 79656 203578 79665
rect 203522 79591 203578 79600
rect 204166 79656 204222 79665
rect 204166 79591 204222 79600
rect 204180 25566 204208 79591
rect 204364 79529 204392 79727
rect 204350 79520 204406 79529
rect 204350 79455 204406 79464
rect 204902 79520 204958 79529
rect 204902 79455 204958 79464
rect 204916 35222 204944 79455
rect 206296 57866 206324 88198
rect 207492 84194 207520 92806
rect 210054 92848 210110 92857
rect 208454 92820 208702 92834
rect 208454 92806 208716 92820
rect 208398 92783 208454 92792
rect 208688 90273 208716 92806
rect 208674 90264 208730 90273
rect 208674 90199 208730 90208
rect 209240 89729 209268 92820
rect 209686 90264 209742 90273
rect 209686 90199 209742 90208
rect 209226 89720 209282 89729
rect 209226 89655 209282 89664
rect 206928 84176 206980 84182
rect 206928 84118 206980 84124
rect 207032 84166 207520 84194
rect 206940 77178 206968 84118
rect 207032 79966 207060 84166
rect 207020 79960 207072 79966
rect 207020 79902 207072 79908
rect 207032 79558 207060 79902
rect 207020 79552 207072 79558
rect 207020 79494 207072 79500
rect 207664 79552 207716 79558
rect 207664 79494 207716 79500
rect 206928 77172 206980 77178
rect 206928 77114 206980 77120
rect 206284 57860 206336 57866
rect 206284 57802 206336 57808
rect 204904 35216 204956 35222
rect 204904 35158 204956 35164
rect 204168 25560 204220 25566
rect 204168 25502 204220 25508
rect 206296 24138 206324 57802
rect 206940 57254 206968 77114
rect 206928 57248 206980 57254
rect 206928 57190 206980 57196
rect 207676 51746 207704 79494
rect 207664 51740 207716 51746
rect 207664 51682 207716 51688
rect 209700 29646 209728 90199
rect 209792 82793 209820 92820
rect 220266 92848 220322 92857
rect 210110 92806 210358 92834
rect 210054 92783 210110 92792
rect 211080 92410 211108 92820
rect 210424 92404 210476 92410
rect 210424 92346 210476 92352
rect 211068 92404 211120 92410
rect 211068 92346 211120 92352
rect 210436 83502 210464 92346
rect 212184 91905 212212 92820
rect 212552 92806 212934 92834
rect 213288 92806 213486 92834
rect 212170 91896 212226 91905
rect 212170 91831 212226 91840
rect 212184 91050 212212 91831
rect 212172 91044 212224 91050
rect 212172 90986 212224 90992
rect 210424 83496 210476 83502
rect 210424 83438 210476 83444
rect 209778 82784 209834 82793
rect 209778 82719 209834 82728
rect 209792 77246 209820 82719
rect 209780 77240 209832 77246
rect 209780 77182 209832 77188
rect 212552 74526 212580 92806
rect 213288 91050 213316 92806
rect 213276 91044 213328 91050
rect 213276 90986 213328 90992
rect 213288 79937 213316 90986
rect 214024 88330 214052 92820
rect 214590 92806 214880 92834
rect 214562 91760 214618 91769
rect 214562 91695 214618 91704
rect 214576 89457 214604 91695
rect 214656 89752 214708 89758
rect 214852 89729 214880 92806
rect 214656 89694 214708 89700
rect 214838 89720 214894 89729
rect 214562 89448 214618 89457
rect 214562 89383 214618 89392
rect 214012 88324 214064 88330
rect 214012 88266 214064 88272
rect 214668 84194 214696 89694
rect 214838 89655 214894 89664
rect 215312 85542 215340 92820
rect 215864 90953 215892 92820
rect 216048 92806 216430 92834
rect 217166 92806 217364 92834
rect 216048 92721 216076 92806
rect 216034 92712 216090 92721
rect 216034 92647 216090 92656
rect 215850 90944 215906 90953
rect 215850 90879 215906 90888
rect 215300 85536 215352 85542
rect 215300 85478 215352 85484
rect 216048 85474 216076 92647
rect 217336 85542 217364 92806
rect 217704 89690 217732 92820
rect 217692 89684 217744 89690
rect 217692 89626 217744 89632
rect 218256 86970 218284 92820
rect 218808 89758 218836 92820
rect 219544 90001 219572 92820
rect 219636 92806 220266 92834
rect 219530 89992 219586 90001
rect 219530 89927 219586 89936
rect 219636 89842 219664 92806
rect 220266 92783 220322 92792
rect 219714 90944 219770 90953
rect 219714 90879 219770 90888
rect 219452 89814 219664 89842
rect 218796 89752 218848 89758
rect 218796 89694 218848 89700
rect 218244 86964 218296 86970
rect 218244 86906 218296 86912
rect 217324 85536 217376 85542
rect 217324 85478 217376 85484
rect 216036 85468 216088 85474
rect 216036 85410 216088 85416
rect 214576 84166 214696 84194
rect 214576 81326 214604 84166
rect 214564 81320 214616 81326
rect 214564 81262 214616 81268
rect 213274 79928 213330 79937
rect 213274 79863 213330 79872
rect 212540 74520 212592 74526
rect 212540 74462 212592 74468
rect 212552 73166 212580 74462
rect 212540 73160 212592 73166
rect 212540 73102 212592 73108
rect 213288 57254 213316 79863
rect 213184 57248 213236 57254
rect 213184 57190 213236 57196
rect 213276 57248 213328 57254
rect 213276 57190 213328 57196
rect 209688 29640 209740 29646
rect 209688 29582 209740 29588
rect 206284 24132 206336 24138
rect 206284 24074 206336 24080
rect 202788 17264 202840 17270
rect 202788 17206 202840 17212
rect 196624 8968 196676 8974
rect 196624 8910 196676 8916
rect 213196 3466 213224 57190
rect 214576 22778 214604 81262
rect 215944 73840 215996 73846
rect 215944 73782 215996 73788
rect 214564 22772 214616 22778
rect 214564 22714 214616 22720
rect 215956 17338 215984 73782
rect 216048 69698 216076 85410
rect 216036 69692 216088 69698
rect 216036 69634 216088 69640
rect 217336 62082 217364 85478
rect 219452 84153 219480 89814
rect 219438 84144 219494 84153
rect 219438 84079 219494 84088
rect 219728 66230 219756 90879
rect 220082 89992 220138 90001
rect 220082 89927 220138 89936
rect 220096 77217 220124 89927
rect 220648 89593 220676 92820
rect 220728 91112 220780 91118
rect 220728 91054 220780 91060
rect 220740 90953 220768 91054
rect 220726 90944 220782 90953
rect 220726 90879 220782 90888
rect 221384 89690 221412 92820
rect 221372 89684 221424 89690
rect 221372 89626 221424 89632
rect 220634 89584 220690 89593
rect 220634 89519 220690 89528
rect 221936 88233 221964 92820
rect 222488 90302 222516 92942
rect 222658 92919 222714 92928
rect 223946 92848 224002 92857
rect 222580 92806 223054 92834
rect 223790 92820 223946 92834
rect 223776 92806 223946 92820
rect 222476 90296 222528 90302
rect 222476 90238 222528 90244
rect 221922 88224 221978 88233
rect 221922 88159 221978 88168
rect 222580 84194 222608 92806
rect 222844 92540 222896 92546
rect 222844 92482 222896 92488
rect 222212 84166 222608 84194
rect 220082 77208 220138 77217
rect 220082 77143 220138 77152
rect 222212 67522 222240 84166
rect 222856 78606 222884 92482
rect 223776 90846 223804 92806
rect 223946 92783 224002 92792
rect 224328 90953 224356 92820
rect 224972 91118 225000 211074
rect 225144 191820 225196 191826
rect 225144 191762 225196 191768
rect 225052 146940 225104 146946
rect 225052 146882 225104 146888
rect 225064 129577 225092 146882
rect 225050 129568 225106 129577
rect 225050 129503 225106 129512
rect 225050 104952 225106 104961
rect 225050 104887 225106 104896
rect 224960 91112 225012 91118
rect 224960 91054 225012 91060
rect 224314 90944 224370 90953
rect 224314 90879 224370 90888
rect 223764 90840 223816 90846
rect 223764 90782 223816 90788
rect 224868 90840 224920 90846
rect 224868 90782 224920 90788
rect 222844 78600 222896 78606
rect 222844 78542 222896 78548
rect 222200 67516 222252 67522
rect 222200 67458 222252 67464
rect 222844 67516 222896 67522
rect 222844 67458 222896 67464
rect 219716 66224 219768 66230
rect 219716 66166 219768 66172
rect 220084 66224 220136 66230
rect 220084 66166 220136 66172
rect 217324 62076 217376 62082
rect 217324 62018 217376 62024
rect 220096 19990 220124 66166
rect 220084 19984 220136 19990
rect 220084 19926 220136 19932
rect 215944 17332 215996 17338
rect 215944 17274 215996 17280
rect 222856 10334 222884 67458
rect 222844 10328 222896 10334
rect 222844 10270 222896 10276
rect 224880 6186 224908 90782
rect 225064 86902 225092 104887
rect 225156 100745 225184 191762
rect 226432 179444 226484 179450
rect 226432 179386 226484 179392
rect 226338 147112 226394 147121
rect 226338 147047 226394 147056
rect 225604 143676 225656 143682
rect 225604 143618 225656 143624
rect 225616 133210 225644 143618
rect 226352 139913 226380 147047
rect 226338 139904 226394 139913
rect 226338 139839 226394 139848
rect 225604 133204 225656 133210
rect 225604 133146 225656 133152
rect 225616 130937 225644 133146
rect 226340 132388 226392 132394
rect 226340 132330 226392 132336
rect 226352 132025 226380 132330
rect 226338 132016 226394 132025
rect 226338 131951 226394 131960
rect 226340 131096 226392 131102
rect 226340 131038 226392 131044
rect 225602 130928 225658 130937
rect 225602 130863 225658 130872
rect 226352 130121 226380 131038
rect 226338 130112 226394 130121
rect 226338 130047 226394 130056
rect 225326 129296 225382 129305
rect 225326 129231 225382 129240
rect 225340 128926 225368 129231
rect 225328 128920 225380 128926
rect 225328 128862 225380 128868
rect 225234 116784 225290 116793
rect 225234 116719 225290 116728
rect 225142 100736 225198 100745
rect 225142 100671 225198 100680
rect 225156 99482 225184 100671
rect 225144 99476 225196 99482
rect 225144 99418 225196 99424
rect 225052 86896 225104 86902
rect 225052 86838 225104 86844
rect 225156 78674 225184 99418
rect 225248 92546 225276 116719
rect 226444 109721 226472 179386
rect 226708 177404 226760 177410
rect 226708 177346 226760 177352
rect 226524 146940 226576 146946
rect 226524 146882 226576 146888
rect 226536 144974 226564 146882
rect 226524 144968 226576 144974
rect 226524 144910 226576 144916
rect 226536 132841 226564 144910
rect 226616 138712 226668 138718
rect 226616 138654 226668 138660
rect 226628 138281 226656 138654
rect 226614 138272 226670 138281
rect 226614 138207 226670 138216
rect 226616 137284 226668 137290
rect 226616 137226 226668 137232
rect 226628 137193 226656 137226
rect 226614 137184 226670 137193
rect 226614 137119 226670 137128
rect 226616 133748 226668 133754
rect 226616 133690 226668 133696
rect 226628 133657 226656 133690
rect 226614 133648 226670 133657
rect 226614 133583 226670 133592
rect 226522 132832 226578 132841
rect 226522 132767 226578 132776
rect 226616 126948 226668 126954
rect 226616 126890 226668 126896
rect 226524 126880 226576 126886
rect 226524 126822 226576 126828
rect 226536 126585 226564 126822
rect 226522 126576 226578 126585
rect 226522 126511 226578 126520
rect 226628 125769 226656 126890
rect 226614 125760 226670 125769
rect 226614 125695 226670 125704
rect 226616 124160 226668 124166
rect 226616 124102 226668 124108
rect 226628 123049 226656 124102
rect 226614 123040 226670 123049
rect 226614 122975 226670 122984
rect 226616 122800 226668 122806
rect 226616 122742 226668 122748
rect 226628 122233 226656 122742
rect 226614 122224 226670 122233
rect 226614 122159 226670 122168
rect 226616 121440 226668 121446
rect 226616 121382 226668 121388
rect 226628 120329 226656 121382
rect 226614 120320 226670 120329
rect 226614 120255 226670 120264
rect 226616 119672 226668 119678
rect 226616 119614 226668 119620
rect 226628 119513 226656 119614
rect 226614 119504 226670 119513
rect 226614 119439 226670 119448
rect 226616 117972 226668 117978
rect 226616 117914 226668 117920
rect 226628 117609 226656 117914
rect 226614 117600 226670 117609
rect 226614 117535 226670 117544
rect 226616 116000 226668 116006
rect 226614 115968 226616 115977
rect 226668 115968 226670 115977
rect 226614 115903 226670 115912
rect 226524 113892 226576 113898
rect 226524 113834 226576 113840
rect 226536 113257 226564 113834
rect 226522 113248 226578 113257
rect 226522 113183 226578 113192
rect 226720 113174 226748 177346
rect 226798 140448 226854 140457
rect 226798 140383 226854 140392
rect 226812 135250 226840 140383
rect 226800 135244 226852 135250
rect 226800 135186 226852 135192
rect 226812 134745 226840 135186
rect 226798 134736 226854 134745
rect 226798 134671 226854 134680
rect 227076 129736 227128 129742
rect 227076 129678 227128 129684
rect 227088 128489 227116 129678
rect 227074 128480 227130 128489
rect 227074 128415 227130 128424
rect 226800 128308 226852 128314
rect 226800 128250 226852 128256
rect 226812 127401 226840 128250
rect 226798 127392 226854 127401
rect 226798 127327 226854 127336
rect 226800 125588 226852 125594
rect 226800 125530 226852 125536
rect 226812 124681 226840 125530
rect 226798 124672 226854 124681
rect 226798 124607 226854 124616
rect 226798 118416 226854 118425
rect 226798 118351 226854 118360
rect 226812 118046 226840 118351
rect 226800 118040 226852 118046
rect 226800 117982 226852 117988
rect 226984 116680 227036 116686
rect 226984 116622 227036 116628
rect 226616 113144 226668 113150
rect 226720 113146 226840 113174
rect 226616 113086 226668 113092
rect 226628 112169 226656 113086
rect 226614 112160 226670 112169
rect 226614 112095 226670 112104
rect 226708 111784 226760 111790
rect 226708 111726 226760 111732
rect 226720 110537 226748 111726
rect 226706 110528 226762 110537
rect 226706 110463 226762 110472
rect 226430 109712 226486 109721
rect 226430 109647 226486 109656
rect 226616 108996 226668 109002
rect 226616 108938 226668 108944
rect 226628 108633 226656 108938
rect 226614 108624 226670 108633
rect 226614 108559 226670 108568
rect 226708 107636 226760 107642
rect 226708 107578 226760 107584
rect 226720 107001 226748 107578
rect 226706 106992 226762 107001
rect 226706 106927 226762 106936
rect 226706 105904 226762 105913
rect 226706 105839 226762 105848
rect 226720 104922 226748 105839
rect 226708 104916 226760 104922
rect 226708 104858 226760 104864
rect 226522 104272 226578 104281
rect 226522 104207 226578 104216
rect 226536 103562 226564 104207
rect 226524 103556 226576 103562
rect 226524 103498 226576 103504
rect 226614 103456 226670 103465
rect 226614 103391 226670 103400
rect 226628 102202 226656 103391
rect 226616 102196 226668 102202
rect 226616 102138 226668 102144
rect 226430 99648 226486 99657
rect 226430 99583 226486 99592
rect 226444 99414 226472 99583
rect 226432 99408 226484 99414
rect 226432 99350 226484 99356
rect 226430 98832 226486 98841
rect 226430 98767 226486 98776
rect 226340 96620 226392 96626
rect 226340 96562 226392 96568
rect 226352 95305 226380 96562
rect 226338 95296 226394 95305
rect 226338 95231 226394 95240
rect 225236 92540 225288 92546
rect 225236 92482 225288 92488
rect 226340 90296 226392 90302
rect 226340 90238 226392 90244
rect 225144 78668 225196 78674
rect 225144 78610 225196 78616
rect 226352 64870 226380 90238
rect 226444 89457 226472 98767
rect 226708 98048 226760 98054
rect 226706 98016 226708 98025
rect 226760 98016 226762 98025
rect 226706 97951 226762 97960
rect 226522 97200 226578 97209
rect 226522 97135 226578 97144
rect 226536 92449 226564 97135
rect 226812 94489 226840 113146
rect 226996 111353 227024 116622
rect 226982 111344 227038 111353
rect 226982 111279 227038 111288
rect 226984 109744 227036 109750
rect 226984 109686 227036 109692
rect 226996 96121 227024 109686
rect 227444 104168 227496 104174
rect 227444 104110 227496 104116
rect 227456 101561 227484 104110
rect 227442 101552 227498 101561
rect 227442 101487 227498 101496
rect 226982 96112 227038 96121
rect 226982 96047 227038 96056
rect 226892 95940 226944 95946
rect 226892 95882 226944 95888
rect 226798 94480 226854 94489
rect 226798 94415 226854 94424
rect 226812 92478 226840 94415
rect 226904 93673 226932 95882
rect 226890 93664 226946 93673
rect 226890 93599 226946 93608
rect 226800 92472 226852 92478
rect 226522 92440 226578 92449
rect 226800 92414 226852 92420
rect 226522 92375 226578 92384
rect 226430 89448 226486 89457
rect 226430 89383 226486 89392
rect 226812 87650 226840 92414
rect 227732 90001 227760 214746
rect 227812 173188 227864 173194
rect 227812 173130 227864 173136
rect 227824 114073 227852 173130
rect 227904 140480 227956 140486
rect 227904 140422 227956 140428
rect 227916 129742 227944 140422
rect 227904 129736 227956 129742
rect 227904 129678 227956 129684
rect 227996 115320 228048 115326
rect 227996 115262 228048 115268
rect 228008 114889 228036 115262
rect 227994 114880 228050 114889
rect 227994 114815 228050 114824
rect 227810 114064 227866 114073
rect 227810 113999 227866 114008
rect 227824 113218 227852 113999
rect 227812 113212 227864 113218
rect 227812 113154 227864 113160
rect 227904 102808 227956 102814
rect 227904 102750 227956 102756
rect 227916 102377 227944 102750
rect 227902 102368 227958 102377
rect 227902 102303 227958 102312
rect 227718 89992 227774 90001
rect 227718 89927 227774 89936
rect 227732 89049 227760 89927
rect 227718 89040 227774 89049
rect 227718 88975 227774 88984
rect 226800 87644 226852 87650
rect 226800 87586 226852 87592
rect 227916 75886 227944 102303
rect 228008 81433 228036 114815
rect 228376 91050 228404 233854
rect 228468 214810 228496 236535
rect 228456 214804 228508 214810
rect 228456 214746 228508 214752
rect 229112 209001 229140 240071
rect 231872 239494 231900 241604
rect 235198 241590 235488 241618
rect 238510 241590 238708 241618
rect 234618 240136 234674 240145
rect 234618 240071 234674 240080
rect 231860 239488 231912 239494
rect 231860 239430 231912 239436
rect 233882 238776 233938 238785
rect 233882 238711 233938 238720
rect 231766 235240 231822 235249
rect 231766 235175 231822 235184
rect 229834 234016 229890 234025
rect 229834 233951 229890 233960
rect 229848 233209 229876 233951
rect 229834 233200 229890 233209
rect 231780 233170 231808 235175
rect 229834 233135 229890 233144
rect 230480 233164 230532 233170
rect 229848 219434 229876 233135
rect 230480 233106 230532 233112
rect 231768 233164 231820 233170
rect 231768 233106 231820 233112
rect 229756 219406 229876 219434
rect 229098 208992 229154 209001
rect 229098 208927 229154 208936
rect 229098 153232 229154 153241
rect 229098 153167 229154 153176
rect 228456 128920 228508 128926
rect 228456 128862 228508 128868
rect 228468 122126 228496 128862
rect 229112 126954 229140 153167
rect 229190 147928 229246 147937
rect 229190 147863 229246 147872
rect 229204 133754 229232 147863
rect 229192 133748 229244 133754
rect 229192 133690 229244 133696
rect 229100 126948 229152 126954
rect 229100 126890 229152 126896
rect 228456 122120 228508 122126
rect 228456 122062 228508 122068
rect 229756 109002 229784 219406
rect 229836 192500 229888 192506
rect 229836 192442 229888 192448
rect 229848 166394 229876 192442
rect 229836 166388 229888 166394
rect 229836 166330 229888 166336
rect 229836 159384 229888 159390
rect 229836 159326 229888 159332
rect 229848 147937 229876 159326
rect 230492 150521 230520 233106
rect 233896 196654 233924 238711
rect 233884 196648 233936 196654
rect 233884 196590 233936 196596
rect 234528 168360 234580 168366
rect 234528 168302 234580 168308
rect 233240 161560 233292 161566
rect 233240 161502 233292 161508
rect 231858 160304 231914 160313
rect 231858 160239 231914 160248
rect 230572 157412 230624 157418
rect 230572 157354 230624 157360
rect 230478 150512 230534 150521
rect 230478 150447 230534 150456
rect 229834 147928 229890 147937
rect 229834 147863 229890 147872
rect 229834 142216 229890 142225
rect 229834 142151 229890 142160
rect 229848 119406 229876 142151
rect 230492 138718 230520 150447
rect 230480 138712 230532 138718
rect 230480 138654 230532 138660
rect 230584 119678 230612 157354
rect 230664 146328 230716 146334
rect 230664 146270 230716 146276
rect 230572 119672 230624 119678
rect 230572 119614 230624 119620
rect 229836 119400 229888 119406
rect 229836 119342 229888 119348
rect 230480 116000 230532 116006
rect 230480 115942 230532 115948
rect 229836 113212 229888 113218
rect 229836 113154 229888 113160
rect 229744 108996 229796 109002
rect 229744 108938 229796 108944
rect 229744 102128 229796 102134
rect 229744 102070 229796 102076
rect 229100 99408 229152 99414
rect 229100 99350 229152 99356
rect 228364 91044 228416 91050
rect 228364 90986 228416 90992
rect 229112 89622 229140 99350
rect 229100 89616 229152 89622
rect 229100 89558 229152 89564
rect 229756 82822 229784 102070
rect 229744 82816 229796 82822
rect 229744 82758 229796 82764
rect 227994 81424 228050 81433
rect 227994 81359 228050 81368
rect 227904 75880 227956 75886
rect 227904 75822 227956 75828
rect 228364 75880 228416 75886
rect 228364 75822 228416 75828
rect 226340 64864 226392 64870
rect 226340 64806 226392 64812
rect 226352 63578 226380 64806
rect 226340 63572 226392 63578
rect 226340 63514 226392 63520
rect 226984 63572 227036 63578
rect 226984 63514 227036 63520
rect 226996 14482 227024 63514
rect 226984 14476 227036 14482
rect 226984 14418 227036 14424
rect 224868 6180 224920 6186
rect 224868 6122 224920 6128
rect 228376 4894 228404 75822
rect 229848 26926 229876 113154
rect 230388 100020 230440 100026
rect 230388 99962 230440 99968
rect 230400 99414 230428 99962
rect 230388 99408 230440 99414
rect 230388 99350 230440 99356
rect 230492 84017 230520 115942
rect 230676 113898 230704 146270
rect 231872 124166 231900 160239
rect 231950 143712 232006 143721
rect 231950 143647 232006 143656
rect 231964 125594 231992 143647
rect 233252 137290 233280 161502
rect 234540 145586 234568 168302
rect 234528 145580 234580 145586
rect 234528 145522 234580 145528
rect 233240 137284 233292 137290
rect 233240 137226 233292 137232
rect 233884 137284 233936 137290
rect 233884 137226 233936 137232
rect 231952 125588 232004 125594
rect 231952 125530 232004 125536
rect 231860 124160 231912 124166
rect 231860 124102 231912 124108
rect 233896 120766 233924 137226
rect 233884 120760 233936 120766
rect 233884 120702 233936 120708
rect 231768 116612 231820 116618
rect 231768 116554 231820 116560
rect 231780 116006 231808 116554
rect 231768 116000 231820 116006
rect 231768 115942 231820 115948
rect 230664 113892 230716 113898
rect 230664 113834 230716 113840
rect 231860 103556 231912 103562
rect 231860 103498 231912 103504
rect 230478 84008 230534 84017
rect 230478 83943 230534 83952
rect 231872 73098 231900 103498
rect 231860 73092 231912 73098
rect 231860 73034 231912 73040
rect 234632 72457 234660 240071
rect 235276 185638 235304 241590
rect 235460 241505 235488 241590
rect 238680 241505 238708 241590
rect 241532 241590 242296 241618
rect 235446 241496 235502 241505
rect 235446 241431 235502 241440
rect 238666 241496 238722 241505
rect 238666 241431 238722 241440
rect 238758 241088 238814 241097
rect 238758 241023 238814 241032
rect 238772 235929 238800 241023
rect 238852 238060 238904 238066
rect 238852 238002 238904 238008
rect 238758 235920 238814 235929
rect 238758 235855 238814 235864
rect 238864 229094 238892 238002
rect 240232 231124 240284 231130
rect 240232 231066 240284 231072
rect 238772 229066 238892 229094
rect 237380 227112 237432 227118
rect 237378 227080 237380 227089
rect 237432 227080 237434 227089
rect 237434 227038 237512 227066
rect 237378 227015 237434 227024
rect 236092 225684 236144 225690
rect 236092 225626 236144 225632
rect 236104 220794 236132 225626
rect 237380 222896 237432 222902
rect 237378 222864 237380 222873
rect 237432 222864 237434 222873
rect 237378 222799 237434 222808
rect 236092 220788 236144 220794
rect 236092 220730 236144 220736
rect 236000 188352 236052 188358
rect 236000 188294 236052 188300
rect 235264 185632 235316 185638
rect 235264 185574 235316 185580
rect 235264 145036 235316 145042
rect 235264 144978 235316 144984
rect 235276 132462 235304 144978
rect 235264 132456 235316 132462
rect 235264 132398 235316 132404
rect 236012 118046 236040 188294
rect 236104 161537 236132 220730
rect 237484 219434 237512 227038
rect 238666 222864 238722 222873
rect 238666 222799 238722 222808
rect 237392 219406 237512 219434
rect 236090 161528 236146 161537
rect 236090 161463 236146 161472
rect 236104 138553 236132 161463
rect 237392 154465 237420 219406
rect 238680 178702 238708 222799
rect 238024 178696 238076 178702
rect 238024 178638 238076 178644
rect 238668 178696 238720 178702
rect 238668 178638 238720 178644
rect 237472 164280 237524 164286
rect 237472 164222 237524 164228
rect 237378 154456 237434 154465
rect 237378 154391 237434 154400
rect 236642 140992 236698 141001
rect 236642 140927 236698 140936
rect 236090 138544 236146 138553
rect 236090 138479 236146 138488
rect 236000 118040 236052 118046
rect 236000 117982 236052 117988
rect 236012 115258 236040 117982
rect 236000 115252 236052 115258
rect 236000 115194 236052 115200
rect 234618 72448 234674 72457
rect 234618 72383 234674 72392
rect 236656 42090 236684 140927
rect 237484 132494 237512 164222
rect 238036 154737 238064 178638
rect 238022 154728 238078 154737
rect 238022 154663 238078 154672
rect 237562 154456 237618 154465
rect 237562 154391 237618 154400
rect 237576 153377 237604 154391
rect 237562 153368 237618 153377
rect 237562 153303 237618 153312
rect 237392 132466 237512 132494
rect 237392 128314 237420 132466
rect 237380 128308 237432 128314
rect 237380 128250 237432 128256
rect 237392 127634 237420 128250
rect 237380 127628 237432 127634
rect 237380 127570 237432 127576
rect 237576 121446 237604 153303
rect 238036 151814 238064 154663
rect 238772 152425 238800 229066
rect 240046 228440 240102 228449
rect 238852 228404 238904 228410
rect 240046 228375 240048 228384
rect 238852 228346 238904 228352
rect 240100 228375 240102 228384
rect 240048 228346 240100 228352
rect 238864 164393 238892 228346
rect 240244 224913 240272 231066
rect 240230 224904 240286 224913
rect 240230 224839 240286 224848
rect 238850 164384 238906 164393
rect 238850 164319 238906 164328
rect 238758 152416 238814 152425
rect 238758 152351 238814 152360
rect 237668 151786 238064 151814
rect 237668 122806 237696 151786
rect 238024 142248 238076 142254
rect 238024 142190 238076 142196
rect 237656 122800 237708 122806
rect 237656 122742 237708 122748
rect 237564 121440 237616 121446
rect 237564 121382 237616 121388
rect 236736 108316 236788 108322
rect 236736 108258 236788 108264
rect 236748 89690 236776 108258
rect 236736 89684 236788 89690
rect 236736 89626 236788 89632
rect 233884 42084 233936 42090
rect 233884 42026 233936 42032
rect 236644 42084 236696 42090
rect 236644 42026 236696 42032
rect 229836 26920 229888 26926
rect 229836 26862 229888 26868
rect 228364 4888 228416 4894
rect 228364 4830 228416 4836
rect 233896 4078 233924 42026
rect 238036 4826 238064 142190
rect 238116 122188 238168 122194
rect 238116 122130 238168 122136
rect 238128 78441 238156 122130
rect 238772 116686 238800 152351
rect 238864 132394 238892 164319
rect 240140 149728 240192 149734
rect 240140 149670 240192 149676
rect 238852 132388 238904 132394
rect 238852 132330 238904 132336
rect 240152 117978 240180 149670
rect 240244 149433 240272 224839
rect 240784 224324 240836 224330
rect 240784 224266 240836 224272
rect 240796 218006 240824 224266
rect 240784 218000 240836 218006
rect 240784 217942 240836 217948
rect 240796 194614 240824 217942
rect 241532 202842 241560 241590
rect 242268 241505 242296 241590
rect 242254 241496 242310 241505
rect 242254 241431 242310 241440
rect 244280 240848 244332 240854
rect 244278 240816 244280 240825
rect 244332 240816 244334 240825
rect 244278 240751 244334 240760
rect 241610 240136 241666 240145
rect 241610 240071 241666 240080
rect 241520 202836 241572 202842
rect 241520 202778 241572 202784
rect 240784 194608 240836 194614
rect 240784 194550 240836 194556
rect 240796 190454 240824 194550
rect 240796 190426 240916 190454
rect 240784 186992 240836 186998
rect 240784 186934 240836 186940
rect 240796 149734 240824 186934
rect 240784 149728 240836 149734
rect 240784 149670 240836 149676
rect 240230 149424 240286 149433
rect 240230 149359 240286 149368
rect 240244 120329 240272 149359
rect 240230 120320 240286 120329
rect 240230 120255 240286 120264
rect 240140 117972 240192 117978
rect 240140 117914 240192 117920
rect 240784 117972 240836 117978
rect 240784 117914 240836 117920
rect 238760 116680 238812 116686
rect 238760 116622 238812 116628
rect 240048 108180 240100 108186
rect 240048 108122 240100 108128
rect 240060 100026 240088 108122
rect 240048 100020 240100 100026
rect 240048 99962 240100 99968
rect 238114 78432 238170 78441
rect 238114 78367 238170 78376
rect 240796 17338 240824 117914
rect 240888 96626 240916 190426
rect 241532 108186 241560 202778
rect 241520 108180 241572 108186
rect 241520 108122 241572 108128
rect 240876 96620 240928 96626
rect 240876 96562 240928 96568
rect 241520 87644 241572 87650
rect 241520 87586 241572 87592
rect 240784 17332 240836 17338
rect 240784 17274 240836 17280
rect 241532 16574 241560 87586
rect 241624 80073 241652 240071
rect 243544 238808 243596 238814
rect 243544 238750 243596 238756
rect 243556 168366 243584 238750
rect 244372 196648 244424 196654
rect 244372 196590 244424 196596
rect 243544 168360 243596 168366
rect 243544 168302 243596 168308
rect 243544 162172 243596 162178
rect 243544 162114 243596 162120
rect 241704 161492 241756 161498
rect 241704 161434 241756 161440
rect 241716 126886 241744 161434
rect 241704 126880 241756 126886
rect 241704 126822 241756 126828
rect 242808 99476 242860 99482
rect 242808 99418 242860 99424
rect 242820 94518 242848 99418
rect 242808 94512 242860 94518
rect 242808 94454 242860 94460
rect 243556 89593 243584 162114
rect 244384 111790 244412 196590
rect 245212 160818 245240 241604
rect 245658 241496 245714 241505
rect 245658 241431 245714 241440
rect 245568 235340 245620 235346
rect 245568 235282 245620 235288
rect 245200 160812 245252 160818
rect 245200 160754 245252 160760
rect 244924 113824 244976 113830
rect 244924 113766 244976 113772
rect 244372 111784 244424 111790
rect 244372 111726 244424 111732
rect 244384 111110 244412 111726
rect 244372 111104 244424 111110
rect 244372 111046 244424 111052
rect 243542 89584 243598 89593
rect 243542 89519 243598 89528
rect 244280 85536 244332 85542
rect 244280 85478 244332 85484
rect 244292 84862 244320 85478
rect 244280 84856 244332 84862
rect 244280 84798 244332 84804
rect 244280 80096 244332 80102
rect 241610 80064 241666 80073
rect 244280 80038 244332 80044
rect 241610 79999 241666 80008
rect 242992 62824 243044 62830
rect 242992 62766 243044 62772
rect 243004 16574 243032 62766
rect 244292 16574 244320 80038
rect 244936 71738 244964 113766
rect 245580 84862 245608 235282
rect 245672 146169 245700 241431
rect 248418 239728 248474 239737
rect 248418 239663 248474 239672
rect 246304 238128 246356 238134
rect 246304 238070 246356 238076
rect 246316 226273 246344 238070
rect 248432 238066 248460 239663
rect 248524 238814 248552 241604
rect 251284 241590 251850 241618
rect 249064 241528 249116 241534
rect 249064 241470 249116 241476
rect 248512 238808 248564 238814
rect 248512 238750 248564 238756
rect 248420 238060 248472 238066
rect 248420 238002 248472 238008
rect 246394 237960 246450 237969
rect 246394 237895 246450 237904
rect 246302 226264 246358 226273
rect 246302 226199 246358 226208
rect 245658 146160 245714 146169
rect 245658 146095 245714 146104
rect 246304 143608 246356 143614
rect 246304 143550 246356 143556
rect 245568 84856 245620 84862
rect 245568 84798 245620 84804
rect 245660 82136 245712 82142
rect 245660 82078 245712 82084
rect 244924 71732 244976 71738
rect 244924 71674 244976 71680
rect 245672 16574 245700 82078
rect 241532 16546 241744 16574
rect 243004 16546 244136 16574
rect 244292 16546 245240 16574
rect 245672 16546 245976 16574
rect 239312 4888 239364 4894
rect 239312 4830 239364 4836
rect 238024 4820 238076 4826
rect 238024 4762 238076 4768
rect 233884 4072 233936 4078
rect 233884 4014 233936 4020
rect 213184 3460 213236 3466
rect 213184 3402 213236 3408
rect 178684 2100 178736 2106
rect 178684 2042 178736 2048
rect 239324 480 239352 4830
rect 240508 4072 240560 4078
rect 240508 4014 240560 4020
rect 240520 480 240548 4014
rect 241716 480 241744 16546
rect 242900 3460 242952 3466
rect 242900 3402 242952 3408
rect 242912 480 242940 3402
rect 244108 480 244136 16546
rect 245212 480 245240 16546
rect 245948 490 245976 16546
rect 246316 3466 246344 143550
rect 246408 122194 246436 237895
rect 248418 226944 248474 226953
rect 248418 226879 248474 226888
rect 246486 146160 246542 146169
rect 246486 146095 246542 146104
rect 246500 144945 246528 146095
rect 246486 144936 246542 144945
rect 246486 144871 246542 144880
rect 246500 124914 246528 144871
rect 246488 124908 246540 124914
rect 246488 124850 246540 124856
rect 246396 122188 246448 122194
rect 246396 122130 246448 122136
rect 248432 73846 248460 226879
rect 249076 199442 249104 241470
rect 250442 240136 250498 240145
rect 250442 240071 250498 240080
rect 250352 238060 250404 238066
rect 250352 238002 250404 238008
rect 250364 232665 250392 238002
rect 250350 232656 250406 232665
rect 250350 232591 250406 232600
rect 250456 228993 250484 240071
rect 251284 239873 251312 241590
rect 251916 241528 251968 241534
rect 251916 241470 251968 241476
rect 251824 240100 251876 240106
rect 251824 240042 251876 240048
rect 251270 239864 251326 239873
rect 251270 239799 251326 239808
rect 250442 228984 250498 228993
rect 250442 228919 250498 228928
rect 250444 215960 250496 215966
rect 250444 215902 250496 215908
rect 249064 199436 249116 199442
rect 249064 199378 249116 199384
rect 250456 170406 250484 215902
rect 250444 170400 250496 170406
rect 250444 170342 250496 170348
rect 250444 158840 250496 158846
rect 250444 158782 250496 158788
rect 249064 139460 249116 139466
rect 249064 139402 249116 139408
rect 248420 73840 248472 73846
rect 248420 73782 248472 73788
rect 248420 50380 248472 50386
rect 248420 50322 248472 50328
rect 247040 24132 247092 24138
rect 247040 24074 247092 24080
rect 247052 16574 247080 24074
rect 247052 16546 247632 16574
rect 246304 3460 246356 3466
rect 246304 3402 246356 3408
rect 246224 598 246436 626
rect 246224 490 246252 598
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 245948 462 246252 490
rect 246408 480 246436 598
rect 247604 480 247632 16546
rect 248432 490 248460 50322
rect 249076 3534 249104 139402
rect 250456 40730 250484 158782
rect 251180 150544 251232 150550
rect 251180 150486 251232 150492
rect 250536 98048 250588 98054
rect 250536 97990 250588 97996
rect 250548 68950 250576 97990
rect 250536 68944 250588 68950
rect 250536 68886 250588 68892
rect 249800 40724 249852 40730
rect 249800 40666 249852 40672
rect 250444 40724 250496 40730
rect 250444 40666 250496 40672
rect 249812 16574 249840 40666
rect 250548 24138 250576 68886
rect 250536 24132 250588 24138
rect 250536 24074 250588 24080
rect 249812 16546 250024 16574
rect 249064 3528 249116 3534
rect 249064 3470 249116 3476
rect 248616 598 248828 626
rect 248616 490 248644 598
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248432 462 248644 490
rect 248800 480 248828 598
rect 249996 480 250024 16546
rect 251192 11830 251220 150486
rect 251284 91905 251312 239799
rect 251836 216034 251864 240042
rect 251928 230489 251956 241470
rect 252468 235272 252520 235278
rect 252468 235214 252520 235220
rect 251914 230480 251970 230489
rect 251914 230415 251970 230424
rect 251824 216028 251876 216034
rect 251824 215970 251876 215976
rect 252480 156738 252508 235214
rect 252664 229945 252692 296398
rect 252940 292574 252968 304982
rect 253204 304360 253256 304366
rect 253204 304302 253256 304308
rect 253020 302252 253072 302258
rect 253020 302194 253072 302200
rect 253032 296585 253060 302194
rect 253216 301580 253244 304302
rect 253308 301578 253336 335310
rect 254596 318073 254624 356662
rect 254768 327752 254820 327758
rect 254768 327694 254820 327700
rect 254582 318064 254638 318073
rect 254582 317999 254638 318008
rect 254582 314120 254638 314129
rect 254582 314055 254638 314064
rect 253938 313984 253994 313993
rect 253938 313919 253994 313928
rect 253664 302184 253716 302190
rect 253664 302126 253716 302132
rect 253296 301572 253348 301578
rect 253296 301514 253348 301520
rect 253112 301368 253164 301374
rect 253676 301345 253704 302126
rect 253112 301310 253164 301316
rect 253662 301336 253718 301345
rect 253124 299033 253152 301310
rect 253662 301271 253718 301280
rect 253110 299024 253166 299033
rect 253110 298959 253166 298968
rect 253124 298246 253152 298959
rect 253112 298240 253164 298246
rect 253112 298182 253164 298188
rect 253202 296984 253258 296993
rect 253202 296919 253258 296928
rect 253018 296576 253074 296585
rect 253018 296511 253074 296520
rect 252940 292546 253152 292574
rect 253124 289814 253152 292546
rect 253216 289921 253244 296919
rect 253202 289912 253258 289921
rect 253202 289847 253258 289856
rect 252848 289786 253152 289814
rect 252848 285433 252876 289786
rect 253846 289640 253902 289649
rect 253846 289575 253902 289584
rect 253664 288788 253716 288794
rect 253664 288730 253716 288736
rect 252834 285424 252890 285433
rect 252834 285359 252890 285368
rect 253676 283937 253704 288730
rect 253860 288454 253888 289575
rect 253848 288448 253900 288454
rect 253848 288390 253900 288396
rect 253662 283928 253718 283937
rect 253662 283863 253718 283872
rect 252926 266384 252982 266393
rect 252926 266319 252982 266328
rect 252834 253192 252890 253201
rect 252834 253127 252890 253136
rect 252848 248414 252876 253127
rect 252756 248386 252876 248414
rect 252756 240009 252784 248386
rect 252940 247110 252968 266319
rect 253952 253745 253980 313919
rect 254214 308544 254270 308553
rect 254214 308479 254270 308488
rect 254124 301572 254176 301578
rect 254124 301514 254176 301520
rect 254136 288794 254164 301514
rect 254124 288788 254176 288794
rect 254124 288730 254176 288736
rect 254122 263256 254178 263265
rect 254122 263191 254178 263200
rect 253938 253736 253994 253745
rect 253938 253671 253994 253680
rect 253938 249520 253994 249529
rect 253938 249455 253994 249464
rect 252928 247104 252980 247110
rect 252928 247046 252980 247052
rect 253204 243568 253256 243574
rect 253204 243510 253256 243516
rect 252834 242856 252890 242865
rect 252834 242791 252890 242800
rect 252742 240000 252798 240009
rect 252742 239935 252798 239944
rect 252848 238754 252876 242791
rect 252926 242448 252982 242457
rect 252926 242383 252982 242392
rect 252940 241534 252968 242383
rect 252928 241528 252980 241534
rect 252928 241470 252980 241476
rect 252756 238726 252876 238754
rect 252650 229936 252706 229945
rect 252650 229871 252706 229880
rect 252756 182889 252784 238726
rect 253216 235346 253244 243510
rect 253204 235340 253256 235346
rect 253204 235282 253256 235288
rect 253204 229764 253256 229770
rect 253204 229706 253256 229712
rect 252742 182880 252798 182889
rect 252742 182815 252798 182824
rect 252468 156732 252520 156738
rect 252468 156674 252520 156680
rect 253216 97986 253244 229706
rect 253952 209098 253980 249455
rect 254032 247104 254084 247110
rect 254032 247046 254084 247052
rect 254044 240106 254072 247046
rect 254032 240100 254084 240106
rect 254032 240042 254084 240048
rect 254136 221474 254164 263191
rect 254228 247489 254256 308479
rect 254596 259593 254624 314055
rect 254780 313993 254808 327694
rect 255332 325694 255360 444751
rect 255424 443465 255452 474710
rect 255596 472048 255648 472054
rect 255596 471990 255648 471996
rect 255608 460934 255636 471990
rect 262220 470620 262272 470626
rect 262220 470562 262272 470568
rect 258078 467936 258134 467945
rect 258078 467871 258134 467880
rect 256700 465180 256752 465186
rect 256700 465122 256752 465128
rect 255608 460906 256096 460934
rect 255962 454064 256018 454073
rect 255962 453999 256018 454008
rect 255976 448905 256004 453999
rect 255962 448896 256018 448905
rect 255962 448831 256018 448840
rect 255686 446176 255742 446185
rect 255686 446111 255742 446120
rect 255700 443698 255728 446111
rect 255688 443692 255740 443698
rect 255688 443634 255740 443640
rect 255410 443456 255466 443465
rect 255410 443391 255466 443400
rect 255424 443018 255452 443391
rect 255412 443012 255464 443018
rect 255412 442954 255464 442960
rect 255412 439544 255464 439550
rect 255412 439486 255464 439492
rect 255424 439113 255452 439486
rect 255410 439104 255466 439113
rect 255410 439039 255466 439048
rect 255504 438864 255556 438870
rect 255504 438806 255556 438812
rect 255516 437753 255544 438806
rect 255502 437744 255558 437753
rect 255502 437679 255558 437688
rect 255504 437436 255556 437442
rect 255504 437378 255556 437384
rect 255516 436801 255544 437378
rect 255502 436792 255558 436801
rect 255502 436727 255558 436736
rect 255412 435396 255464 435402
rect 255412 435338 255464 435344
rect 255424 435033 255452 435338
rect 255410 435024 255466 435033
rect 255410 434959 255466 434968
rect 255412 434648 255464 434654
rect 255412 434590 255464 434596
rect 255424 433673 255452 434590
rect 255410 433664 255466 433673
rect 255410 433599 255466 433608
rect 255976 432682 256004 448831
rect 256068 446185 256096 460906
rect 256054 446176 256110 446185
rect 256054 446111 256110 446120
rect 255964 432676 256016 432682
rect 255964 432618 256016 432624
rect 255594 430672 255650 430681
rect 255594 430607 255650 430616
rect 255410 427952 255466 427961
rect 255410 427887 255466 427896
rect 255424 427854 255452 427887
rect 255412 427848 255464 427854
rect 255412 427790 255464 427796
rect 255504 427780 255556 427786
rect 255504 427722 255556 427728
rect 255516 426601 255544 427722
rect 255502 426592 255558 426601
rect 255502 426527 255558 426536
rect 255608 426442 255636 430607
rect 256606 429312 256662 429321
rect 256712 429298 256740 465122
rect 256792 458244 256844 458250
rect 256792 458186 256844 458192
rect 256662 429270 256740 429298
rect 256606 429247 256662 429256
rect 255424 426414 255636 426442
rect 255424 387734 255452 426414
rect 256606 425232 256662 425241
rect 256804 425218 256832 458186
rect 258092 434654 258120 467871
rect 259552 463820 259604 463826
rect 259552 463762 259604 463768
rect 258264 459604 258316 459610
rect 258264 459546 258316 459552
rect 258170 452704 258226 452713
rect 258170 452639 258226 452648
rect 258080 434648 258132 434654
rect 258080 434590 258132 434596
rect 256662 425190 256832 425218
rect 256606 425167 256662 425176
rect 256804 424386 256832 425190
rect 256792 424380 256844 424386
rect 256792 424322 256844 424328
rect 255502 423600 255558 423609
rect 255502 423535 255558 423544
rect 255516 422346 255544 423535
rect 255504 422340 255556 422346
rect 255504 422282 255556 422288
rect 255502 422240 255558 422249
rect 255502 422175 255558 422184
rect 255516 420986 255544 422175
rect 255504 420980 255556 420986
rect 255504 420922 255556 420928
rect 255594 420880 255650 420889
rect 255594 420815 255650 420824
rect 255608 419558 255636 420815
rect 255596 419552 255648 419558
rect 255502 419520 255558 419529
rect 255596 419494 255648 419500
rect 255502 419455 255558 419464
rect 255516 418198 255544 419455
rect 255504 418192 255556 418198
rect 255504 418134 255556 418140
rect 255594 418160 255650 418169
rect 255594 418095 255650 418104
rect 255608 416906 255636 418095
rect 255596 416900 255648 416906
rect 255596 416842 255648 416848
rect 255504 416832 255556 416838
rect 255502 416800 255504 416809
rect 255556 416800 255558 416809
rect 255502 416735 255558 416744
rect 256606 415168 256662 415177
rect 256662 415126 256740 415154
rect 256606 415103 256662 415112
rect 255502 412448 255558 412457
rect 255502 412383 255558 412392
rect 255516 411602 255544 412383
rect 255504 411596 255556 411602
rect 255504 411538 255556 411544
rect 255502 411088 255558 411097
rect 255502 411023 255558 411032
rect 255516 409970 255544 411023
rect 255504 409964 255556 409970
rect 255504 409906 255556 409912
rect 255502 409728 255558 409737
rect 255502 409663 255558 409672
rect 255516 408542 255544 409663
rect 255504 408536 255556 408542
rect 255504 408478 255556 408484
rect 255502 408368 255558 408377
rect 255502 408303 255558 408312
rect 255516 407250 255544 408303
rect 255504 407244 255556 407250
rect 255504 407186 255556 407192
rect 255502 407008 255558 407017
rect 255502 406943 255558 406952
rect 255516 405754 255544 406943
rect 255504 405748 255556 405754
rect 255504 405690 255556 405696
rect 255502 404016 255558 404025
rect 255502 403951 255558 403960
rect 255516 403442 255544 403951
rect 255504 403436 255556 403442
rect 255504 403378 255556 403384
rect 255502 401296 255558 401305
rect 255502 401231 255558 401240
rect 255516 400246 255544 401231
rect 255504 400240 255556 400246
rect 255504 400182 255556 400188
rect 255502 399936 255558 399945
rect 255502 399871 255558 399880
rect 255516 398886 255544 399871
rect 255504 398880 255556 398886
rect 255504 398822 255556 398828
rect 255502 398576 255558 398585
rect 255502 398511 255558 398520
rect 255516 397526 255544 398511
rect 255504 397520 255556 397526
rect 255504 397462 255556 397468
rect 255502 396944 255558 396953
rect 255502 396879 255558 396888
rect 255412 387728 255464 387734
rect 255412 387670 255464 387676
rect 255424 329118 255452 387670
rect 255516 375290 255544 396879
rect 255594 394224 255650 394233
rect 255594 394159 255650 394168
rect 255608 393378 255636 394159
rect 255596 393372 255648 393378
rect 255596 393314 255648 393320
rect 256712 378146 256740 415126
rect 258080 411596 258132 411602
rect 258080 411538 258132 411544
rect 257344 403436 257396 403442
rect 257344 403378 257396 403384
rect 256700 378140 256752 378146
rect 256700 378082 256752 378088
rect 256698 377360 256754 377369
rect 256698 377295 256754 377304
rect 256712 376786 256740 377295
rect 257356 376786 257384 403378
rect 258092 390998 258120 411538
rect 258080 390992 258132 390998
rect 258080 390934 258132 390940
rect 258078 386472 258134 386481
rect 258078 386407 258134 386416
rect 256700 376780 256752 376786
rect 256700 376722 256752 376728
rect 257344 376780 257396 376786
rect 257344 376722 257396 376728
rect 255504 375284 255556 375290
rect 255504 375226 255556 375232
rect 255412 329112 255464 329118
rect 255412 329054 255464 329060
rect 255516 328409 255544 375226
rect 255502 328400 255558 328409
rect 255502 328335 255558 328344
rect 256700 327208 256752 327214
rect 256700 327150 256752 327156
rect 255332 325666 255728 325694
rect 255700 323610 255728 325666
rect 255688 323604 255740 323610
rect 255688 323546 255740 323552
rect 254766 313984 254822 313993
rect 254766 313919 254822 313928
rect 255412 310616 255464 310622
rect 255412 310558 255464 310564
rect 255424 292641 255452 310558
rect 255504 309800 255556 309806
rect 255504 309742 255556 309748
rect 255516 293865 255544 309742
rect 255596 308440 255648 308446
rect 255596 308382 255648 308388
rect 255608 295089 255636 308382
rect 255594 295080 255650 295089
rect 255594 295015 255650 295024
rect 255502 293856 255558 293865
rect 255502 293791 255558 293800
rect 255410 292632 255466 292641
rect 255410 292567 255466 292576
rect 255412 292256 255464 292262
rect 255410 292224 255412 292233
rect 255464 292224 255466 292233
rect 255410 292159 255466 292168
rect 255410 290864 255466 290873
rect 255410 290799 255466 290808
rect 255424 290562 255452 290799
rect 255412 290556 255464 290562
rect 255412 290498 255464 290504
rect 255516 290442 255544 293791
rect 255700 293457 255728 323546
rect 256606 300792 256662 300801
rect 256606 300727 256662 300736
rect 256514 300384 256570 300393
rect 256514 300319 256570 300328
rect 256528 299538 256556 300319
rect 256620 299606 256648 300727
rect 256608 299600 256660 299606
rect 256608 299542 256660 299548
rect 256516 299532 256568 299538
rect 256516 299474 256568 299480
rect 256606 298344 256662 298353
rect 256606 298279 256662 298288
rect 256620 298178 256648 298279
rect 256608 298172 256660 298178
rect 256608 298114 256660 298120
rect 256606 297936 256662 297945
rect 256606 297871 256662 297880
rect 256514 297528 256570 297537
rect 255872 297492 255924 297498
rect 256514 297463 256570 297472
rect 255872 297434 255924 297440
rect 255884 297129 255912 297434
rect 256528 297430 256556 297463
rect 256516 297424 256568 297430
rect 256516 297366 256568 297372
rect 255870 297120 255926 297129
rect 255870 297055 255926 297064
rect 256620 296993 256648 297871
rect 256606 296984 256662 296993
rect 256606 296919 256662 296928
rect 256608 295996 256660 296002
rect 256608 295938 256660 295944
rect 256620 295497 256648 295938
rect 256606 295488 256662 295497
rect 256606 295423 256662 295432
rect 256606 295080 256662 295089
rect 256606 295015 256608 295024
rect 256660 295015 256662 295024
rect 256608 294986 256660 294992
rect 256606 294264 256662 294273
rect 256606 294199 256662 294208
rect 256620 294030 256648 294199
rect 256608 294024 256660 294030
rect 256608 293966 256660 293972
rect 255686 293448 255742 293457
rect 255686 293383 255742 293392
rect 256606 293040 256662 293049
rect 256606 292975 256662 292984
rect 256620 292942 256648 292975
rect 256608 292936 256660 292942
rect 256608 292878 256660 292884
rect 255424 290414 255544 290442
rect 255320 288380 255372 288386
rect 255320 288322 255372 288328
rect 255332 287609 255360 288322
rect 255318 287600 255374 287609
rect 255318 287535 255374 287544
rect 255424 287054 255452 290414
rect 255504 289808 255556 289814
rect 255504 289750 255556 289756
rect 255516 288833 255544 289750
rect 255502 288824 255558 288833
rect 255502 288759 255558 288768
rect 255504 288312 255556 288318
rect 255504 288254 255556 288260
rect 255516 287201 255544 288254
rect 255502 287192 255558 287201
rect 255502 287127 255558 287136
rect 255332 287026 255452 287054
rect 255044 263288 255096 263294
rect 255042 263256 255044 263265
rect 255096 263256 255098 263265
rect 255042 263191 255098 263200
rect 254582 259584 254638 259593
rect 254582 259519 254638 259528
rect 254596 258505 254624 259519
rect 254582 258496 254638 258505
rect 254582 258431 254638 258440
rect 255226 254824 255282 254833
rect 255226 254759 255282 254768
rect 255240 254425 255268 254759
rect 255226 254416 255282 254425
rect 255226 254351 255282 254360
rect 254952 249756 255004 249762
rect 254952 249698 255004 249704
rect 254964 249529 254992 249698
rect 254950 249520 255006 249529
rect 254950 249455 255006 249464
rect 254582 248704 254638 248713
rect 254582 248639 254638 248648
rect 254214 247480 254270 247489
rect 254214 247415 254270 247424
rect 254228 247110 254256 247415
rect 254216 247104 254268 247110
rect 254216 247046 254268 247052
rect 254596 232558 254624 248639
rect 255332 233918 255360 287026
rect 255504 287020 255556 287026
rect 255504 286962 255556 286968
rect 255412 286952 255464 286958
rect 255412 286894 255464 286900
rect 255424 285977 255452 286894
rect 255516 286385 255544 286962
rect 255502 286376 255558 286385
rect 255502 286311 255558 286320
rect 255410 285968 255466 285977
rect 255410 285903 255466 285912
rect 255410 285560 255466 285569
rect 255410 285495 255466 285504
rect 255424 284345 255452 285495
rect 255410 284336 255466 284345
rect 255410 284271 255466 284280
rect 255504 284300 255556 284306
rect 255504 284242 255556 284248
rect 255516 283121 255544 284242
rect 255502 283112 255558 283121
rect 255502 283047 255558 283056
rect 255504 282872 255556 282878
rect 255504 282814 255556 282820
rect 255516 282713 255544 282814
rect 255502 282704 255558 282713
rect 255502 282639 255558 282648
rect 255412 281920 255464 281926
rect 255410 281888 255412 281897
rect 255464 281888 255466 281897
rect 255410 281823 255466 281832
rect 255412 281376 255464 281382
rect 255410 281344 255412 281353
rect 255464 281344 255466 281353
rect 255410 281279 255466 281288
rect 255412 281240 255464 281246
rect 255412 281182 255464 281188
rect 255424 280537 255452 281182
rect 255410 280528 255466 280537
rect 255410 280463 255466 280472
rect 255412 280152 255464 280158
rect 255410 280120 255412 280129
rect 255464 280120 255466 280129
rect 255410 280055 255466 280064
rect 255504 280084 255556 280090
rect 255504 280026 255556 280032
rect 255516 278905 255544 280026
rect 256712 279313 256740 327150
rect 256790 325816 256846 325825
rect 256790 325751 256846 325760
rect 256804 290057 256832 325751
rect 256884 315308 256936 315314
rect 256884 315250 256936 315256
rect 256790 290048 256846 290057
rect 256790 289983 256846 289992
rect 256896 284753 256924 315250
rect 256976 314084 257028 314090
rect 256976 314026 257028 314032
rect 256988 298761 257016 314026
rect 256974 298752 257030 298761
rect 256974 298687 257030 298696
rect 258092 294642 258120 386407
rect 258184 351218 258212 452639
rect 258276 439550 258304 459546
rect 259460 452736 259512 452742
rect 259460 452678 259512 452684
rect 258816 443012 258868 443018
rect 258816 442954 258868 442960
rect 258264 439544 258316 439550
rect 258264 439486 258316 439492
rect 258828 429894 258856 442954
rect 258724 429888 258776 429894
rect 258724 429830 258776 429836
rect 258816 429888 258868 429894
rect 258816 429830 258868 429836
rect 258264 409964 258316 409970
rect 258264 409906 258316 409912
rect 258276 375329 258304 409906
rect 258736 403617 258764 429830
rect 258722 403608 258778 403617
rect 258722 403543 258778 403552
rect 258356 398880 258408 398886
rect 258356 398822 258408 398828
rect 258368 382265 258396 398822
rect 258354 382256 258410 382265
rect 258354 382191 258410 382200
rect 258262 375320 258318 375329
rect 258262 375255 258318 375264
rect 258172 351212 258224 351218
rect 258172 351154 258224 351160
rect 258172 341624 258224 341630
rect 258172 341566 258224 341572
rect 258184 295882 258212 341566
rect 258264 329112 258316 329118
rect 258264 329054 258316 329060
rect 258276 296002 258304 329054
rect 259472 316742 259500 452678
rect 259564 435402 259592 463762
rect 260930 461000 260986 461009
rect 260930 460935 260986 460944
rect 260840 456884 260892 456890
rect 260840 456826 260892 456832
rect 260104 455524 260156 455530
rect 260104 455466 260156 455472
rect 259552 435396 259604 435402
rect 259552 435338 259604 435344
rect 259552 407244 259604 407250
rect 259552 407186 259604 407192
rect 259564 384334 259592 407186
rect 259552 384328 259604 384334
rect 259552 384270 259604 384276
rect 259552 362976 259604 362982
rect 259552 362918 259604 362924
rect 259460 316736 259512 316742
rect 259460 316678 259512 316684
rect 259472 316577 259500 316678
rect 259458 316568 259514 316577
rect 259458 316503 259514 316512
rect 258356 308508 258408 308514
rect 258356 308450 258408 308456
rect 258368 306374 258396 308450
rect 258368 306346 258488 306374
rect 258264 295996 258316 296002
rect 258264 295938 258316 295944
rect 258184 295854 258304 295882
rect 258276 294794 258304 295854
rect 258184 294766 258304 294794
rect 258080 294636 258132 294642
rect 258080 294578 258132 294584
rect 257066 291816 257122 291825
rect 257066 291751 257122 291760
rect 256882 284744 256938 284753
rect 256882 284679 256938 284688
rect 256698 279304 256754 279313
rect 256698 279239 256754 279248
rect 255502 278896 255558 278905
rect 255502 278831 255558 278840
rect 255412 278724 255464 278730
rect 255412 278666 255464 278672
rect 255424 277681 255452 278666
rect 255410 277672 255466 277681
rect 255410 277607 255466 277616
rect 255412 277364 255464 277370
rect 255412 277306 255464 277312
rect 255424 276457 255452 277306
rect 255504 277296 255556 277302
rect 255504 277238 255556 277244
rect 255410 276448 255466 276457
rect 255410 276383 255466 276392
rect 255516 276049 255544 277238
rect 255502 276040 255558 276049
rect 255412 276004 255464 276010
rect 255502 275975 255558 275984
rect 255412 275946 255464 275952
rect 255424 275233 255452 275946
rect 255410 275224 255466 275233
rect 255410 275159 255466 275168
rect 255410 274816 255466 274825
rect 255410 274751 255466 274760
rect 255424 274718 255452 274751
rect 255412 274712 255464 274718
rect 255412 274654 255464 274660
rect 255504 274644 255556 274650
rect 255504 274586 255556 274592
rect 255412 274576 255464 274582
rect 255412 274518 255464 274524
rect 255424 274417 255452 274518
rect 255410 274408 255466 274417
rect 255410 274343 255466 274352
rect 255516 274009 255544 274586
rect 255502 274000 255558 274009
rect 255502 273935 255558 273944
rect 255504 273216 255556 273222
rect 255410 273184 255466 273193
rect 255504 273158 255556 273164
rect 255410 273119 255412 273128
rect 255464 273119 255466 273128
rect 255412 273090 255464 273096
rect 255516 272785 255544 273158
rect 255502 272776 255558 272785
rect 255502 272711 255558 272720
rect 256882 271960 256938 271969
rect 256882 271895 256938 271904
rect 255412 271856 255464 271862
rect 255412 271798 255464 271804
rect 255424 271425 255452 271798
rect 255410 271416 255466 271425
rect 255410 271351 255466 271360
rect 255410 270600 255466 270609
rect 255410 270535 255412 270544
rect 255464 270535 255466 270544
rect 255412 270506 255464 270512
rect 255504 270496 255556 270502
rect 255504 270438 255556 270444
rect 255516 270201 255544 270438
rect 255502 270192 255558 270201
rect 255502 270127 255558 270136
rect 255410 269784 255466 269793
rect 255410 269719 255466 269728
rect 255424 269142 255452 269719
rect 256698 269376 256754 269385
rect 256698 269311 256754 269320
rect 255412 269136 255464 269142
rect 255412 269078 255464 269084
rect 255412 269000 255464 269006
rect 255410 268968 255412 268977
rect 255464 268968 255466 268977
rect 255410 268903 255466 268912
rect 255504 268932 255556 268938
rect 255504 268874 255556 268880
rect 255516 268161 255544 268874
rect 255502 268152 255558 268161
rect 255502 268087 255558 268096
rect 255502 267744 255558 267753
rect 255502 267679 255558 267688
rect 255412 267028 255464 267034
rect 255412 266970 255464 266976
rect 255424 266937 255452 266970
rect 255410 266928 255466 266937
rect 255410 266863 255466 266872
rect 255516 266422 255544 267679
rect 255504 266416 255556 266422
rect 255504 266358 255556 266364
rect 255412 266348 255464 266354
rect 255412 266290 255464 266296
rect 255424 265305 255452 266290
rect 255502 266112 255558 266121
rect 255502 266047 255558 266056
rect 255410 265296 255466 265305
rect 255410 265231 255466 265240
rect 255516 264994 255544 266047
rect 255504 264988 255556 264994
rect 255504 264930 255556 264936
rect 255594 264888 255650 264897
rect 255594 264823 255650 264832
rect 255410 264480 255466 264489
rect 255410 264415 255466 264424
rect 255424 264246 255452 264415
rect 255412 264240 255464 264246
rect 255412 264182 255464 264188
rect 255410 264072 255466 264081
rect 255410 264007 255466 264016
rect 255424 263634 255452 264007
rect 255502 263800 255558 263809
rect 255502 263735 255558 263744
rect 255412 263628 255464 263634
rect 255412 263570 255464 263576
rect 255516 262449 255544 263735
rect 255608 262886 255636 264823
rect 255596 262880 255648 262886
rect 255596 262822 255648 262828
rect 255502 262440 255558 262449
rect 255502 262375 255558 262384
rect 255412 260840 255464 260846
rect 255412 260782 255464 260788
rect 255424 260681 255452 260782
rect 255410 260672 255466 260681
rect 255410 260607 255466 260616
rect 255594 260264 255650 260273
rect 255594 260199 255650 260208
rect 255504 259480 255556 259486
rect 255410 259448 255466 259457
rect 255504 259422 255556 259428
rect 255410 259383 255412 259392
rect 255464 259383 255466 259392
rect 255412 259354 255464 259360
rect 255516 258641 255544 259422
rect 255608 258777 255636 260199
rect 255594 258768 255650 258777
rect 255594 258703 255650 258712
rect 255502 258632 255558 258641
rect 255502 258567 255558 258576
rect 255412 257440 255464 257446
rect 255410 257408 255412 257417
rect 255464 257408 255466 257417
rect 255410 257343 255466 257352
rect 255410 257000 255466 257009
rect 255410 256935 255466 256944
rect 255424 256766 255452 256935
rect 255412 256760 255464 256766
rect 255412 256702 255464 256708
rect 255410 256592 255466 256601
rect 255410 256527 255466 256536
rect 255424 256018 255452 256527
rect 255594 256184 255650 256193
rect 255594 256119 255650 256128
rect 255504 256080 255556 256086
rect 255504 256022 255556 256028
rect 255412 256012 255464 256018
rect 255412 255954 255464 255960
rect 255516 255377 255544 256022
rect 255502 255368 255558 255377
rect 255502 255303 255558 255312
rect 255504 255264 255556 255270
rect 255504 255206 255556 255212
rect 255410 254552 255466 254561
rect 255410 254487 255466 254496
rect 255424 253978 255452 254487
rect 255516 254153 255544 255206
rect 255608 254561 255636 256119
rect 255594 254552 255650 254561
rect 255594 254487 255650 254496
rect 255502 254144 255558 254153
rect 255502 254079 255558 254088
rect 255412 253972 255464 253978
rect 255412 253914 255464 253920
rect 255412 253292 255464 253298
rect 255412 253234 255464 253240
rect 255424 252929 255452 253234
rect 255410 252920 255466 252929
rect 255410 252855 255466 252864
rect 255410 252512 255466 252521
rect 255410 252447 255466 252456
rect 255424 251870 255452 252447
rect 255502 252104 255558 252113
rect 255502 252039 255558 252048
rect 255412 251864 255464 251870
rect 255412 251806 255464 251812
rect 255516 251258 255544 252039
rect 255504 251252 255556 251258
rect 255504 251194 255556 251200
rect 255502 251152 255558 251161
rect 255502 251087 255558 251096
rect 255516 249830 255544 251087
rect 255872 249960 255924 249966
rect 255870 249928 255872 249937
rect 255924 249928 255926 249937
rect 255870 249863 255926 249872
rect 255504 249824 255556 249830
rect 255504 249766 255556 249772
rect 255410 249112 255466 249121
rect 255410 249047 255412 249056
rect 255464 249047 255466 249056
rect 255412 249018 255464 249024
rect 255504 247716 255556 247722
rect 255504 247658 255556 247664
rect 255516 247081 255544 247658
rect 255502 247072 255558 247081
rect 255502 247007 255558 247016
rect 255410 246664 255466 246673
rect 255410 246599 255466 246608
rect 255424 246362 255452 246599
rect 255412 246356 255464 246362
rect 255412 246298 255464 246304
rect 255686 246256 255742 246265
rect 255686 246191 255742 246200
rect 255410 245848 255466 245857
rect 255410 245783 255412 245792
rect 255464 245783 255466 245792
rect 255412 245754 255464 245760
rect 255412 245608 255464 245614
rect 255412 245550 255464 245556
rect 255424 245449 255452 245550
rect 255410 245440 255466 245449
rect 255410 245375 255466 245384
rect 255594 245032 255650 245041
rect 255594 244967 255650 244976
rect 255502 244624 255558 244633
rect 255502 244559 255558 244568
rect 255516 244322 255544 244559
rect 255504 244316 255556 244322
rect 255504 244258 255556 244264
rect 255412 244248 255464 244254
rect 255410 244216 255412 244225
rect 255464 244216 255466 244225
rect 255410 244151 255466 244160
rect 255502 243808 255558 243817
rect 255502 243743 255558 243752
rect 255410 240952 255466 240961
rect 255410 240887 255466 240896
rect 255424 240854 255452 240887
rect 255412 240848 255464 240854
rect 255412 240790 255464 240796
rect 255516 238754 255544 243743
rect 255608 242321 255636 244967
rect 255594 242312 255650 242321
rect 255594 242247 255650 242256
rect 255594 240816 255650 240825
rect 255700 240802 255728 246191
rect 256054 242176 256110 242185
rect 256054 242111 256110 242120
rect 255650 240774 255728 240802
rect 255594 240751 255596 240760
rect 255648 240751 255650 240760
rect 255596 240722 255648 240728
rect 256068 239290 256096 242111
rect 256056 239284 256108 239290
rect 256056 239226 256108 239232
rect 255424 238726 255544 238754
rect 255424 236609 255452 238726
rect 255410 236600 255466 236609
rect 255410 236535 255466 236544
rect 255320 233912 255372 233918
rect 255320 233854 255372 233860
rect 254584 232552 254636 232558
rect 254584 232494 254636 232500
rect 254124 221468 254176 221474
rect 254124 221410 254176 221416
rect 254596 218754 254624 232494
rect 254584 218748 254636 218754
rect 254584 218690 254636 218696
rect 255962 214568 256018 214577
rect 255962 214503 256018 214512
rect 254584 211812 254636 211818
rect 254584 211754 254636 211760
rect 253940 209092 253992 209098
rect 253940 209034 253992 209040
rect 253294 140040 253350 140049
rect 253294 139975 253350 139984
rect 253204 97980 253256 97986
rect 253204 97922 253256 97928
rect 251270 91896 251326 91905
rect 251270 91831 251326 91840
rect 251284 91225 251312 91831
rect 251270 91216 251326 91225
rect 251270 91151 251326 91160
rect 251822 91216 251878 91225
rect 251822 91151 251878 91160
rect 251836 43450 251864 91151
rect 253204 44872 253256 44878
rect 253204 44814 253256 44820
rect 251824 43444 251876 43450
rect 251824 43386 251876 43392
rect 251180 11824 251232 11830
rect 251180 11766 251232 11772
rect 252376 11824 252428 11830
rect 252376 11766 252428 11772
rect 251180 6248 251232 6254
rect 251180 6190 251232 6196
rect 251192 480 251220 6190
rect 252388 480 252416 11766
rect 253216 3398 253244 44814
rect 253308 18630 253336 139975
rect 254596 113830 254624 211754
rect 255976 205057 256004 214503
rect 256054 207632 256110 207641
rect 256054 207567 256110 207576
rect 255318 205048 255374 205057
rect 255318 204983 255374 204992
rect 255962 205048 256018 205057
rect 255962 204983 256018 204992
rect 254584 113824 254636 113830
rect 254584 113766 254636 113772
rect 255332 90953 255360 204983
rect 255964 156732 256016 156738
rect 255964 156674 256016 156680
rect 255318 90944 255374 90953
rect 255318 90879 255374 90888
rect 253296 18624 253348 18630
rect 253296 18566 253348 18572
rect 255976 9042 256004 156674
rect 256068 153105 256096 207567
rect 256712 207058 256740 269311
rect 256896 240038 256924 271895
rect 257080 241602 257108 291751
rect 258184 283529 258212 294766
rect 258264 294636 258316 294642
rect 258264 294578 258316 294584
rect 258170 283520 258226 283529
rect 258170 283455 258226 283464
rect 258276 280809 258304 294578
rect 258460 290562 258488 306346
rect 259460 305652 259512 305658
rect 259460 305594 259512 305600
rect 259368 296676 259420 296682
rect 259368 296618 259420 296624
rect 259380 292262 259408 296618
rect 259368 292256 259420 292262
rect 259368 292198 259420 292204
rect 258448 290556 258500 290562
rect 258448 290498 258500 290504
rect 258724 290488 258776 290494
rect 258724 290430 258776 290436
rect 258262 280800 258318 280809
rect 258262 280735 258318 280744
rect 258736 279721 258764 290430
rect 259092 284232 259144 284238
rect 259092 284174 259144 284180
rect 259104 281382 259132 284174
rect 259472 281926 259500 305594
rect 259564 297430 259592 362918
rect 259644 329928 259696 329934
rect 259644 329870 259696 329876
rect 259552 297424 259604 297430
rect 259552 297366 259604 297372
rect 259656 292942 259684 329870
rect 260116 305833 260144 455466
rect 260852 334626 260880 456826
rect 260944 427786 260972 460935
rect 262232 438870 262260 470562
rect 269120 452668 269172 452674
rect 269120 452610 269172 452616
rect 263598 450256 263654 450265
rect 263598 450191 263654 450200
rect 262864 449948 262916 449954
rect 262864 449890 262916 449896
rect 262220 438864 262272 438870
rect 262220 438806 262272 438812
rect 262232 437510 262260 438806
rect 262220 437504 262272 437510
rect 262220 437446 262272 437452
rect 262220 432676 262272 432682
rect 262220 432618 262272 432624
rect 260932 427780 260984 427786
rect 260932 427722 260984 427728
rect 262128 427780 262180 427786
rect 262128 427722 262180 427728
rect 262140 427106 262168 427722
rect 262128 427100 262180 427106
rect 262128 427042 262180 427048
rect 262128 417444 262180 417450
rect 262128 417386 262180 417392
rect 262140 416906 262168 417386
rect 260932 416900 260984 416906
rect 260932 416842 260984 416848
rect 262128 416900 262180 416906
rect 262128 416842 262180 416848
rect 260944 376553 260972 416842
rect 260930 376544 260986 376553
rect 260930 376479 260986 376488
rect 261482 376544 261538 376553
rect 261482 376479 261538 376488
rect 261496 363089 261524 376479
rect 262232 373318 262260 432618
rect 262220 373312 262272 373318
rect 262220 373254 262272 373260
rect 261482 363080 261538 363089
rect 261482 363015 261538 363024
rect 260932 359508 260984 359514
rect 260932 359450 260984 359456
rect 260840 334620 260892 334626
rect 260840 334562 260892 334568
rect 260102 305824 260158 305833
rect 260102 305759 260158 305768
rect 259734 302832 259790 302841
rect 259734 302767 259790 302776
rect 259644 292936 259696 292942
rect 259644 292878 259696 292884
rect 259460 281920 259512 281926
rect 259460 281862 259512 281868
rect 259092 281376 259144 281382
rect 259092 281318 259144 281324
rect 259748 281246 259776 302767
rect 260840 302320 260892 302326
rect 260840 302262 260892 302268
rect 260748 292936 260800 292942
rect 260748 292878 260800 292884
rect 260760 291854 260788 292878
rect 260748 291848 260800 291854
rect 260748 291790 260800 291796
rect 259736 281240 259788 281246
rect 259736 281182 259788 281188
rect 258814 280936 258870 280945
rect 258814 280871 258870 280880
rect 258722 279712 258778 279721
rect 258722 279647 258778 279656
rect 258078 276856 258134 276865
rect 258078 276791 258134 276800
rect 257342 269784 257398 269793
rect 257342 269719 257398 269728
rect 257356 249966 257384 269719
rect 257344 249960 257396 249966
rect 257344 249902 257396 249908
rect 257356 248414 257384 249902
rect 257264 248386 257384 248414
rect 257068 241596 257120 241602
rect 257068 241538 257120 241544
rect 256884 240032 256936 240038
rect 256884 239974 256936 239980
rect 257264 239737 257292 248386
rect 257342 240816 257398 240825
rect 257342 240751 257398 240760
rect 257250 239728 257306 239737
rect 257250 239663 257306 239672
rect 256792 239284 256844 239290
rect 256792 239226 256844 239232
rect 256804 235249 256832 239226
rect 256790 235240 256846 235249
rect 256790 235175 256846 235184
rect 256700 207052 256752 207058
rect 256700 206994 256752 207000
rect 256054 153096 256110 153105
rect 256054 153031 256110 153040
rect 256712 89729 256740 206994
rect 257356 201482 257384 240751
rect 258092 213217 258120 276791
rect 258262 270600 258318 270609
rect 258262 270535 258264 270544
rect 258316 270535 258318 270544
rect 258264 270506 258316 270512
rect 258724 269068 258776 269074
rect 258724 269010 258776 269016
rect 258172 258120 258224 258126
rect 258172 258062 258224 258068
rect 258184 255270 258212 258062
rect 258172 255264 258224 255270
rect 258172 255206 258224 255212
rect 258540 253224 258592 253230
rect 258540 253166 258592 253172
rect 258264 251864 258316 251870
rect 258264 251806 258316 251812
rect 258172 247104 258224 247110
rect 258172 247046 258224 247052
rect 258184 224330 258212 247046
rect 258276 241097 258304 251806
rect 258552 251569 258580 253166
rect 258538 251560 258594 251569
rect 258538 251495 258594 251504
rect 258262 241088 258318 241097
rect 258262 241023 258318 241032
rect 258172 224324 258224 224330
rect 258172 224266 258224 224272
rect 258078 213208 258134 213217
rect 258078 213143 258134 213152
rect 258736 212537 258764 269010
rect 258828 268938 258856 280871
rect 259550 277264 259606 277273
rect 259550 277199 259606 277208
rect 259458 273184 259514 273193
rect 259458 273119 259460 273128
rect 259512 273119 259514 273128
rect 259460 273090 259512 273096
rect 259368 269816 259420 269822
rect 259368 269758 259420 269764
rect 259380 269006 259408 269758
rect 259368 269000 259420 269006
rect 259368 268942 259420 268948
rect 258816 268932 258868 268938
rect 258816 268874 258868 268880
rect 259274 265568 259330 265577
rect 259274 265503 259330 265512
rect 259288 263294 259316 265503
rect 259276 263288 259328 263294
rect 259276 263230 259328 263236
rect 258816 260908 258868 260914
rect 258816 260850 258868 260856
rect 258828 257446 258856 260850
rect 258816 257440 258868 257446
rect 258816 257382 258868 257388
rect 258816 227112 258868 227118
rect 258816 227054 258868 227060
rect 258722 212528 258778 212537
rect 258722 212463 258778 212472
rect 257344 201476 257396 201482
rect 257344 201418 257396 201424
rect 258724 141432 258776 141438
rect 258724 141374 258776 141380
rect 256698 89720 256754 89729
rect 256698 89655 256754 89664
rect 256056 84856 256108 84862
rect 256056 84798 256108 84804
rect 255964 9036 256016 9042
rect 255964 8978 256016 8984
rect 256068 6186 256096 84798
rect 256700 17332 256752 17338
rect 256700 17274 256752 17280
rect 254676 6180 254728 6186
rect 254676 6122 254728 6128
rect 256056 6180 256108 6186
rect 256056 6122 256108 6128
rect 253480 3460 253532 3466
rect 253480 3402 253532 3408
rect 253204 3392 253256 3398
rect 253204 3334 253256 3340
rect 253492 480 253520 3402
rect 254688 480 254716 6122
rect 255872 3528 255924 3534
rect 255872 3470 255924 3476
rect 255884 480 255912 3470
rect 256712 490 256740 17274
rect 258264 8968 258316 8974
rect 258264 8910 258316 8916
rect 256896 598 257108 626
rect 256896 490 256924 598
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 256712 462 256924 490
rect 257080 480 257108 598
rect 258276 480 258304 8910
rect 258736 3058 258764 141374
rect 258828 102814 258856 227054
rect 259472 153202 259500 273090
rect 259564 212566 259592 277199
rect 259734 265704 259790 265713
rect 259734 265639 259790 265648
rect 259644 245812 259696 245818
rect 259644 245754 259696 245760
rect 259656 215966 259684 245754
rect 259748 240961 259776 265639
rect 260746 259448 260802 259457
rect 260746 259383 260748 259392
rect 260800 259383 260802 259392
rect 260748 259354 260800 259360
rect 259734 240952 259790 240961
rect 259734 240887 259790 240896
rect 260852 229770 260880 302262
rect 260944 273873 260972 359450
rect 262312 337408 262364 337414
rect 262312 337350 262364 337356
rect 261024 322992 261076 322998
rect 261024 322934 261076 322940
rect 261036 288318 261064 322934
rect 261114 312488 261170 312497
rect 261114 312423 261170 312432
rect 261024 288312 261076 288318
rect 261024 288254 261076 288260
rect 261128 278730 261156 312423
rect 262220 307080 262272 307086
rect 262220 307022 262272 307028
rect 262232 286958 262260 307022
rect 262220 286952 262272 286958
rect 262220 286894 262272 286900
rect 261116 278724 261168 278730
rect 261116 278666 261168 278672
rect 262324 277273 262352 337350
rect 262876 313993 262904 449890
rect 263612 320113 263640 450191
rect 267740 446412 267792 446418
rect 267740 446354 267792 446360
rect 263692 437504 263744 437510
rect 263692 437446 263744 437452
rect 263598 320104 263654 320113
rect 263598 320039 263654 320048
rect 263704 318889 263732 437446
rect 265072 434648 265124 434654
rect 265072 434590 265124 434596
rect 264980 427848 265032 427854
rect 264980 427790 265032 427796
rect 263784 417512 263836 417518
rect 263784 417454 263836 417460
rect 263796 416838 263824 417454
rect 263784 416832 263836 416838
rect 263784 416774 263836 416780
rect 263796 386345 263824 416774
rect 263782 386336 263838 386345
rect 263782 386271 263838 386280
rect 263876 322244 263928 322250
rect 263876 322186 263928 322192
rect 263782 320104 263838 320113
rect 263782 320039 263838 320048
rect 263796 319025 263824 320039
rect 263782 319016 263838 319025
rect 263782 318951 263838 318960
rect 263690 318880 263746 318889
rect 263690 318815 263746 318824
rect 262862 313984 262918 313993
rect 262862 313919 262918 313928
rect 262404 311976 262456 311982
rect 262404 311918 262456 311924
rect 262416 302234 262444 311918
rect 262864 309800 262916 309806
rect 262864 309742 262916 309748
rect 262876 304366 262904 309742
rect 262864 304360 262916 304366
rect 262864 304302 262916 304308
rect 262416 302206 262536 302234
rect 262404 298240 262456 298246
rect 262404 298182 262456 298188
rect 262416 293282 262444 298182
rect 262508 296682 262536 302206
rect 262496 296676 262548 296682
rect 262496 296618 262548 296624
rect 262496 295044 262548 295050
rect 262496 294986 262548 294992
rect 262404 293276 262456 293282
rect 262404 293218 262456 293224
rect 262508 292574 262536 294986
rect 262416 292546 262536 292574
rect 262310 277264 262366 277273
rect 262310 277199 262366 277208
rect 260930 273864 260986 273873
rect 260930 273799 260986 273808
rect 261024 270564 261076 270570
rect 261024 270506 261076 270512
rect 260932 266416 260984 266422
rect 260932 266358 260984 266364
rect 260840 229764 260892 229770
rect 260840 229706 260892 229712
rect 260944 227050 260972 266358
rect 261036 231810 261064 270506
rect 261116 256760 261168 256766
rect 261116 256702 261168 256708
rect 261128 238134 261156 256702
rect 262312 250504 262364 250510
rect 262312 250446 262364 250452
rect 262324 249830 262352 250446
rect 262312 249824 262364 249830
rect 262312 249766 262364 249772
rect 261116 238128 261168 238134
rect 261116 238070 261168 238076
rect 261024 231804 261076 231810
rect 261024 231746 261076 231752
rect 260932 227044 260984 227050
rect 260932 226986 260984 226992
rect 259644 215960 259696 215966
rect 259644 215902 259696 215908
rect 259552 212560 259604 212566
rect 259552 212502 259604 212508
rect 259460 153196 259512 153202
rect 259460 153138 259512 153144
rect 259564 108322 259592 212502
rect 260104 147688 260156 147694
rect 260104 147630 260156 147636
rect 259552 108316 259604 108322
rect 259552 108258 259604 108264
rect 258816 102808 258868 102814
rect 258816 102750 258868 102756
rect 259550 86184 259606 86193
rect 259550 86119 259606 86128
rect 259564 6914 259592 86119
rect 259472 6886 259592 6914
rect 258724 3052 258776 3058
rect 258724 2994 258776 3000
rect 259472 480 259500 6886
rect 260116 3534 260144 147630
rect 261036 116618 261064 231746
rect 262324 207641 262352 249766
rect 262416 243574 262444 292546
rect 263598 290728 263654 290737
rect 263598 290663 263654 290672
rect 262588 290556 262640 290562
rect 262588 290498 262640 290504
rect 262496 264988 262548 264994
rect 262496 264930 262548 264936
rect 262404 243568 262456 243574
rect 262404 243510 262456 243516
rect 262508 237318 262536 264930
rect 262496 237312 262548 237318
rect 262496 237254 262548 237260
rect 262310 207632 262366 207641
rect 262310 207567 262366 207576
rect 262600 204950 262628 290498
rect 262678 247888 262734 247897
rect 262678 247823 262734 247832
rect 262692 247722 262720 247823
rect 262680 247716 262732 247722
rect 262680 247658 262732 247664
rect 262864 228404 262916 228410
rect 262864 228346 262916 228352
rect 262220 204944 262272 204950
rect 262220 204886 262272 204892
rect 262588 204944 262640 204950
rect 262588 204886 262640 204892
rect 261024 116612 261076 116618
rect 261024 116554 261076 116560
rect 262232 94761 262260 204886
rect 262218 94752 262274 94761
rect 262218 94687 262274 94696
rect 262876 77178 262904 228346
rect 262864 77172 262916 77178
rect 262864 77114 262916 77120
rect 262218 76528 262274 76537
rect 262218 76463 262274 76472
rect 260840 26920 260892 26926
rect 260840 26862 260892 26868
rect 260852 16574 260880 26862
rect 262232 16574 262260 76463
rect 260852 16546 261800 16574
rect 262232 16546 262536 16574
rect 260104 3528 260156 3534
rect 260104 3470 260156 3476
rect 260656 3052 260708 3058
rect 260656 2994 260708 3000
rect 260668 480 260696 2994
rect 261772 480 261800 16546
rect 262508 490 262536 16546
rect 263612 6254 263640 290663
rect 263704 285569 263732 318815
rect 263690 285560 263746 285569
rect 263690 285495 263746 285504
rect 263704 284374 263732 285495
rect 263692 284368 263744 284374
rect 263692 284310 263744 284316
rect 263690 277944 263746 277953
rect 263690 277879 263746 277888
rect 263704 277574 263732 277879
rect 263692 277568 263744 277574
rect 263692 277510 263744 277516
rect 263704 209778 263732 277510
rect 263796 270881 263824 318951
rect 263888 288289 263916 322186
rect 264992 309806 265020 427790
rect 265084 318782 265112 434590
rect 266360 424380 266412 424386
rect 266360 424322 266412 424328
rect 265164 329180 265216 329186
rect 265164 329122 265216 329128
rect 265072 318776 265124 318782
rect 265072 318718 265124 318724
rect 264980 309800 265032 309806
rect 264980 309742 265032 309748
rect 265070 305688 265126 305697
rect 265070 305623 265126 305632
rect 264886 296984 264942 296993
rect 264886 296919 264942 296928
rect 264900 291922 264928 296919
rect 264888 291916 264940 291922
rect 264888 291858 264940 291864
rect 263874 288280 263930 288289
rect 263874 288215 263930 288224
rect 264888 284368 264940 284374
rect 264940 284316 265020 284322
rect 264888 284310 265020 284316
rect 264900 284294 265020 284310
rect 263782 270872 263838 270881
rect 263782 270807 263838 270816
rect 263874 263800 263930 263809
rect 263874 263735 263930 263744
rect 263784 257372 263836 257378
rect 263784 257314 263836 257320
rect 263796 256086 263824 257314
rect 263784 256080 263836 256086
rect 263784 256022 263836 256028
rect 263692 209772 263744 209778
rect 263692 209714 263744 209720
rect 263704 109750 263732 209714
rect 263796 191146 263824 256022
rect 263888 225622 263916 263735
rect 263876 225616 263928 225622
rect 263876 225558 263928 225564
rect 263784 191140 263836 191146
rect 263784 191082 263836 191088
rect 264992 146946 265020 284294
rect 265084 270502 265112 305623
rect 265176 274582 265204 329122
rect 265256 321632 265308 321638
rect 265256 321574 265308 321580
rect 265268 288386 265296 321574
rect 265348 318776 265400 318782
rect 265348 318718 265400 318724
rect 265360 317558 265388 318718
rect 265348 317552 265400 317558
rect 265348 317494 265400 317500
rect 265256 288380 265308 288386
rect 265256 288322 265308 288328
rect 265360 285433 265388 317494
rect 266372 311030 266400 424322
rect 266452 419552 266504 419558
rect 266452 419494 266504 419500
rect 266464 387705 266492 419494
rect 266450 387696 266506 387705
rect 266450 387631 266506 387640
rect 266450 339552 266506 339561
rect 266450 339487 266452 339496
rect 266504 339487 266506 339496
rect 266452 339458 266504 339464
rect 266452 326460 266504 326466
rect 266452 326402 266504 326408
rect 266360 311024 266412 311030
rect 266360 310966 266412 310972
rect 266358 298072 266414 298081
rect 266358 298007 266414 298016
rect 266372 297498 266400 298007
rect 266360 297492 266412 297498
rect 266360 297434 266412 297440
rect 265346 285424 265402 285433
rect 265346 285359 265402 285368
rect 265360 284345 265388 285359
rect 265346 284336 265402 284345
rect 265346 284271 265402 284280
rect 266358 284336 266414 284345
rect 266464 284306 266492 326402
rect 266544 313336 266596 313342
rect 266544 313278 266596 313284
rect 266358 284271 266414 284280
rect 266452 284300 266504 284306
rect 265164 274576 265216 274582
rect 265164 274518 265216 274524
rect 265072 270496 265124 270502
rect 265072 270438 265124 270444
rect 265164 262880 265216 262886
rect 265164 262822 265216 262828
rect 265070 258904 265126 258913
rect 265070 258839 265126 258848
rect 265084 258641 265112 258839
rect 265070 258632 265126 258641
rect 265070 258567 265126 258576
rect 265084 189689 265112 258567
rect 265176 236706 265204 262822
rect 265622 242856 265678 242865
rect 265622 242791 265678 242800
rect 265164 236700 265216 236706
rect 265164 236642 265216 236648
rect 265636 224262 265664 242791
rect 265624 224256 265676 224262
rect 265624 224198 265676 224204
rect 265070 189680 265126 189689
rect 265070 189615 265126 189624
rect 264980 146940 265032 146946
rect 264980 146882 265032 146888
rect 266372 131102 266400 284271
rect 266452 284242 266504 284248
rect 266556 284238 266584 313278
rect 266636 311024 266688 311030
rect 266636 310966 266688 310972
rect 266648 310554 266676 310966
rect 266636 310548 266688 310554
rect 266636 310490 266688 310496
rect 266544 284232 266596 284238
rect 266544 284174 266596 284180
rect 266450 283520 266506 283529
rect 266450 283455 266506 283464
rect 266464 207670 266492 283455
rect 266648 278361 266676 310490
rect 267752 309369 267780 446354
rect 267832 387116 267884 387122
rect 267832 387058 267884 387064
rect 267738 309360 267794 309369
rect 267738 309295 267794 309304
rect 266634 278352 266690 278361
rect 266634 278287 266690 278296
rect 267752 272241 267780 309295
rect 267844 289814 267872 387058
rect 268016 314696 268068 314702
rect 268016 314638 268068 314644
rect 267922 308408 267978 308417
rect 267922 308343 267978 308352
rect 267936 291825 267964 308343
rect 267922 291816 267978 291825
rect 267922 291751 267978 291760
rect 267832 289808 267884 289814
rect 267832 289750 267884 289756
rect 267832 284300 267884 284306
rect 267832 284242 267884 284248
rect 267738 272232 267794 272241
rect 267738 272167 267794 272176
rect 266818 267064 266874 267073
rect 266818 266999 266820 267008
rect 266872 266999 266874 267008
rect 267648 267028 267700 267034
rect 266820 266970 266872 266976
rect 267648 266970 267700 266976
rect 267660 266370 267688 266970
rect 267660 266342 267780 266370
rect 267186 264888 267242 264897
rect 267186 264823 267242 264832
rect 267200 263634 267228 264823
rect 266544 263628 266596 263634
rect 266544 263570 266596 263576
rect 267188 263628 267240 263634
rect 267188 263570 267240 263576
rect 266452 207664 266504 207670
rect 266452 207606 266504 207612
rect 266360 131096 266412 131102
rect 266360 131038 266412 131044
rect 263692 109744 263744 109750
rect 263692 109686 263744 109692
rect 266464 95946 266492 207606
rect 266556 192506 266584 263570
rect 266910 255232 266966 255241
rect 266910 255167 266966 255176
rect 266924 253978 266952 255167
rect 266636 253972 266688 253978
rect 266636 253914 266688 253920
rect 266912 253972 266964 253978
rect 266912 253914 266964 253920
rect 266648 227089 266676 253914
rect 266634 227080 266690 227089
rect 266634 227015 266690 227024
rect 266544 192500 266596 192506
rect 266544 192442 266596 192448
rect 267752 166326 267780 266342
rect 267844 214606 267872 284242
rect 267832 214600 267884 214606
rect 267832 214542 267884 214548
rect 267740 166320 267792 166326
rect 267740 166262 267792 166268
rect 267844 104174 267872 214542
rect 267936 211818 267964 291751
rect 268028 282878 268056 314638
rect 269132 309097 269160 452610
rect 270500 450016 270552 450022
rect 270500 449958 270552 449964
rect 269304 378208 269356 378214
rect 269304 378150 269356 378156
rect 269118 309088 269174 309097
rect 269118 309023 269174 309032
rect 269118 305008 269174 305017
rect 269118 304943 269174 304952
rect 269132 295361 269160 304943
rect 269118 295352 269174 295361
rect 269118 295287 269174 295296
rect 269120 294024 269172 294030
rect 269120 293966 269172 293972
rect 268016 282872 268068 282878
rect 268016 282814 268068 282820
rect 268014 268016 268070 268025
rect 268014 267951 268070 267960
rect 268028 234598 268056 267951
rect 269028 249076 269080 249082
rect 269028 249018 269080 249024
rect 269040 248470 269068 249018
rect 269028 248464 269080 248470
rect 269026 248432 269028 248441
rect 269080 248432 269082 248441
rect 269026 248367 269082 248376
rect 268016 234592 268068 234598
rect 268016 234534 268068 234540
rect 267924 211812 267976 211818
rect 267924 211754 267976 211760
rect 267924 122120 267976 122126
rect 267924 122062 267976 122068
rect 267832 104168 267884 104174
rect 267832 104110 267884 104116
rect 266452 95940 266504 95946
rect 266452 95882 266504 95888
rect 267004 83564 267056 83570
rect 267004 83506 267056 83512
rect 266360 69692 266412 69698
rect 266360 69634 266412 69640
rect 264980 21412 265032 21418
rect 264980 21354 265032 21360
rect 263600 6248 263652 6254
rect 263600 6190 263652 6196
rect 264152 3392 264204 3398
rect 264152 3334 264204 3340
rect 262784 598 262996 626
rect 262784 490 262812 598
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262508 462 262812 490
rect 262968 480 262996 598
rect 264164 480 264192 3334
rect 264992 490 265020 21354
rect 266372 16574 266400 69634
rect 266372 16546 266584 16574
rect 265176 598 265388 626
rect 265176 490 265204 598
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 264992 462 265204 490
rect 265360 480 265388 598
rect 266556 480 266584 16546
rect 267016 3466 267044 83506
rect 267936 16574 267964 122062
rect 269132 75857 269160 293966
rect 269212 288448 269264 288454
rect 269212 288390 269264 288396
rect 269224 92585 269252 288390
rect 269316 277574 269344 378150
rect 270512 320210 270540 449958
rect 270592 429888 270644 429894
rect 270592 429830 270644 429836
rect 270604 321609 270632 429830
rect 271156 417518 271184 702850
rect 273352 455456 273404 455462
rect 273352 455398 273404 455404
rect 271880 442264 271932 442270
rect 271880 442206 271932 442212
rect 271144 417512 271196 417518
rect 271144 417454 271196 417460
rect 270684 338156 270736 338162
rect 270684 338098 270736 338104
rect 270590 321600 270646 321609
rect 270590 321535 270646 321544
rect 270500 320204 270552 320210
rect 270500 320146 270552 320152
rect 269394 309088 269450 309097
rect 269394 309023 269450 309032
rect 269408 307873 269436 309023
rect 269394 307864 269450 307873
rect 269394 307799 269450 307808
rect 269304 277568 269356 277574
rect 269304 277510 269356 277516
rect 269408 277302 269436 307799
rect 270512 287065 270540 320146
rect 270604 287473 270632 321535
rect 270590 287464 270646 287473
rect 270590 287399 270646 287408
rect 270498 287056 270554 287065
rect 270498 286991 270554 287000
rect 269396 277296 269448 277302
rect 269396 277238 269448 277244
rect 269408 276078 269436 277238
rect 269396 276072 269448 276078
rect 269396 276014 269448 276020
rect 269304 274576 269356 274582
rect 269304 274518 269356 274524
rect 269316 222154 269344 274518
rect 270590 273864 270646 273873
rect 270590 273799 270646 273808
rect 270498 272232 270554 272241
rect 270498 272167 270554 272176
rect 269856 264240 269908 264246
rect 269856 264182 269908 264188
rect 269868 263673 269896 264182
rect 269854 263664 269910 263673
rect 269854 263599 269910 263608
rect 270408 253904 270460 253910
rect 270408 253846 270460 253852
rect 270420 253298 270448 253846
rect 269396 253292 269448 253298
rect 269396 253234 269448 253240
rect 270408 253292 270460 253298
rect 270408 253234 270460 253240
rect 269408 252657 269436 253234
rect 269394 252648 269450 252657
rect 269394 252583 269450 252592
rect 270408 251864 270460 251870
rect 270408 251806 270460 251812
rect 270420 251258 270448 251806
rect 269396 251252 269448 251258
rect 269396 251194 269448 251200
rect 270408 251252 270460 251258
rect 270408 251194 270460 251200
rect 269408 233238 269436 251194
rect 269396 233232 269448 233238
rect 269396 233174 269448 233180
rect 269304 222148 269356 222154
rect 269304 222090 269356 222096
rect 270512 151745 270540 272167
rect 270604 209846 270632 273799
rect 270696 271862 270724 338098
rect 271892 320657 271920 442206
rect 271972 393372 272024 393378
rect 271972 393314 272024 393320
rect 271984 360874 272012 393314
rect 271972 360868 272024 360874
rect 271972 360810 272024 360816
rect 271878 320648 271934 320657
rect 271878 320583 271934 320592
rect 270774 289096 270830 289105
rect 270774 289031 270830 289040
rect 270684 271856 270736 271862
rect 270684 271798 270736 271804
rect 270682 259584 270738 259593
rect 270682 259519 270738 259528
rect 270696 259486 270724 259519
rect 270684 259480 270736 259486
rect 270684 259422 270736 259428
rect 270682 254416 270738 254425
rect 270682 254351 270738 254360
rect 270696 238066 270724 254351
rect 270684 238060 270736 238066
rect 270684 238002 270736 238008
rect 270788 228410 270816 289031
rect 271880 276072 271932 276078
rect 271880 276014 271932 276020
rect 271788 260772 271840 260778
rect 271788 260714 271840 260720
rect 271800 259486 271828 260714
rect 271788 259480 271840 259486
rect 271788 259422 271840 259428
rect 270776 228404 270828 228410
rect 270776 228346 270828 228352
rect 270592 209840 270644 209846
rect 270592 209782 270644 209788
rect 270498 151736 270554 151745
rect 270498 151671 270554 151680
rect 270604 97481 270632 209782
rect 271892 149054 271920 276014
rect 271984 276010 272012 360810
rect 272154 320648 272210 320657
rect 272154 320583 272210 320592
rect 272168 320249 272196 320583
rect 272154 320240 272210 320249
rect 272154 320175 272210 320184
rect 272062 298072 272118 298081
rect 272062 298007 272118 298016
rect 271972 276004 272024 276010
rect 271972 275946 272024 275952
rect 271970 251152 272026 251161
rect 271970 251087 272026 251096
rect 271984 250617 272012 251087
rect 271970 250608 272026 250617
rect 271970 250543 272026 250552
rect 271984 204270 272012 250543
rect 272076 235278 272104 298007
rect 272168 265577 272196 320175
rect 272524 319456 272576 319462
rect 272524 319398 272576 319404
rect 272536 299470 272564 319398
rect 273258 299568 273314 299577
rect 273258 299503 273314 299512
rect 272524 299464 272576 299470
rect 272522 299432 272524 299441
rect 272576 299432 272578 299441
rect 272522 299367 272578 299376
rect 272536 299341 272564 299367
rect 272154 265568 272210 265577
rect 272154 265503 272210 265512
rect 272154 250744 272210 250753
rect 272154 250679 272210 250688
rect 272064 235272 272116 235278
rect 272064 235214 272116 235220
rect 272168 217938 272196 250679
rect 272156 217932 272208 217938
rect 272156 217874 272208 217880
rect 271972 204264 272024 204270
rect 271972 204206 272024 204212
rect 271880 149048 271932 149054
rect 271880 148990 271932 148996
rect 271788 105596 271840 105602
rect 271788 105538 271840 105544
rect 271800 104922 271828 105538
rect 271788 104916 271840 104922
rect 271788 104858 271840 104864
rect 270590 97472 270646 97481
rect 270590 97407 270646 97416
rect 269210 92576 269266 92585
rect 269210 92511 269266 92520
rect 269118 75848 269174 75857
rect 269118 75783 269174 75792
rect 269120 58676 269172 58682
rect 269120 58618 269172 58624
rect 269132 16574 269160 58618
rect 270500 53100 270552 53106
rect 270500 53042 270552 53048
rect 270512 16574 270540 53042
rect 267936 16546 268424 16574
rect 269132 16546 269988 16574
rect 270512 16546 270816 16574
rect 267740 3528 267792 3534
rect 267740 3470 267792 3476
rect 267004 3460 267056 3466
rect 267004 3402 267056 3408
rect 267752 480 267780 3470
rect 268396 490 268424 16546
rect 269960 2666 269988 16546
rect 270040 4820 270092 4826
rect 270040 4762 270092 4768
rect 270052 2854 270080 4762
rect 270040 2848 270092 2854
rect 270040 2790 270092 2796
rect 269960 2638 270080 2666
rect 268672 598 268884 626
rect 268672 490 268700 598
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268396 462 268700 490
rect 268856 480 268884 598
rect 270052 480 270080 2638
rect 270788 490 270816 16546
rect 271800 9654 271828 104858
rect 273272 56574 273300 299503
rect 273364 245614 273392 455398
rect 273916 389094 273944 703258
rect 282184 703044 282236 703050
rect 282184 702986 282236 702992
rect 280804 702704 280856 702710
rect 280804 702646 280856 702652
rect 276020 454164 276072 454170
rect 276020 454106 276072 454112
rect 274640 435396 274692 435402
rect 274640 435338 274692 435344
rect 273904 389088 273956 389094
rect 273904 389030 273956 389036
rect 273536 382288 273588 382294
rect 273536 382230 273588 382236
rect 273444 380928 273496 380934
rect 273444 380870 273496 380876
rect 273456 274650 273484 380870
rect 273548 277370 273576 382230
rect 273536 277364 273588 277370
rect 273536 277306 273588 277312
rect 273444 274644 273496 274650
rect 273444 274586 273496 274592
rect 274652 274582 274680 435338
rect 274732 405748 274784 405754
rect 274732 405690 274784 405696
rect 274744 369850 274772 405690
rect 274732 369844 274784 369850
rect 274732 369786 274784 369792
rect 274744 280090 274772 369786
rect 274824 332716 274876 332722
rect 274824 332658 274876 332664
rect 274836 290494 274864 332658
rect 274824 290488 274876 290494
rect 274824 290430 274876 290436
rect 274824 289808 274876 289814
rect 274824 289750 274876 289756
rect 274732 280084 274784 280090
rect 274732 280026 274784 280032
rect 273904 274576 273956 274582
rect 273904 274518 273956 274524
rect 274640 274576 274692 274582
rect 274640 274518 274692 274524
rect 273534 255640 273590 255649
rect 273534 255575 273590 255584
rect 273352 245608 273404 245614
rect 273352 245550 273404 245556
rect 273364 244934 273392 245550
rect 273352 244928 273404 244934
rect 273352 244870 273404 244876
rect 273352 244316 273404 244322
rect 273352 244258 273404 244264
rect 273364 234569 273392 244258
rect 273444 241460 273496 241466
rect 273444 241402 273496 241408
rect 273350 234560 273406 234569
rect 273350 234495 273406 234504
rect 273364 78577 273392 234495
rect 273456 133210 273484 241402
rect 273548 220289 273576 255575
rect 273916 241466 273944 274518
rect 273904 241460 273956 241466
rect 273904 241402 273956 241408
rect 274836 227118 274864 289750
rect 274914 280800 274970 280809
rect 274914 280735 274970 280744
rect 274824 227112 274876 227118
rect 274824 227054 274876 227060
rect 273534 220280 273590 220289
rect 273534 220215 273590 220224
rect 274928 209774 274956 280735
rect 276032 262886 276060 454106
rect 277400 451308 277452 451314
rect 277400 451250 277452 451256
rect 276112 422340 276164 422346
rect 276112 422282 276164 422288
rect 276124 321570 276152 422282
rect 276204 408536 276256 408542
rect 276204 408478 276256 408484
rect 276216 380905 276244 408478
rect 276202 380896 276258 380905
rect 276202 380831 276258 380840
rect 276216 379545 276244 380831
rect 276202 379536 276258 379545
rect 276202 379471 276258 379480
rect 276112 321564 276164 321570
rect 276112 321506 276164 321512
rect 276124 287026 276152 321506
rect 276296 306400 276348 306406
rect 276296 306342 276348 306348
rect 276112 287020 276164 287026
rect 276112 286962 276164 286968
rect 276202 277944 276258 277953
rect 276202 277879 276258 277888
rect 276020 262880 276072 262886
rect 276020 262822 276072 262828
rect 274652 209746 274956 209774
rect 274652 206310 274680 209746
rect 274640 206304 274692 206310
rect 274640 206246 274692 206252
rect 274652 162178 274680 206246
rect 274640 162172 274692 162178
rect 274640 162114 274692 162120
rect 276018 135960 276074 135969
rect 276018 135895 276074 135904
rect 273444 133204 273496 133210
rect 273444 133146 273496 133152
rect 273350 78568 273406 78577
rect 273350 78503 273406 78512
rect 273260 56568 273312 56574
rect 273260 56510 273312 56516
rect 273272 55894 273300 56510
rect 273260 55888 273312 55894
rect 273260 55830 273312 55836
rect 274640 51740 274692 51746
rect 274640 51682 274692 51688
rect 274652 16574 274680 51682
rect 276032 16574 276060 135895
rect 276216 125594 276244 277879
rect 276308 186998 276336 306342
rect 276388 295996 276440 296002
rect 276388 295938 276440 295944
rect 276296 186992 276348 186998
rect 276296 186934 276348 186940
rect 276400 129742 276428 295938
rect 277412 268433 277440 451250
rect 279332 427100 279384 427106
rect 279332 427042 279384 427048
rect 279344 426494 279372 427042
rect 279332 426488 279384 426494
rect 279332 426430 279384 426436
rect 279344 422294 279372 426430
rect 279344 422266 279464 422294
rect 277492 400240 277544 400246
rect 277492 400182 277544 400188
rect 277504 376582 277532 400182
rect 277492 376576 277544 376582
rect 277492 376518 277544 376524
rect 277504 269822 277532 376518
rect 278872 324964 278924 324970
rect 278872 324906 278924 324912
rect 277584 316056 277636 316062
rect 277584 315998 277636 316004
rect 277596 282169 277624 315998
rect 277674 306504 277730 306513
rect 277674 306439 277730 306448
rect 277582 282160 277638 282169
rect 277582 282095 277638 282104
rect 277492 269816 277544 269822
rect 277492 269758 277544 269764
rect 277398 268424 277454 268433
rect 277398 268359 277454 268368
rect 277398 266792 277454 266801
rect 277398 266727 277454 266736
rect 277412 230450 277440 266727
rect 277584 253224 277636 253230
rect 277584 253166 277636 253172
rect 277400 230444 277452 230450
rect 277400 230386 277452 230392
rect 276388 129736 276440 129742
rect 276388 129678 276440 129684
rect 276204 125588 276256 125594
rect 276204 125530 276256 125536
rect 277412 115326 277440 230386
rect 277492 220108 277544 220114
rect 277492 220050 277544 220056
rect 277400 115320 277452 115326
rect 277400 115262 277452 115268
rect 277504 113150 277532 220050
rect 277596 160750 277624 253166
rect 277688 220114 277716 306439
rect 278778 302424 278834 302433
rect 278778 302359 278834 302368
rect 278136 262268 278188 262274
rect 278136 262210 278188 262216
rect 278044 259412 278096 259418
rect 278044 259354 278096 259360
rect 278056 249762 278084 259354
rect 278148 258777 278176 262210
rect 278134 258768 278190 258777
rect 278134 258703 278190 258712
rect 278148 253230 278176 258703
rect 278136 253224 278188 253230
rect 278136 253166 278188 253172
rect 278044 249756 278096 249762
rect 278044 249698 278096 249704
rect 277676 220108 277728 220114
rect 277676 220050 277728 220056
rect 277584 160744 277636 160750
rect 277584 160686 277636 160692
rect 278792 135250 278820 302359
rect 278884 295225 278912 324906
rect 278964 311908 279016 311914
rect 278964 311850 279016 311856
rect 278870 295216 278926 295225
rect 278870 295151 278926 295160
rect 278884 294001 278912 295151
rect 278870 293992 278926 294001
rect 278870 293927 278926 293936
rect 278870 287464 278926 287473
rect 278870 287399 278926 287408
rect 278884 146305 278912 287399
rect 278976 280158 279004 311850
rect 278964 280152 279016 280158
rect 278964 280094 279016 280100
rect 278962 254552 279018 254561
rect 278962 254487 279018 254496
rect 278976 231130 279004 254487
rect 279436 253162 279464 422266
rect 280160 420980 280212 420986
rect 280160 420922 280212 420928
rect 279424 253156 279476 253162
rect 279424 253098 279476 253104
rect 280172 246362 280200 420922
rect 280436 324352 280488 324358
rect 280436 324294 280488 324300
rect 280250 311264 280306 311273
rect 280250 311199 280306 311208
rect 280264 250510 280292 311199
rect 280342 311128 280398 311137
rect 280342 311063 280398 311072
rect 280356 260846 280384 311063
rect 280448 296721 280476 324294
rect 280816 311137 280844 702646
rect 281632 448996 281684 449002
rect 281632 448938 281684 448944
rect 281446 311264 281502 311273
rect 281446 311199 281502 311208
rect 281460 311166 281488 311199
rect 281448 311160 281500 311166
rect 280802 311128 280858 311137
rect 281448 311102 281500 311108
rect 280802 311063 280858 311072
rect 280434 296712 280490 296721
rect 280434 296647 280490 296656
rect 280448 295361 280476 296647
rect 280434 295352 280490 295361
rect 280434 295287 280490 295296
rect 281540 293276 281592 293282
rect 281540 293218 281592 293224
rect 280804 291916 280856 291922
rect 280804 291858 280856 291864
rect 280344 260840 280396 260846
rect 280344 260782 280396 260788
rect 280252 250504 280304 250510
rect 280252 250446 280304 250452
rect 280160 246356 280212 246362
rect 280160 246298 280212 246304
rect 278964 231124 279016 231130
rect 278964 231066 279016 231072
rect 278870 146296 278926 146305
rect 278870 146231 278926 146240
rect 278780 135244 278832 135250
rect 278780 135186 278832 135192
rect 280068 135244 280120 135250
rect 280068 135186 280120 135192
rect 280080 134570 280108 135186
rect 280068 134564 280120 134570
rect 280068 134506 280120 134512
rect 278044 129736 278096 129742
rect 278044 129678 278096 129684
rect 277492 113144 277544 113150
rect 277492 113086 277544 113092
rect 278056 102814 278084 129678
rect 280172 124166 280200 246298
rect 280816 132462 280844 291858
rect 280896 142180 280948 142186
rect 280896 142122 280948 142128
rect 280804 132456 280856 132462
rect 280804 132398 280856 132404
rect 280816 131782 280844 132398
rect 280804 131776 280856 131782
rect 280804 131718 280856 131724
rect 280160 124160 280212 124166
rect 280160 124102 280212 124108
rect 278688 113144 278740 113150
rect 278688 113086 278740 113092
rect 278700 112470 278728 113086
rect 278688 112464 278740 112470
rect 278688 112406 278740 112412
rect 278044 102808 278096 102814
rect 278044 102750 278096 102756
rect 277400 94512 277452 94518
rect 277400 94454 277452 94460
rect 277412 16574 277440 94454
rect 280804 57248 280856 57254
rect 280804 57190 280856 57196
rect 278780 29640 278832 29646
rect 278780 29582 278832 29588
rect 278792 16574 278820 29582
rect 274652 16546 274864 16574
rect 276032 16546 276704 16574
rect 277412 16546 278360 16574
rect 278792 16546 279096 16574
rect 271788 9648 271840 9654
rect 271788 9590 271840 9596
rect 273628 3460 273680 3466
rect 273628 3402 273680 3408
rect 272432 2848 272484 2854
rect 272432 2790 272484 2796
rect 271064 598 271276 626
rect 271064 490 271092 598
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 270788 462 271092 490
rect 271248 480 271276 598
rect 272444 480 272472 2790
rect 273640 480 273668 3402
rect 274836 480 274864 16546
rect 276020 9648 276072 9654
rect 276020 9590 276072 9596
rect 276032 480 276060 9590
rect 276676 490 276704 16546
rect 276952 598 277164 626
rect 276952 490 276980 598
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 276676 462 276980 490
rect 277136 480 277164 598
rect 278332 480 278360 16546
rect 279068 490 279096 16546
rect 280712 15904 280764 15910
rect 280712 15846 280764 15852
rect 279344 598 279556 626
rect 279344 490 279372 598
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279068 462 279372 490
rect 279528 480 279556 598
rect 280724 480 280752 15846
rect 280816 3534 280844 57190
rect 280908 33794 280936 142122
rect 281552 82793 281580 293218
rect 281644 259418 281672 448938
rect 282196 388385 282224 702986
rect 300136 702982 300164 703520
rect 332520 703186 332548 703520
rect 348804 703322 348832 703520
rect 348792 703316 348844 703322
rect 348792 703258 348844 703264
rect 364996 703254 365024 703520
rect 364984 703248 365036 703254
rect 364984 703190 365036 703196
rect 332508 703180 332560 703186
rect 332508 703122 332560 703128
rect 300124 702976 300176 702982
rect 300124 702918 300176 702924
rect 397472 702778 397500 703520
rect 413664 703118 413692 703520
rect 413652 703112 413704 703118
rect 413652 703054 413704 703060
rect 429856 702846 429884 703520
rect 462332 703050 462360 703520
rect 462320 703044 462372 703050
rect 462320 702986 462372 702992
rect 478524 702914 478552 703520
rect 478512 702908 478564 702914
rect 478512 702850 478564 702856
rect 429844 702840 429896 702846
rect 429844 702782 429896 702788
rect 397460 702772 397512 702778
rect 397460 702714 397512 702720
rect 494808 702506 494836 703520
rect 527192 702658 527220 703520
rect 543476 702710 543504 703520
rect 527100 702642 527220 702658
rect 543464 702704 543516 702710
rect 543464 702646 543516 702652
rect 527088 702636 527220 702642
rect 527140 702630 527220 702636
rect 527088 702578 527140 702584
rect 559668 702545 559696 703520
rect 580908 702568 580960 702574
rect 559654 702536 559710 702545
rect 494796 702500 494848 702506
rect 580908 702510 580960 702516
rect 559654 702471 559710 702480
rect 494796 702442 494848 702448
rect 580920 697241 580948 702510
rect 580906 697232 580962 697241
rect 580906 697167 580962 697176
rect 582378 683904 582434 683913
rect 582378 683839 582434 683848
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 291200 462392 291252 462398
rect 291200 462334 291252 462340
rect 285680 461644 285732 461650
rect 285680 461586 285732 461592
rect 285692 460970 285720 461586
rect 285680 460964 285732 460970
rect 285732 460912 285904 460934
rect 285680 460906 285904 460912
rect 284390 458416 284446 458425
rect 284390 458351 284446 458360
rect 284300 443692 284352 443698
rect 284300 443634 284352 443640
rect 283012 432608 283064 432614
rect 283012 432550 283064 432556
rect 282182 388376 282238 388385
rect 282182 388311 282238 388320
rect 281724 385076 281776 385082
rect 281724 385018 281776 385024
rect 281736 273222 281764 385018
rect 282920 382968 282972 382974
rect 282918 382936 282920 382945
rect 282972 382936 282974 382945
rect 282918 382871 282974 382880
rect 281816 342916 281868 342922
rect 281816 342858 281868 342864
rect 281724 273216 281776 273222
rect 281724 273158 281776 273164
rect 281722 271144 281778 271153
rect 281722 271079 281778 271088
rect 281632 259412 281684 259418
rect 281632 259354 281684 259360
rect 281632 253156 281684 253162
rect 281632 253098 281684 253104
rect 281644 126954 281672 253098
rect 281736 150414 281764 271079
rect 281828 244254 281856 342858
rect 282918 303648 282974 303657
rect 282918 303583 282974 303592
rect 281816 244248 281868 244254
rect 281816 244190 281868 244196
rect 281724 150408 281776 150414
rect 281724 150350 281776 150356
rect 281632 126948 281684 126954
rect 281632 126890 281684 126896
rect 282184 120760 282236 120766
rect 282184 120702 282236 120708
rect 281538 82784 281594 82793
rect 281538 82719 281594 82728
rect 281552 82142 281580 82719
rect 281540 82136 281592 82142
rect 281540 82078 281592 82084
rect 280896 33788 280948 33794
rect 280896 33730 280948 33736
rect 281540 13116 281592 13122
rect 281540 13058 281592 13064
rect 280804 3528 280856 3534
rect 280804 3470 280856 3476
rect 281552 490 281580 13058
rect 282196 2990 282224 120702
rect 282932 73166 282960 303583
rect 283024 247761 283052 432550
rect 283104 382968 283156 382974
rect 283104 382910 283156 382916
rect 283116 255649 283144 382910
rect 283102 255640 283158 255649
rect 283102 255575 283158 255584
rect 283010 247752 283066 247761
rect 283010 247687 283066 247696
rect 283024 225690 283052 247687
rect 284312 239426 284340 443634
rect 284404 262274 284432 458351
rect 285680 418192 285732 418198
rect 285680 418134 285732 418140
rect 285692 386345 285720 418134
rect 285678 386336 285734 386345
rect 285678 386271 285734 386280
rect 284574 367704 284630 367713
rect 284574 367639 284630 367648
rect 284482 295352 284538 295361
rect 284482 295287 284538 295296
rect 284392 262268 284444 262274
rect 284392 262210 284444 262216
rect 284390 242856 284446 242865
rect 284390 242791 284446 242800
rect 284404 242185 284432 242791
rect 284390 242176 284446 242185
rect 284390 242111 284446 242120
rect 284300 239420 284352 239426
rect 284300 239362 284352 239368
rect 283012 225684 283064 225690
rect 283012 225626 283064 225632
rect 284404 88097 284432 242111
rect 284496 163441 284524 295287
rect 284588 242865 284616 367639
rect 285772 298172 285824 298178
rect 285772 298114 285824 298120
rect 285678 293992 285734 294001
rect 285678 293927 285734 293936
rect 284668 262200 284720 262206
rect 284668 262142 284720 262148
rect 284680 260914 284708 262142
rect 284668 260908 284720 260914
rect 284668 260850 284720 260856
rect 284574 242856 284630 242865
rect 284574 242791 284630 242800
rect 284680 233209 284708 260850
rect 284666 233200 284722 233209
rect 284666 233135 284722 233144
rect 284482 163432 284538 163441
rect 284482 163367 284538 163376
rect 284390 88088 284446 88097
rect 284390 88023 284446 88032
rect 284300 79348 284352 79354
rect 284300 79290 284352 79296
rect 282920 73160 282972 73166
rect 282920 73102 282972 73108
rect 282932 72486 282960 73102
rect 282920 72480 282972 72486
rect 282920 72422 282972 72428
rect 282184 2984 282236 2990
rect 282184 2926 282236 2932
rect 283104 2984 283156 2990
rect 283104 2926 283156 2932
rect 281736 598 281948 626
rect 281736 490 281764 598
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281552 462 281764 490
rect 281920 480 281948 598
rect 283116 480 283144 2926
rect 284312 480 284340 79290
rect 285692 60625 285720 293927
rect 285784 67590 285812 298114
rect 285876 257378 285904 460906
rect 287058 456920 287114 456929
rect 287058 456855 287114 456864
rect 288346 456920 288402 456929
rect 288346 456855 288402 456864
rect 286048 418804 286100 418810
rect 286048 418746 286100 418752
rect 286060 418198 286088 418746
rect 286048 418192 286100 418198
rect 286048 418134 286100 418140
rect 287072 258126 287100 456855
rect 288360 456822 288388 456855
rect 288348 456816 288400 456822
rect 288348 456758 288400 456764
rect 288438 453112 288494 453121
rect 288438 453047 288494 453056
rect 287150 451344 287206 451353
rect 287150 451279 287206 451288
rect 285956 258120 286008 258126
rect 285956 258062 286008 258068
rect 287060 258120 287112 258126
rect 287060 258062 287112 258068
rect 285864 257372 285916 257378
rect 285864 257314 285916 257320
rect 285968 146985 285996 258062
rect 287164 253910 287192 451279
rect 287336 309800 287388 309806
rect 287336 309742 287388 309748
rect 287244 297424 287296 297430
rect 287244 297366 287296 297372
rect 287152 253904 287204 253910
rect 287152 253846 287204 253852
rect 285954 146976 286010 146985
rect 285954 146911 286010 146920
rect 287256 103514 287284 297366
rect 287348 126886 287376 309742
rect 287704 256012 287756 256018
rect 287704 255954 287756 255960
rect 287716 159390 287744 255954
rect 288452 219434 288480 453047
rect 288624 439544 288676 439550
rect 288624 439486 288676 439492
rect 288532 299600 288584 299606
rect 288532 299542 288584 299548
rect 288440 219428 288492 219434
rect 288440 219370 288492 219376
rect 288452 219201 288480 219370
rect 288438 219192 288494 219201
rect 288438 219127 288494 219136
rect 287704 159384 287756 159390
rect 287704 159326 287756 159332
rect 287336 126880 287388 126886
rect 287336 126822 287388 126828
rect 288348 126880 288400 126886
rect 288348 126822 288400 126828
rect 288360 126274 288388 126822
rect 288348 126268 288400 126274
rect 288348 126210 288400 126216
rect 288544 107642 288572 299542
rect 288636 256018 288664 439486
rect 289728 399492 289780 399498
rect 289728 399434 289780 399440
rect 289740 398886 289768 399434
rect 288716 398880 288768 398886
rect 288716 398822 288768 398828
rect 289728 398880 289780 398886
rect 289728 398822 289780 398828
rect 288728 262206 288756 398822
rect 291108 398132 291160 398138
rect 291108 398074 291160 398080
rect 291120 397526 291148 398074
rect 289820 397520 289872 397526
rect 289820 397462 289872 397468
rect 291108 397520 291160 397526
rect 291108 397462 291160 397468
rect 289832 367033 289860 397462
rect 289818 367024 289874 367033
rect 289818 366959 289874 366968
rect 289832 364334 289860 366959
rect 289832 364306 289952 364334
rect 289820 299532 289872 299538
rect 289820 299474 289872 299480
rect 288716 262200 288768 262206
rect 288716 262142 288768 262148
rect 288624 256012 288676 256018
rect 288624 255954 288676 255960
rect 288624 244248 288676 244254
rect 288624 244190 288676 244196
rect 288532 107636 288584 107642
rect 288532 107578 288584 107584
rect 287072 103486 287284 103514
rect 287072 102134 287100 103486
rect 287060 102128 287112 102134
rect 287060 102070 287112 102076
rect 288348 102128 288400 102134
rect 288348 102070 288400 102076
rect 288360 101454 288388 102070
rect 288348 101448 288400 101454
rect 288348 101390 288400 101396
rect 288636 86873 288664 244190
rect 289084 140820 289136 140826
rect 289084 140762 289136 140768
rect 288622 86864 288678 86873
rect 288622 86799 288678 86808
rect 288438 71088 288494 71097
rect 288438 71023 288494 71032
rect 285772 67584 285824 67590
rect 285772 67526 285824 67532
rect 285784 66910 285812 67526
rect 285772 66904 285824 66910
rect 285772 66846 285824 66852
rect 285678 60616 285734 60625
rect 285678 60551 285734 60560
rect 286414 60616 286470 60625
rect 286414 60551 286470 60560
rect 286428 60042 286456 60551
rect 286416 60036 286468 60042
rect 286416 59978 286468 59984
rect 285680 40724 285732 40730
rect 285680 40666 285732 40672
rect 284392 19984 284444 19990
rect 284392 19926 284444 19932
rect 284404 16574 284432 19926
rect 285692 16574 285720 40666
rect 288452 16574 288480 71023
rect 284404 16546 284984 16574
rect 285692 16546 286640 16574
rect 288452 16546 289032 16574
rect 284956 490 284984 16546
rect 285232 598 285444 626
rect 285232 490 285260 598
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 284956 462 285260 490
rect 285416 480 285444 598
rect 286612 480 286640 16546
rect 287796 3528 287848 3534
rect 287796 3470 287848 3476
rect 287808 480 287836 3470
rect 289004 480 289032 16546
rect 289096 3330 289124 140762
rect 289728 107636 289780 107642
rect 289728 107578 289780 107584
rect 289740 106962 289768 107578
rect 289728 106956 289780 106962
rect 289728 106898 289780 106904
rect 289726 86864 289782 86873
rect 289726 86799 289782 86808
rect 289740 85649 289768 86799
rect 289726 85640 289782 85649
rect 289726 85575 289782 85584
rect 289832 64802 289860 299474
rect 289924 260778 289952 364306
rect 291212 291922 291240 462334
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456822 580212 458079
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 582392 437442 582420 683839
rect 582654 670712 582710 670721
rect 582654 670647 582710 670656
rect 582470 644056 582526 644065
rect 582470 643991 582526 644000
rect 582380 437436 582432 437442
rect 582380 437378 582432 437384
rect 582378 431624 582434 431633
rect 582378 431559 582434 431568
rect 291292 376780 291344 376786
rect 291292 376722 291344 376728
rect 291200 291916 291252 291922
rect 291200 291858 291252 291864
rect 291304 270502 291332 376722
rect 582392 376689 582420 431559
rect 582484 398138 582512 643991
rect 582562 630864 582618 630873
rect 582562 630799 582618 630808
rect 582472 398132 582524 398138
rect 582472 398074 582524 398080
rect 582576 390561 582604 630799
rect 582668 458833 582696 670647
rect 582838 617536 582894 617545
rect 582838 617471 582894 617480
rect 582746 591016 582802 591025
rect 582746 590951 582802 590960
rect 582654 458824 582710 458833
rect 582654 458759 582710 458768
rect 582656 426488 582708 426494
rect 582656 426430 582708 426436
rect 582562 390552 582618 390561
rect 582562 390487 582618 390496
rect 582470 383888 582526 383897
rect 582470 383823 582526 383832
rect 582484 378457 582512 383823
rect 582470 378448 582526 378457
rect 582470 378383 582526 378392
rect 582378 376680 582434 376689
rect 582378 376615 582434 376624
rect 582378 365120 582434 365129
rect 582378 365055 582434 365064
rect 293960 362228 294012 362234
rect 293960 362170 294012 362176
rect 291384 331900 291436 331906
rect 291384 331842 291436 331848
rect 291292 270496 291344 270502
rect 291292 270438 291344 270444
rect 291396 266354 291424 331842
rect 291476 291848 291528 291854
rect 291476 291790 291528 291796
rect 291384 266348 291436 266354
rect 291384 266290 291436 266296
rect 289912 260772 289964 260778
rect 289912 260714 289964 260720
rect 291292 244928 291344 244934
rect 291292 244870 291344 244876
rect 291304 158710 291332 244870
rect 291292 158704 291344 158710
rect 291292 158646 291344 158652
rect 291304 158030 291332 158646
rect 291292 158024 291344 158030
rect 291292 157966 291344 157972
rect 291488 105602 291516 291790
rect 291660 270496 291712 270502
rect 291660 270438 291712 270444
rect 291672 269793 291700 270438
rect 291658 269784 291714 269793
rect 291658 269719 291714 269728
rect 293972 269074 294000 362170
rect 580262 325272 580318 325281
rect 580262 325207 580318 325216
rect 580276 311166 580304 325207
rect 580264 311160 580316 311166
rect 580264 311102 580316 311108
rect 295432 304292 295484 304298
rect 295432 304234 295484 304240
rect 293960 269068 294012 269074
rect 293960 269010 294012 269016
rect 295340 153264 295392 153270
rect 295340 153206 295392 153212
rect 291844 111104 291896 111110
rect 291844 111046 291896 111052
rect 291476 105596 291528 105602
rect 291476 105538 291528 105544
rect 289820 64796 289872 64802
rect 289820 64738 289872 64744
rect 289832 64190 289860 64738
rect 289820 64184 289872 64190
rect 289820 64126 289872 64132
rect 289820 42084 289872 42090
rect 289820 42026 289872 42032
rect 289084 3324 289136 3330
rect 289084 3266 289136 3272
rect 289832 490 289860 42026
rect 291200 36576 291252 36582
rect 291200 36518 291252 36524
rect 291212 16574 291240 36518
rect 291212 16546 291424 16574
rect 290016 598 290228 626
rect 290016 490 290044 598
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 289832 462 290044 490
rect 290200 480 290228 598
rect 291396 480 291424 16546
rect 291856 4486 291884 111046
rect 292672 60036 292724 60042
rect 292672 59978 292724 59984
rect 292684 16574 292712 59978
rect 295352 16574 295380 153206
rect 295444 144129 295472 304234
rect 580172 299464 580224 299470
rect 580172 299406 580224 299412
rect 580184 298761 580212 299406
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 580184 270502 580212 272167
rect 580172 270496 580224 270502
rect 580172 270438 580224 270444
rect 580172 259412 580224 259418
rect 580172 259354 580224 259360
rect 580184 258913 580212 259354
rect 580170 258904 580226 258913
rect 580170 258839 580226 258848
rect 582392 251870 582420 365055
rect 582668 351937 582696 426430
rect 582760 399498 582788 590951
rect 582852 585818 582880 617471
rect 582840 585812 582892 585818
rect 582840 585754 582892 585760
rect 582930 564360 582986 564369
rect 582930 564295 582986 564304
rect 582838 524512 582894 524521
rect 582838 524447 582894 524456
rect 582748 399492 582800 399498
rect 582748 399434 582800 399440
rect 582852 382974 582880 524447
rect 582944 439550 582972 564295
rect 583022 537840 583078 537849
rect 583022 537775 583078 537784
rect 582932 439544 582984 439550
rect 582932 439486 582984 439492
rect 583036 418810 583064 537775
rect 583206 511320 583262 511329
rect 583206 511255 583262 511264
rect 583114 471472 583170 471481
rect 583114 471407 583170 471416
rect 583024 418804 583076 418810
rect 583024 418746 583076 418752
rect 582930 418296 582986 418305
rect 582930 418231 582986 418240
rect 582840 382968 582892 382974
rect 582840 382910 582892 382916
rect 582944 379506 582972 418231
rect 583128 417450 583156 471407
rect 583220 461650 583248 511255
rect 583208 461644 583260 461650
rect 583208 461586 583260 461592
rect 583206 451344 583262 451353
rect 583206 451279 583262 451288
rect 583116 417444 583168 417450
rect 583116 417386 583168 417392
rect 583220 404977 583248 451279
rect 583206 404968 583262 404977
rect 583206 404903 583262 404912
rect 582932 379500 582984 379506
rect 582932 379442 582984 379448
rect 582654 351928 582710 351937
rect 582654 351863 582710 351872
rect 582562 312080 582618 312089
rect 582562 312015 582618 312024
rect 582470 302288 582526 302297
rect 582470 302223 582526 302232
rect 582380 251864 582432 251870
rect 582380 251806 582432 251812
rect 582380 248464 582432 248470
rect 582380 248406 582432 248412
rect 582392 245585 582420 248406
rect 582378 245576 582434 245585
rect 582378 245511 582434 245520
rect 580172 232552 580224 232558
rect 580172 232494 580224 232500
rect 580184 232393 580212 232494
rect 580170 232384 580226 232393
rect 580170 232319 580226 232328
rect 580264 225616 580316 225622
rect 580264 225558 580316 225564
rect 579896 219428 579948 219434
rect 579896 219370 579948 219376
rect 579908 219065 579936 219370
rect 579894 219056 579950 219065
rect 579894 218991 579950 219000
rect 580276 205737 580304 225558
rect 582378 215928 582434 215937
rect 582378 215863 582434 215872
rect 580262 205728 580318 205737
rect 580262 205663 580318 205672
rect 580172 194608 580224 194614
rect 580172 194550 580224 194556
rect 574744 193860 574796 193866
rect 574744 193802 574796 193808
rect 317420 171148 317472 171154
rect 317420 171090 317472 171096
rect 300124 164348 300176 164354
rect 300124 164290 300176 164296
rect 295430 144120 295486 144129
rect 295430 144055 295486 144064
rect 298100 124908 298152 124914
rect 298100 124850 298152 124856
rect 292684 16546 293264 16574
rect 295352 16546 295656 16574
rect 292488 6180 292540 6186
rect 292488 6122 292540 6128
rect 291844 4480 291896 4486
rect 291844 4422 291896 4428
rect 292500 2990 292528 6122
rect 292580 3324 292632 3330
rect 292580 3266 292632 3272
rect 292488 2984 292540 2990
rect 292488 2926 292540 2932
rect 292592 480 292620 3266
rect 293236 490 293264 16546
rect 294880 2984 294932 2990
rect 294880 2926 294932 2932
rect 293512 598 293724 626
rect 293512 490 293540 598
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293236 462 293540 490
rect 293696 480 293724 598
rect 294892 480 294920 2926
rect 295628 490 295656 16546
rect 297272 4480 297324 4486
rect 297272 4422 297324 4428
rect 295904 598 296116 626
rect 295904 490 295932 598
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 295628 462 295932 490
rect 296088 480 296116 598
rect 297284 480 297312 4422
rect 298112 490 298140 124850
rect 299480 102808 299532 102814
rect 299480 102750 299532 102756
rect 299492 3534 299520 102750
rect 300136 5642 300164 164290
rect 303618 163432 303674 163441
rect 303618 163367 303674 163376
rect 302238 144120 302294 144129
rect 302238 144055 302294 144064
rect 301962 7576 302018 7585
rect 301962 7511 302018 7520
rect 300124 5636 300176 5642
rect 300124 5578 300176 5584
rect 299480 3528 299532 3534
rect 299480 3470 299532 3476
rect 300768 3528 300820 3534
rect 300768 3470 300820 3476
rect 299664 3120 299716 3126
rect 299664 3062 299716 3068
rect 298296 598 298508 626
rect 298296 490 298324 598
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298112 462 298324 490
rect 298480 480 298508 598
rect 299676 480 299704 3062
rect 300780 480 300808 3470
rect 301976 480 302004 7511
rect 302252 3126 302280 144055
rect 303632 16574 303660 163367
rect 316040 138780 316092 138786
rect 316040 138722 316092 138728
rect 307024 134564 307076 134570
rect 307024 134506 307076 134512
rect 305644 131776 305696 131782
rect 305644 131718 305696 131724
rect 304264 115252 304316 115258
rect 304264 115194 304316 115200
rect 303632 16546 303936 16574
rect 303160 14476 303212 14482
rect 303160 14418 303212 14424
rect 302424 9036 302476 9042
rect 302424 8978 302476 8984
rect 302436 3534 302464 8978
rect 302424 3528 302476 3534
rect 302424 3470 302476 3476
rect 302240 3120 302292 3126
rect 302240 3062 302292 3068
rect 303172 480 303200 14418
rect 303908 490 303936 16546
rect 304276 3058 304304 115194
rect 305656 6225 305684 131718
rect 305736 39364 305788 39370
rect 305736 39306 305788 39312
rect 305642 6216 305698 6225
rect 305642 6151 305698 6160
rect 305748 5574 305776 39306
rect 306748 5636 306800 5642
rect 306748 5578 306800 5584
rect 305736 5568 305788 5574
rect 305736 5510 305788 5516
rect 305552 3528 305604 3534
rect 305552 3470 305604 3476
rect 304264 3052 304316 3058
rect 304264 2994 304316 3000
rect 304184 598 304396 626
rect 304184 490 304212 598
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 303908 462 304212 490
rect 304368 480 304396 598
rect 305564 480 305592 3470
rect 306760 480 306788 5578
rect 307036 4214 307064 134506
rect 313280 119400 313332 119406
rect 313280 119342 313332 119348
rect 309782 84280 309838 84289
rect 309782 84215 309838 84224
rect 309140 68332 309192 68338
rect 309140 68274 309192 68280
rect 309152 6914 309180 68274
rect 309796 16574 309824 84215
rect 313292 16574 313320 119342
rect 316052 16574 316080 138722
rect 317432 16574 317460 171090
rect 335358 155272 335414 155281
rect 335358 155207 335414 155216
rect 331864 127628 331916 127634
rect 331864 127570 331916 127576
rect 324320 112464 324372 112470
rect 324320 112406 324372 112412
rect 323584 103556 323636 103562
rect 323584 103498 323636 103504
rect 321652 101448 321704 101454
rect 321652 101390 321704 101396
rect 320824 100020 320876 100026
rect 320824 99962 320876 99968
rect 320180 66904 320232 66910
rect 320180 66846 320232 66852
rect 320192 16574 320220 66846
rect 309796 16546 309916 16574
rect 313292 16546 313872 16574
rect 316052 16546 316264 16574
rect 317432 16546 318104 16574
rect 320192 16546 320496 16574
rect 309152 6886 309824 6914
rect 309048 5568 309100 5574
rect 309048 5510 309100 5516
rect 307024 4208 307076 4214
rect 307024 4150 307076 4156
rect 307944 3052 307996 3058
rect 307944 2994 307996 3000
rect 307956 480 307984 2994
rect 309060 480 309088 5510
rect 309796 490 309824 6886
rect 309888 3398 309916 16546
rect 312176 11756 312228 11762
rect 312176 11698 312228 11704
rect 309876 3392 309928 3398
rect 309876 3334 309928 3340
rect 311440 3392 311492 3398
rect 311440 3334 311492 3340
rect 310072 598 310284 626
rect 310072 490 310100 598
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 309796 462 310100 490
rect 310256 480 310284 598
rect 311452 480 311480 3334
rect 312188 490 312216 11698
rect 312464 598 312676 626
rect 312464 490 312492 598
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312188 462 312492 490
rect 312648 480 312676 598
rect 313844 480 313872 16546
rect 315028 4208 315080 4214
rect 315028 4150 315080 4156
rect 315040 480 315068 4150
rect 316236 480 316264 16546
rect 317328 3256 317380 3262
rect 317328 3198 317380 3204
rect 317340 480 317368 3198
rect 318076 490 318104 16546
rect 319718 6216 319774 6225
rect 319718 6151 319774 6160
rect 318352 598 318564 626
rect 318352 490 318380 598
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 462 318380 490
rect 318536 480 318564 598
rect 319732 480 319760 6151
rect 320468 490 320496 16546
rect 320836 3466 320864 99962
rect 321560 17264 321612 17270
rect 321560 17206 321612 17212
rect 320824 3460 320876 3466
rect 320824 3402 320876 3408
rect 321572 3074 321600 17206
rect 321664 3262 321692 101390
rect 322940 82136 322992 82142
rect 322940 82078 322992 82084
rect 321652 3256 321704 3262
rect 321652 3198 321704 3204
rect 321572 3046 322152 3074
rect 320744 598 320956 626
rect 320744 490 320772 598
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320468 462 320772 490
rect 320928 480 320956 598
rect 322124 480 322152 3046
rect 322952 490 322980 82078
rect 323596 4826 323624 103498
rect 323584 4820 323636 4826
rect 323584 4762 323636 4768
rect 324332 3534 324360 112406
rect 327078 80744 327134 80753
rect 327078 80679 327134 80688
rect 325700 33788 325752 33794
rect 325700 33730 325752 33736
rect 324412 25560 324464 25566
rect 324412 25502 324464 25508
rect 324320 3528 324372 3534
rect 324320 3470 324372 3476
rect 323136 598 323348 626
rect 323136 490 323164 598
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 322952 462 323164 490
rect 323320 480 323348 598
rect 324424 480 324452 25502
rect 325712 16574 325740 33730
rect 327092 16574 327120 80679
rect 328460 28280 328512 28286
rect 328460 28222 328512 28228
rect 328472 16574 328500 28222
rect 331220 24132 331272 24138
rect 331220 24074 331272 24080
rect 325712 16546 326384 16574
rect 327092 16546 328040 16574
rect 328472 16546 328776 16574
rect 325608 3528 325660 3534
rect 325608 3470 325660 3476
rect 325620 480 325648 3470
rect 326356 490 326384 16546
rect 326632 598 326844 626
rect 326632 490 326660 598
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326356 462 326660 490
rect 326816 480 326844 598
rect 328012 480 328040 16546
rect 328748 490 328776 16546
rect 330392 4820 330444 4826
rect 330392 4762 330444 4768
rect 329024 598 329236 626
rect 329024 490 329052 598
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 328748 462 329052 490
rect 329208 480 329236 598
rect 330404 480 330432 4762
rect 331232 490 331260 24074
rect 331876 4554 331904 127570
rect 333980 72480 334032 72486
rect 333980 72422 334032 72428
rect 332692 37936 332744 37942
rect 332692 37878 332744 37884
rect 332704 11762 332732 37878
rect 333992 16574 334020 72422
rect 335372 16574 335400 155207
rect 340144 145580 340196 145586
rect 340144 145522 340196 145528
rect 338120 47592 338172 47598
rect 338120 47534 338172 47540
rect 338132 16574 338160 47534
rect 333992 16546 334664 16574
rect 335372 16546 336320 16574
rect 338132 16546 338712 16574
rect 332692 11756 332744 11762
rect 332692 11698 332744 11704
rect 333888 11756 333940 11762
rect 333888 11698 333940 11704
rect 331864 4548 331916 4554
rect 331864 4490 331916 4496
rect 332692 3460 332744 3466
rect 332692 3402 332744 3408
rect 331416 598 331628 626
rect 331416 490 331444 598
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331232 462 331444 490
rect 331600 480 331628 598
rect 332704 480 332732 3402
rect 333900 480 333928 11698
rect 334636 490 334664 16546
rect 334716 10328 334768 10334
rect 334716 10270 334768 10276
rect 334728 3466 334756 10270
rect 334716 3460 334768 3466
rect 334716 3402 334768 3408
rect 334912 598 335124 626
rect 334912 490 334940 598
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 462 334940 490
rect 335096 480 335124 598
rect 336292 480 336320 16546
rect 337476 4548 337528 4554
rect 337476 4490 337528 4496
rect 337488 480 337516 4490
rect 338684 480 338712 16546
rect 340156 3534 340184 145522
rect 353300 126268 353352 126274
rect 353300 126210 353352 126216
rect 342904 106956 342956 106962
rect 342904 106898 342956 106904
rect 340972 55888 341024 55894
rect 340972 55830 341024 55836
rect 340236 35216 340288 35222
rect 340236 35158 340288 35164
rect 340144 3528 340196 3534
rect 340144 3470 340196 3476
rect 339868 3460 339920 3466
rect 339868 3402 339920 3408
rect 339880 480 339908 3402
rect 340248 3330 340276 35158
rect 340236 3324 340288 3330
rect 340236 3266 340288 3272
rect 340984 480 341012 55830
rect 342260 31068 342312 31074
rect 342260 31010 342312 31016
rect 342272 6914 342300 31010
rect 342916 16574 342944 106898
rect 345020 64184 345072 64190
rect 345020 64126 345072 64132
rect 344284 18624 344336 18630
rect 344284 18566 344336 18572
rect 342916 16546 343036 16574
rect 342272 6886 342944 6914
rect 342168 3528 342220 3534
rect 342168 3470 342220 3476
rect 342180 480 342208 3470
rect 342916 490 342944 6886
rect 343008 4146 343036 16546
rect 342996 4140 343048 4146
rect 342996 4082 343048 4088
rect 344296 3466 344324 18566
rect 345032 16574 345060 64126
rect 349804 43444 349856 43450
rect 349804 43386 349856 43392
rect 347044 22772 347096 22778
rect 347044 22714 347096 22720
rect 345032 16546 345336 16574
rect 344284 3460 344336 3466
rect 344284 3402 344336 3408
rect 344560 3324 344612 3330
rect 344560 3266 344612 3272
rect 343192 598 343404 626
rect 343192 490 343220 598
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 462 343220 490
rect 343376 480 343404 598
rect 344572 480 344600 3266
rect 345308 490 345336 16546
rect 346952 4140 347004 4146
rect 346952 4082 347004 4088
rect 345584 598 345796 626
rect 345584 490 345612 598
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345308 462 345612 490
rect 345768 480 345796 598
rect 346964 480 346992 4082
rect 347056 3126 347084 22714
rect 349816 5574 349844 43386
rect 349804 5568 349856 5574
rect 349804 5510 349856 5516
rect 351644 5568 351696 5574
rect 351644 5510 351696 5516
rect 348054 3496 348110 3505
rect 348054 3431 348110 3440
rect 350448 3460 350500 3466
rect 347044 3120 347096 3126
rect 347044 3062 347096 3068
rect 348068 480 348096 3431
rect 350448 3402 350500 3408
rect 349252 3120 349304 3126
rect 349252 3062 349304 3068
rect 349264 480 349292 3062
rect 350460 480 350488 3402
rect 351656 480 351684 5510
rect 353312 3505 353340 126210
rect 353298 3496 353354 3505
rect 574756 3466 574784 193802
rect 580184 192545 580212 194550
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580184 178702 580212 179143
rect 580172 178696 580224 178702
rect 580172 178638 580224 178644
rect 580262 89040 580318 89049
rect 580262 88975 580318 88984
rect 580276 73001 580304 88975
rect 580262 72992 580318 73001
rect 580262 72927 580318 72936
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 353298 3431 353354 3440
rect 574744 3460 574796 3466
rect 574744 3402 574796 3408
rect 582196 3460 582248 3466
rect 582196 3402 582248 3408
rect 581000 3256 581052 3262
rect 581000 3198 581052 3204
rect 581012 480 581040 3198
rect 582208 480 582236 3402
rect 582392 3074 582420 215863
rect 582484 3262 582512 302223
rect 582576 250481 582604 312015
rect 582562 250472 582618 250481
rect 582562 250407 582618 250416
rect 582564 240780 582616 240786
rect 582564 240722 582616 240728
rect 582576 152697 582604 240722
rect 582748 170400 582800 170406
rect 582748 170342 582800 170348
rect 582656 156664 582708 156670
rect 582656 156606 582708 156612
rect 582562 152688 582618 152697
rect 582562 152623 582618 152632
rect 582564 138712 582616 138718
rect 582564 138654 582616 138660
rect 582576 19825 582604 138654
rect 582668 112849 582696 156606
rect 582760 139369 582788 170342
rect 582838 165880 582894 165889
rect 582838 165815 582894 165824
rect 582746 139360 582802 139369
rect 582746 139295 582802 139304
rect 582852 124166 582880 165815
rect 582932 158024 582984 158030
rect 582932 157966 582984 157972
rect 582944 126041 582972 157966
rect 583022 140856 583078 140865
rect 583022 140791 583078 140800
rect 582930 126032 582986 126041
rect 582930 125967 582986 125976
rect 582840 124160 582892 124166
rect 582840 124102 582892 124108
rect 582654 112840 582710 112849
rect 582654 112775 582710 112784
rect 582654 99512 582710 99521
rect 582654 99447 582710 99456
rect 582668 78577 582696 99447
rect 582930 87544 582986 87553
rect 582930 87479 582986 87488
rect 582840 83496 582892 83502
rect 582840 83438 582892 83444
rect 582654 78568 582710 78577
rect 582654 78503 582710 78512
rect 582852 33153 582880 83438
rect 582838 33144 582894 33153
rect 582838 33079 582894 33088
rect 582562 19816 582618 19825
rect 582562 19751 582618 19760
rect 582944 6633 582972 87479
rect 583036 59673 583064 140791
rect 583022 59664 583078 59673
rect 583022 59599 583078 59608
rect 582930 6624 582986 6633
rect 582930 6559 582986 6568
rect 582472 3256 582524 3262
rect 582472 3198 582524 3204
rect 582392 3046 583432 3074
rect 583404 480 583432 3046
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3514 671200 3570 671256
rect 3422 658144 3478 658200
rect 3422 632032 3478 632088
rect 2778 606056 2834 606112
rect 3514 619112 3570 619168
rect 8114 581032 8170 581088
rect 3514 579944 3570 580000
rect 3422 566888 3478 566944
rect 3330 553832 3386 553888
rect 14462 541048 14518 541104
rect 3514 527876 3570 527912
rect 3514 527856 3516 527876
rect 3516 527856 3568 527876
rect 3568 527856 3570 527876
rect 3514 514820 3570 514856
rect 3514 514800 3516 514820
rect 3516 514800 3568 514820
rect 3568 514800 3570 514820
rect 3422 501744 3478 501800
rect 2778 475632 2834 475688
rect 3146 449520 3202 449576
rect 2962 410488 3018 410544
rect 3514 462576 3570 462632
rect 3514 423580 3516 423600
rect 3516 423580 3568 423600
rect 3568 423580 3570 423600
rect 3514 423544 3570 423580
rect 3514 397432 3570 397488
rect 3514 386280 3570 386336
rect 3422 371320 3478 371376
rect 11702 389136 11758 389192
rect 3238 358400 3294 358456
rect 3422 345364 3478 345400
rect 3422 345344 3424 345364
rect 3424 345344 3476 345364
rect 3476 345344 3478 345364
rect 4066 319232 4122 319288
rect 1306 309168 1362 309224
rect 3238 306176 3294 306232
rect 3422 293120 3478 293176
rect 3146 254088 3202 254144
rect 3514 283192 3570 283248
rect 3514 267144 3570 267200
rect 3514 241032 3570 241088
rect 6826 232464 6882 232520
rect 4066 220088 4122 220144
rect 3422 214920 3478 214976
rect 3238 201864 3294 201920
rect 3422 188808 3478 188864
rect 3422 162868 3424 162888
rect 3424 162868 3476 162888
rect 3476 162868 3478 162888
rect 3422 162832 3478 162868
rect 3330 149776 3386 149832
rect 3238 136720 3294 136776
rect 3422 110608 3478 110664
rect 3422 97552 3478 97608
rect 3146 84632 3202 84688
rect 3422 83408 3478 83464
rect 3422 71576 3478 71632
rect 2962 58520 3018 58576
rect 3422 45500 3424 45520
rect 3424 45500 3476 45520
rect 3476 45500 3478 45520
rect 3422 45464 3478 45500
rect 3514 32408 3570 32464
rect 3422 19352 3478 19408
rect 3422 6432 3478 6488
rect 10966 146920 11022 146976
rect 32402 388320 32458 388376
rect 22006 324400 22062 324456
rect 17866 307808 17922 307864
rect 16486 297336 16542 297392
rect 15106 236544 15162 236600
rect 19246 221448 19302 221504
rect 33782 314744 33838 314800
rect 22742 313248 22798 313304
rect 30286 311888 30342 311944
rect 26146 302504 26202 302560
rect 24766 233824 24822 233880
rect 23386 203496 23442 203552
rect 32402 306720 32458 306776
rect 31666 200640 31722 200696
rect 33046 152360 33102 152416
rect 34426 202136 34482 202192
rect 44086 453192 44142 453248
rect 45466 434832 45522 434888
rect 37094 214512 37150 214568
rect 41142 310528 41198 310584
rect 39946 298152 40002 298208
rect 38566 224168 38622 224224
rect 39946 235184 40002 235240
rect 41234 260072 41290 260128
rect 42706 197920 42762 197976
rect 44086 255856 44142 255912
rect 48226 399472 48282 399528
rect 46846 253952 46902 254008
rect 45466 204856 45522 204912
rect 53562 433336 53618 433392
rect 50802 261432 50858 261488
rect 49606 229744 49662 229800
rect 48226 225528 48282 225584
rect 50710 151000 50766 151056
rect 52366 255176 52422 255232
rect 52366 253952 52422 254008
rect 53470 237360 53526 237416
rect 53654 237360 53710 237416
rect 52366 209616 52422 209672
rect 53470 158752 53526 158808
rect 50894 90344 50950 90400
rect 53746 158752 53802 158808
rect 55126 391448 55182 391504
rect 57702 422184 57758 422240
rect 56414 357992 56470 358048
rect 55126 289176 55182 289232
rect 53746 148280 53802 148336
rect 55126 189624 55182 189680
rect 56414 151136 56470 151192
rect 57702 242120 57758 242176
rect 57242 136720 57298 136776
rect 60554 537376 60610 537432
rect 61750 439456 61806 439512
rect 60646 425040 60702 425096
rect 59174 389272 59230 389328
rect 60462 270680 60518 270736
rect 58622 135360 58678 135416
rect 59266 258168 59322 258224
rect 59174 138080 59230 138136
rect 61658 311072 61714 311128
rect 61842 436056 61898 436112
rect 62762 438096 62818 438152
rect 61842 311072 61898 311128
rect 61842 285640 61898 285696
rect 60646 269184 60702 269240
rect 61934 265104 61990 265160
rect 60646 167592 60702 167648
rect 61842 162832 61898 162888
rect 63406 405728 63462 405784
rect 65982 567568 66038 567624
rect 65890 550840 65946 550896
rect 65798 544040 65854 544096
rect 66534 579944 66590 580000
rect 67546 578584 67602 578640
rect 67454 577224 67510 577280
rect 66534 573144 66590 573200
rect 66534 571784 66590 571840
rect 66902 570152 66958 570208
rect 67362 568792 67418 568848
rect 66166 566752 66222 566808
rect 66534 564712 66590 564768
rect 66534 563352 66590 563408
rect 66718 560632 66774 560688
rect 66718 559272 66774 559328
rect 66718 557912 66774 557968
rect 66074 555192 66130 555248
rect 65982 522280 66038 522336
rect 66534 553696 66590 553752
rect 66534 549616 66590 549672
rect 66810 548120 66866 548176
rect 66718 545400 66774 545456
rect 67270 543360 67326 543416
rect 66442 540096 66498 540152
rect 65982 475360 66038 475416
rect 65798 438096 65854 438152
rect 63130 265104 63186 265160
rect 62118 252728 62174 252784
rect 62026 240216 62082 240272
rect 61750 81096 61806 81152
rect 63222 161608 63278 161664
rect 64602 291760 64658 291816
rect 63406 252728 63462 252784
rect 65798 433336 65854 433392
rect 65890 393388 65892 393408
rect 65892 393388 65944 393408
rect 65944 393388 65946 393408
rect 65890 393352 65946 393388
rect 66074 442992 66130 443048
rect 66074 387368 66130 387424
rect 65890 373904 65946 373960
rect 65798 288360 65854 288416
rect 64786 261432 64842 261488
rect 65890 259528 65946 259584
rect 64786 235320 64842 235376
rect 66074 288360 66130 288416
rect 66074 287272 66130 287328
rect 66258 431432 66314 431488
rect 67178 430344 67234 430400
rect 66258 428168 66314 428224
rect 66902 427352 66958 427408
rect 66626 425176 66682 425232
rect 66810 424088 66866 424144
rect 66626 423272 66682 423328
rect 66810 422220 66812 422240
rect 66812 422220 66864 422240
rect 66864 422220 66866 422240
rect 66810 422184 66866 422220
rect 66902 420008 66958 420064
rect 66810 418920 66866 418976
rect 66994 417016 67050 417072
rect 66902 415928 66958 415984
rect 66718 414840 66774 414896
rect 67270 414024 67326 414080
rect 66258 412936 66314 412992
rect 66810 411848 66866 411904
rect 66902 410760 66958 410816
rect 66810 408856 66866 408912
rect 66810 407768 66866 407824
rect 67454 418104 67510 418160
rect 67362 405592 67418 405648
rect 66902 404504 66958 404560
rect 66810 403688 66866 403744
rect 67270 401648 67326 401704
rect 66718 401512 66774 401568
rect 67178 395256 67234 395312
rect 66810 394440 66866 394496
rect 66258 392264 66314 392320
rect 67362 400424 67418 400480
rect 67178 372544 67234 372600
rect 67638 575864 67694 575920
rect 71778 585112 71834 585168
rect 73526 582528 73582 582584
rect 75366 581032 75422 581088
rect 80242 581168 80298 581224
rect 85486 582664 85542 582720
rect 82726 581032 82782 581088
rect 70858 580760 70914 580816
rect 79874 580760 79930 580816
rect 84198 580760 84254 580816
rect 92110 583752 92166 583808
rect 88890 580760 88946 580816
rect 92570 580760 92626 580816
rect 67730 575320 67786 575376
rect 95238 574776 95294 574832
rect 94686 558592 94742 558648
rect 67730 556552 67786 556608
rect 67822 552200 67878 552256
rect 94686 552200 94742 552256
rect 68926 535472 68982 535528
rect 67638 474000 67694 474056
rect 67638 418104 67694 418160
rect 67546 402600 67602 402656
rect 67546 401648 67602 401704
rect 67546 399608 67602 399664
rect 68926 471824 68982 471880
rect 68926 470600 68982 470656
rect 69662 465160 69718 465216
rect 69018 440272 69074 440328
rect 68926 437144 68982 437200
rect 68558 436192 68614 436248
rect 67822 433608 67878 433664
rect 68926 436056 68982 436112
rect 70490 442992 70546 443048
rect 71134 442992 71190 443048
rect 76746 539552 76802 539608
rect 71778 460128 71834 460184
rect 71686 442856 71742 442912
rect 71594 437144 71650 437200
rect 73802 535472 73858 535528
rect 73158 472504 73214 472560
rect 71870 436056 71926 436112
rect 72698 436056 72754 436112
rect 72606 434968 72662 435024
rect 72514 434424 72570 434480
rect 75366 444896 75422 444952
rect 80058 536016 80114 536072
rect 84014 536152 84070 536208
rect 78034 455640 78090 455696
rect 75918 439456 75974 439512
rect 75642 434560 75698 434616
rect 71134 433608 71190 433664
rect 74722 433608 74778 433664
rect 76378 433608 76434 433664
rect 87602 536016 87658 536072
rect 81346 438232 81402 438288
rect 80334 436192 80390 436248
rect 79874 433744 79930 433800
rect 81346 434832 81402 434888
rect 78218 433608 78274 433664
rect 81898 433608 81954 433664
rect 82910 439456 82966 439512
rect 82818 438096 82874 438152
rect 85762 453192 85818 453248
rect 84658 433608 84714 433664
rect 85854 435240 85910 435296
rect 94318 539688 94374 539744
rect 88522 440272 88578 440328
rect 86866 435240 86922 435296
rect 86866 434832 86922 434888
rect 93950 538872 94006 538928
rect 93398 536016 93454 536072
rect 92386 464344 92442 464400
rect 89718 436192 89774 436248
rect 92570 449928 92626 449984
rect 92478 434560 92534 434616
rect 94778 542952 94834 543008
rect 95606 567160 95662 567216
rect 95422 563624 95478 563680
rect 95146 446392 95202 446448
rect 95514 558592 95570 558648
rect 97170 578856 97226 578912
rect 97170 577496 97226 577552
rect 97906 576408 97962 576464
rect 97906 573416 97962 573472
rect 96802 572056 96858 572112
rect 97262 571376 97318 571432
rect 96710 568656 96766 568712
rect 97906 570016 97962 570072
rect 97906 568676 97962 568712
rect 97906 568656 97908 568676
rect 97908 568656 97960 568676
rect 97960 568656 97962 568676
rect 96710 565800 96766 565856
rect 97262 565800 97318 565856
rect 96618 552472 96674 552528
rect 96802 562264 96858 562320
rect 96894 560904 96950 560960
rect 96802 559544 96858 559600
rect 96802 556824 96858 556880
rect 95606 534656 95662 534712
rect 96986 555464 97042 555520
rect 96986 552744 97042 552800
rect 97906 550704 97962 550760
rect 96986 545672 97042 545728
rect 95422 523640 95478 523696
rect 97078 544312 97134 544368
rect 97170 541592 97226 541648
rect 96618 456048 96674 456104
rect 95330 440816 95386 440872
rect 99378 436464 99434 436520
rect 99746 436464 99802 436520
rect 107014 582528 107070 582584
rect 101218 436328 101274 436384
rect 104254 536152 104310 536208
rect 104438 535472 104494 535528
rect 107014 467880 107070 467936
rect 107566 467880 107622 467936
rect 106646 437008 106702 437064
rect 91466 433744 91522 433800
rect 96710 433744 96766 433800
rect 100482 433744 100538 433800
rect 85946 433608 86002 433664
rect 87234 433608 87290 433664
rect 89994 433608 90050 433664
rect 91190 433608 91246 433664
rect 92938 433608 92994 433664
rect 96342 433608 96398 433664
rect 98182 433608 98238 433664
rect 98458 433608 98514 433664
rect 99838 433608 99894 433664
rect 104714 433608 104770 433664
rect 106738 433608 106794 433664
rect 107658 436056 107714 436112
rect 111062 449112 111118 449168
rect 110418 448568 110474 448624
rect 111062 448568 111118 448624
rect 109682 437280 109738 437336
rect 108394 436056 108450 436112
rect 109038 433608 109094 433664
rect 110694 433608 110750 433664
rect 111798 433608 111854 433664
rect 68650 433064 68706 433120
rect 67822 429800 67878 429856
rect 67730 397468 67732 397488
rect 67732 397468 67784 397488
rect 67784 397468 67786 397488
rect 67730 397432 67786 397468
rect 67730 396344 67786 396400
rect 67546 391992 67602 392048
rect 67546 391176 67602 391232
rect 67546 387368 67602 387424
rect 67086 283736 67142 283792
rect 66810 282956 66812 282976
rect 66812 282956 66864 282976
rect 66864 282956 66866 282976
rect 66810 282920 66866 282956
rect 67086 282140 67088 282160
rect 67088 282140 67140 282160
rect 67140 282140 67142 282160
rect 67086 282104 67142 282140
rect 67270 281560 67326 281616
rect 66534 281424 66590 281480
rect 66902 280472 66958 280528
rect 66626 278840 66682 278896
rect 66810 278044 66866 278080
rect 66810 278024 66812 278044
rect 66812 278024 66864 278044
rect 66864 278024 66866 278044
rect 66902 276392 66958 276448
rect 66166 275576 66222 275632
rect 66074 274760 66130 274816
rect 65982 239808 66038 239864
rect 65798 226344 65854 226400
rect 65798 144880 65854 144936
rect 64694 139576 64750 139632
rect 64602 89528 64658 89584
rect 66534 273964 66590 274000
rect 66534 273944 66536 273964
rect 66536 273944 66588 273964
rect 66588 273944 66590 273964
rect 66626 272312 66682 272368
rect 66258 271496 66314 271552
rect 66902 269048 66958 269104
rect 66810 268232 66866 268288
rect 66626 267416 66682 267472
rect 66442 266600 66498 266656
rect 66810 265784 66866 265840
rect 66810 264152 66866 264208
rect 67086 263336 67142 263392
rect 66902 262520 66958 262576
rect 66258 261704 66314 261760
rect 66810 260072 66866 260128
rect 66810 258440 66866 258496
rect 66258 257896 66314 257952
rect 66626 256844 66628 256864
rect 66628 256844 66680 256864
rect 66680 256844 66682 256864
rect 66626 256808 66682 256844
rect 66810 254360 66866 254416
rect 66994 253544 67050 253600
rect 66810 251912 66866 251968
rect 66442 251096 66498 251152
rect 66810 250280 66866 250336
rect 66626 249464 66682 249520
rect 66166 248648 66222 248704
rect 66074 123800 66130 123856
rect 65982 110200 66038 110256
rect 65890 107752 65946 107808
rect 66810 244568 66866 244624
rect 66626 243752 66682 243808
rect 66810 242936 66866 242992
rect 66258 131960 66314 132016
rect 66350 131144 66406 131200
rect 66258 130600 66314 130656
rect 67362 277208 67418 277264
rect 67546 283736 67602 283792
rect 67546 279656 67602 279712
rect 67454 263336 67510 263392
rect 67454 247016 67510 247072
rect 67362 246200 67418 246256
rect 113270 436736 113326 436792
rect 113270 416744 113326 416800
rect 113178 414840 113234 414896
rect 112718 406952 112774 407008
rect 112718 401784 112774 401840
rect 72514 390904 72570 390960
rect 73986 390904 74042 390960
rect 71134 390768 71190 390824
rect 70674 388184 70730 388240
rect 71226 387776 71282 387832
rect 69662 383696 69718 383752
rect 68558 283464 68614 283520
rect 68282 281424 68338 281480
rect 68190 258712 68246 258768
rect 67178 129784 67234 129840
rect 66258 128968 66314 129024
rect 66902 127608 66958 127664
rect 66810 126828 66812 126848
rect 66812 126828 66864 126848
rect 66864 126828 66866 126848
rect 66810 126792 66866 126828
rect 66902 125976 66958 126032
rect 66810 125160 66866 125216
rect 66810 122984 66866 123040
rect 66350 122168 66406 122224
rect 66810 121388 66812 121408
rect 66812 121388 66864 121408
rect 66864 121388 66866 121408
rect 66810 121352 66866 121388
rect 66902 120536 66958 120592
rect 66810 120028 66812 120048
rect 66812 120028 66864 120048
rect 66864 120028 66866 120048
rect 66810 119992 66866 120028
rect 66902 119176 66958 119232
rect 66902 118360 66958 118416
rect 66810 117544 66866 117600
rect 66626 116184 66682 116240
rect 66810 115368 66866 115424
rect 66902 114552 66958 114608
rect 66810 113736 66866 113792
rect 66902 113192 66958 113248
rect 66902 111560 66958 111616
rect 67178 110744 67234 110800
rect 66810 109384 66866 109440
rect 66810 106936 66866 106992
rect 66626 105596 66682 105632
rect 66626 105576 66628 105596
rect 66628 105576 66680 105596
rect 66680 105576 66682 105596
rect 66810 104796 66812 104816
rect 66812 104796 66864 104816
rect 66864 104796 66866 104816
rect 66810 104760 66866 104796
rect 67270 103944 67326 104000
rect 66810 102584 66866 102640
rect 66534 101768 66590 101824
rect 66810 100952 66866 101008
rect 66718 100136 66774 100192
rect 66074 85448 66130 85504
rect 66258 99592 66314 99648
rect 67546 149116 67602 149152
rect 67546 149096 67548 149116
rect 67548 149096 67600 149116
rect 67600 149096 67602 149116
rect 72422 389000 72478 389056
rect 72974 389000 73030 389056
rect 72514 387504 72570 387560
rect 69386 283464 69442 283520
rect 74446 388864 74502 388920
rect 76654 390904 76710 390960
rect 77206 384920 77262 384976
rect 73066 356632 73122 356688
rect 72422 338136 72478 338192
rect 73066 338156 73122 338192
rect 73066 338136 73068 338156
rect 73068 338136 73120 338156
rect 73120 338136 73122 338156
rect 73066 326304 73122 326360
rect 69754 283328 69810 283384
rect 72054 287000 72110 287056
rect 71042 283056 71098 283112
rect 71318 283464 71374 283520
rect 72422 284280 72478 284336
rect 73158 289856 73214 289912
rect 73066 287000 73122 287056
rect 73158 284144 73214 284200
rect 79138 389000 79194 389056
rect 79966 389000 80022 389056
rect 77390 320184 77446 320240
rect 75182 304952 75238 305008
rect 74538 289992 74594 290048
rect 74906 284280 74962 284336
rect 75918 285776 75974 285832
rect 76010 284824 76066 284880
rect 80150 389000 80206 389056
rect 80978 389000 81034 389056
rect 79966 368328 80022 368384
rect 79966 294480 80022 294536
rect 79322 289176 79378 289232
rect 79690 289040 79746 289096
rect 82082 390632 82138 390688
rect 81254 388320 81310 388376
rect 81346 382880 81402 382936
rect 80150 291760 80206 291816
rect 80886 291216 80942 291272
rect 89258 390496 89314 390552
rect 83186 387504 83242 387560
rect 83462 369688 83518 369744
rect 86866 320728 86922 320784
rect 84842 318688 84898 318744
rect 82726 317484 82782 317520
rect 82726 317464 82728 317484
rect 82728 317464 82780 317484
rect 82780 317464 82782 317484
rect 82726 316784 82782 316840
rect 82910 312432 82966 312488
rect 83094 291896 83150 291952
rect 82634 289992 82690 290048
rect 83186 290400 83242 290456
rect 75366 283056 75422 283112
rect 83462 304952 83518 305008
rect 86222 316648 86278 316704
rect 85854 291216 85910 291272
rect 86774 291216 86830 291272
rect 89166 387504 89222 387560
rect 88982 384240 89038 384296
rect 89534 381520 89590 381576
rect 87050 300736 87106 300792
rect 86406 287408 86462 287464
rect 86866 287408 86922 287464
rect 87510 285640 87566 285696
rect 88982 307944 89038 308000
rect 87602 284144 87658 284200
rect 89534 302776 89590 302832
rect 89166 284416 89222 284472
rect 88614 283464 88670 283520
rect 91098 386960 91154 387016
rect 91006 383696 91062 383752
rect 90914 319368 90970 319424
rect 89718 300736 89774 300792
rect 90914 289856 90970 289912
rect 89626 284416 89682 284472
rect 91926 390360 91982 390416
rect 94318 388184 94374 388240
rect 94778 387912 94834 387968
rect 91098 292576 91154 292632
rect 90914 285640 90970 285696
rect 91926 285776 91982 285832
rect 83462 283328 83518 283384
rect 95146 320184 95202 320240
rect 95054 318008 95110 318064
rect 93766 294480 93822 294536
rect 93858 285640 93914 285696
rect 95330 390632 95386 390688
rect 96710 390632 96766 390688
rect 95238 304952 95294 305008
rect 104254 390632 104310 390688
rect 100942 390496 100998 390552
rect 96986 390360 97042 390416
rect 96894 389000 96950 389056
rect 97630 389000 97686 389056
rect 99470 389272 99526 389328
rect 99562 388456 99618 388512
rect 96526 305632 96582 305688
rect 97906 323584 97962 323640
rect 96618 298696 96674 298752
rect 95790 287136 95846 287192
rect 99286 319368 99342 319424
rect 97446 284280 97502 284336
rect 102046 390224 102102 390280
rect 102414 389408 102470 389464
rect 102046 389136 102102 389192
rect 101494 384240 101550 384296
rect 100758 320184 100814 320240
rect 100022 291896 100078 291952
rect 97906 283056 97962 283112
rect 85302 282920 85358 282976
rect 98918 282784 98974 282840
rect 98090 258440 98146 258496
rect 69478 241712 69534 241768
rect 72698 241712 72754 241768
rect 73250 241712 73306 241768
rect 73802 241712 73858 241768
rect 69662 241440 69718 241496
rect 70306 241440 70362 241496
rect 69202 239944 69258 240000
rect 69294 139440 69350 139496
rect 67822 132776 67878 132832
rect 67730 112376 67786 112432
rect 67730 110744 67786 110800
rect 67454 97960 67510 98016
rect 67362 97144 67418 97200
rect 66902 95784 66958 95840
rect 66810 94968 66866 95024
rect 67270 94152 67326 94208
rect 67546 92540 67602 92576
rect 67546 92520 67548 92540
rect 67548 92520 67600 92540
rect 67600 92520 67602 92540
rect 67362 86672 67418 86728
rect 67822 103128 67878 103184
rect 69570 134988 69572 135008
rect 69572 134988 69624 135008
rect 69624 134988 69626 135008
rect 69570 134952 69626 134988
rect 70812 241304 70868 241360
rect 71318 241304 71374 241360
rect 71318 240080 71374 240136
rect 72238 240080 72294 240136
rect 71686 237496 71742 237552
rect 70030 138216 70086 138272
rect 69846 137264 69902 137320
rect 72882 156440 72938 156496
rect 71686 139304 71742 139360
rect 71134 138488 71190 138544
rect 71042 138352 71098 138408
rect 71686 138488 71742 138544
rect 74906 240080 74962 240136
rect 74814 239808 74870 239864
rect 73066 134680 73122 134736
rect 74538 164328 74594 164384
rect 83738 241712 83794 241768
rect 86590 241712 86646 241768
rect 87142 241712 87198 241768
rect 75458 239808 75514 239864
rect 77574 236680 77630 236736
rect 75918 215328 75974 215384
rect 75182 157392 75238 157448
rect 76194 142704 76250 142760
rect 75550 137672 75606 137728
rect 75826 136720 75882 136776
rect 76654 216008 76710 216064
rect 76654 215328 76710 215384
rect 78034 217232 78090 217288
rect 78770 238584 78826 238640
rect 78678 213152 78734 213208
rect 80334 235864 80390 235920
rect 80058 142840 80114 142896
rect 78678 142704 78734 142760
rect 80610 140800 80666 140856
rect 79874 137944 79930 138000
rect 81346 149096 81402 149152
rect 81346 141344 81402 141400
rect 81346 140800 81402 140856
rect 82174 238856 82230 238912
rect 84106 241168 84162 241224
rect 84106 238720 84162 238776
rect 81438 138760 81494 138816
rect 81438 138624 81494 138680
rect 80702 137264 80758 137320
rect 81346 136856 81402 136912
rect 81990 144064 82046 144120
rect 85946 241576 86002 241632
rect 86590 241440 86646 241496
rect 86866 241440 86922 241496
rect 86774 239808 86830 239864
rect 84842 238856 84898 238912
rect 90362 241712 90418 241768
rect 91558 241712 91614 241768
rect 87510 239944 87566 240000
rect 88062 241440 88118 241496
rect 88062 241168 88118 241224
rect 88246 240080 88302 240136
rect 88154 239944 88210 240000
rect 89626 241168 89682 241224
rect 88706 240080 88762 240136
rect 88982 239808 89038 239864
rect 84842 173984 84898 174040
rect 83462 156032 83518 156088
rect 83002 149232 83058 149288
rect 82910 136720 82966 136776
rect 83554 152496 83610 152552
rect 83646 137672 83702 137728
rect 86958 165688 87014 165744
rect 86222 154536 86278 154592
rect 84842 137944 84898 138000
rect 85486 136720 85542 136776
rect 86222 136856 86278 136912
rect 87142 160112 87198 160168
rect 91006 240216 91062 240272
rect 93766 241712 93822 241768
rect 93766 241168 93822 241224
rect 95146 238040 95202 238096
rect 94226 237496 94282 237552
rect 94134 233960 94190 234016
rect 88982 175888 89038 175944
rect 89166 137264 89222 137320
rect 89810 168408 89866 168464
rect 92478 169768 92534 169824
rect 91742 135360 91798 135416
rect 92294 135360 92350 135416
rect 93122 144744 93178 144800
rect 97722 241596 97778 241632
rect 96894 240080 96950 240136
rect 97722 241576 97724 241596
rect 97724 241576 97776 241596
rect 97776 241576 97778 241596
rect 95238 135496 95294 135552
rect 94778 108704 94834 108760
rect 67270 63416 67326 63472
rect 63222 3304 63278 3360
rect 69708 92656 69764 92712
rect 69846 92520 69902 92576
rect 71180 92656 71236 92712
rect 70306 77832 70362 77888
rect 72836 92656 72892 92712
rect 71778 91024 71834 91080
rect 73066 90344 73122 90400
rect 71778 86536 71834 86592
rect 73066 77968 73122 78024
rect 78402 89664 78458 89720
rect 77574 81232 77630 81288
rect 77298 80008 77354 80064
rect 79506 85312 79562 85368
rect 81438 92384 81494 92440
rect 83554 92248 83610 92304
rect 84106 89392 84162 89448
rect 86682 88032 86738 88088
rect 86130 86808 86186 86864
rect 82818 82456 82874 82512
rect 75826 75112 75882 75168
rect 73802 6160 73858 6216
rect 76562 73752 76618 73808
rect 84106 61376 84162 61432
rect 81346 14456 81402 14512
rect 91788 92656 91844 92712
rect 93260 92656 93316 92712
rect 94778 93064 94834 93120
rect 92386 92112 92442 92168
rect 93122 91704 93178 91760
rect 92754 88168 92810 88224
rect 91098 84088 91154 84144
rect 89994 82592 90050 82648
rect 89902 77152 89958 77208
rect 91006 72392 91062 72448
rect 88246 48864 88302 48920
rect 95422 127608 95478 127664
rect 95330 120264 95386 120320
rect 94778 87896 94834 87952
rect 95146 86808 95202 86864
rect 96710 135904 96766 135960
rect 96710 133048 96766 133104
rect 96618 132232 96674 132288
rect 96710 131416 96766 131472
rect 96710 130872 96766 130928
rect 96618 130056 96674 130112
rect 96526 98232 96582 98288
rect 96710 129240 96766 129296
rect 96710 125432 96766 125488
rect 97170 119448 97226 119504
rect 97170 115676 97172 115696
rect 97172 115676 97224 115696
rect 97224 115676 97226 115696
rect 97170 115640 97226 115676
rect 96710 111868 96712 111888
rect 96712 111868 96764 111888
rect 96764 111868 96766 111888
rect 96710 111832 96766 111868
rect 96710 111016 96766 111072
rect 97078 110236 97080 110256
rect 97080 110236 97132 110256
rect 97132 110236 97134 110256
rect 97078 110200 97134 110236
rect 96802 105032 96858 105088
rect 96710 102076 96712 102096
rect 96712 102076 96764 102096
rect 96764 102076 96766 102096
rect 96710 102040 96766 102076
rect 96710 101224 96766 101280
rect 96710 96600 96766 96656
rect 97630 127064 97686 127120
rect 97906 126248 97962 126304
rect 97906 125468 97908 125488
rect 97908 125468 97960 125488
rect 97960 125468 97962 125488
rect 97906 125432 97962 125468
rect 97814 124616 97870 124672
rect 97906 124108 97908 124128
rect 97908 124108 97960 124128
rect 97960 124108 97962 124128
rect 97906 124072 97962 124108
rect 97722 123392 97778 123448
rect 97446 123256 97502 123312
rect 97446 121624 97502 121680
rect 97630 120808 97686 120864
rect 97538 120264 97594 120320
rect 97354 116592 97410 116648
rect 97906 122440 97962 122496
rect 97906 118632 97962 118688
rect 97814 117816 97870 117872
rect 97906 117000 97962 117056
rect 97722 116456 97778 116512
rect 97538 114824 97594 114880
rect 97354 114008 97410 114064
rect 97262 94968 97318 95024
rect 96986 94424 97042 94480
rect 96618 91704 96674 91760
rect 95330 83408 95386 83464
rect 97538 113464 97594 113520
rect 97906 112648 97962 112704
rect 97906 109656 97962 109712
rect 100114 287408 100170 287464
rect 100022 269728 100078 269784
rect 100298 284824 100354 284880
rect 100758 282684 100760 282704
rect 100760 282684 100812 282704
rect 100812 282684 100814 282704
rect 100758 282648 100814 282684
rect 100850 281016 100906 281072
rect 100758 280200 100814 280256
rect 100758 279384 100814 279440
rect 100758 277752 100814 277808
rect 100850 276664 100906 276720
rect 100758 276120 100814 276176
rect 100758 273672 100814 273728
rect 100758 272856 100814 272912
rect 100850 272040 100906 272096
rect 100298 268368 100354 268424
rect 100114 267824 100170 267880
rect 99286 258168 99342 258224
rect 99194 248376 99250 248432
rect 98274 248240 98330 248296
rect 98734 240080 98790 240136
rect 97906 107208 97962 107264
rect 97906 104216 97962 104272
rect 97814 103420 97870 103456
rect 97814 103400 97816 103420
rect 97816 103400 97868 103420
rect 97868 103400 97870 103420
rect 97906 102856 97962 102912
rect 97446 100408 97502 100464
rect 97906 99592 97962 99648
rect 97906 99068 97962 99104
rect 97906 99048 97908 99068
rect 97908 99048 97960 99068
rect 97960 99048 97962 99068
rect 97906 98232 97962 98288
rect 99194 179444 99250 179480
rect 99194 179424 99196 179444
rect 99196 179424 99248 179444
rect 99248 179424 99250 179444
rect 100114 257352 100170 257408
rect 100022 251096 100078 251152
rect 97814 96056 97870 96112
rect 97906 95260 97962 95296
rect 97906 95240 97908 95260
rect 97908 95240 97960 95260
rect 97960 95240 97962 95260
rect 97906 93644 97908 93664
rect 97908 93644 97960 93664
rect 97960 93644 97962 93664
rect 97906 93608 97962 93644
rect 100206 247560 100262 247616
rect 100758 271224 100814 271280
rect 100758 270444 100760 270464
rect 100760 270444 100812 270464
rect 100812 270444 100814 270464
rect 100758 270408 100814 270444
rect 100758 268776 100814 268832
rect 100758 267960 100814 268016
rect 100758 267144 100814 267200
rect 100942 266328 100998 266384
rect 100758 265512 100814 265568
rect 100850 264696 100906 264752
rect 100758 263880 100814 263936
rect 100758 263064 100814 263120
rect 100942 262792 100998 262848
rect 100758 262268 100814 262304
rect 100758 262248 100760 262268
rect 100760 262248 100812 262268
rect 100812 262248 100814 262268
rect 100850 261432 100906 261488
rect 100850 260616 100906 260672
rect 100758 259800 100814 259856
rect 102782 388456 102838 388512
rect 102690 320184 102746 320240
rect 101494 276936 101550 276992
rect 101494 274488 101550 274544
rect 101678 304136 101734 304192
rect 103886 389272 103942 389328
rect 102138 285640 102194 285696
rect 101678 278568 101734 278624
rect 101586 269592 101642 269648
rect 101402 258168 101458 258224
rect 100850 256536 100906 256592
rect 101402 255720 101458 255776
rect 100850 254940 100852 254960
rect 100852 254940 100904 254960
rect 100904 254940 100906 254960
rect 100850 254904 100906 254940
rect 100850 254088 100906 254144
rect 100850 253272 100906 253328
rect 100850 250824 100906 250880
rect 100850 249192 100906 249248
rect 100850 246744 100906 246800
rect 100850 245928 100906 245984
rect 100850 245112 100906 245168
rect 100942 244296 100998 244352
rect 100850 243480 100906 243536
rect 101678 252456 101734 252512
rect 101954 250008 102010 250064
rect 98826 89528 98882 89584
rect 100758 98640 100814 98696
rect 102966 285640 103022 285696
rect 102322 242664 102378 242720
rect 102230 241596 102286 241632
rect 102230 241576 102232 241596
rect 102232 241576 102284 241596
rect 102284 241576 102286 241596
rect 102782 238584 102838 238640
rect 105082 390632 105138 390688
rect 107750 390632 107806 390688
rect 105266 390496 105322 390552
rect 105174 389000 105230 389056
rect 104806 385600 104862 385656
rect 104162 291216 104218 291272
rect 106094 389000 106150 389056
rect 105910 383560 105966 383616
rect 106002 382880 106058 382936
rect 104898 289992 104954 290048
rect 104254 241848 104310 241904
rect 104162 236000 104218 236056
rect 103518 235864 103574 235920
rect 100114 88032 100170 88088
rect 100022 86672 100078 86728
rect 102782 149232 102838 149288
rect 98734 82592 98790 82648
rect 101402 77968 101458 78024
rect 98642 69536 98698 69592
rect 95146 54440 95202 54496
rect 104806 240080 104862 240136
rect 104714 236680 104770 236736
rect 104254 141480 104310 141536
rect 104806 211792 104862 211848
rect 104162 90480 104218 90536
rect 104346 90344 104402 90400
rect 104346 80008 104402 80064
rect 104990 267824 105046 267880
rect 106094 270544 106150 270600
rect 111982 390632 112038 390688
rect 107934 389000 107990 389056
rect 108854 389000 108910 389056
rect 108670 387640 108726 387696
rect 106462 380704 106518 380760
rect 106462 291760 106518 291816
rect 106370 236680 106426 236736
rect 105542 221584 105598 221640
rect 105542 217232 105598 217288
rect 104898 143384 104954 143440
rect 106922 241304 106978 241360
rect 106554 236000 106610 236056
rect 106922 231104 106978 231160
rect 106554 144064 106610 144120
rect 105542 90616 105598 90672
rect 105542 81232 105598 81288
rect 107658 235864 107714 235920
rect 107014 219136 107070 219192
rect 107014 161472 107070 161528
rect 107566 144064 107622 144120
rect 107014 135904 107070 135960
rect 100298 3304 100354 3360
rect 110418 389136 110474 389192
rect 109038 379344 109094 379400
rect 109682 379344 109738 379400
rect 111062 320728 111118 320784
rect 111154 284416 111210 284472
rect 108302 145560 108358 145616
rect 108302 128424 108358 128480
rect 107750 98640 107806 98696
rect 108302 98640 108358 98696
rect 108302 91704 108358 91760
rect 110326 226888 110382 226944
rect 109682 160248 109738 160304
rect 111154 260072 111210 260128
rect 115018 433336 115074 433392
rect 115294 458496 115350 458552
rect 114650 429256 114706 429312
rect 113454 425992 113510 426048
rect 113362 402328 113418 402384
rect 114650 421912 114706 421968
rect 114558 420824 114614 420880
rect 115294 431160 115350 431216
rect 115294 425992 115350 426048
rect 115294 424940 115296 424960
rect 115296 424940 115348 424960
rect 115348 424940 115350 424960
rect 115294 424904 115350 424940
rect 115110 424088 115166 424144
rect 115202 418920 115258 418976
rect 115018 414024 115074 414080
rect 115018 412664 115074 412720
rect 115202 406408 115258 406464
rect 114742 400424 114798 400480
rect 114834 391176 114890 391232
rect 113822 387368 113878 387424
rect 113454 384240 113510 384296
rect 113822 298152 113878 298208
rect 113822 285504 113878 285560
rect 113822 281560 113878 281616
rect 115846 430072 115902 430128
rect 115846 428168 115902 428224
rect 115846 427080 115902 427136
rect 115846 423000 115902 423056
rect 115846 420008 115902 420064
rect 115846 416744 115902 416800
rect 115846 415656 115902 415712
rect 115846 413788 115848 413808
rect 115848 413788 115900 413808
rect 115900 413788 115902 413808
rect 115846 413752 115902 413788
rect 115846 410488 115902 410544
rect 115846 409672 115902 409728
rect 115846 408584 115902 408640
rect 115846 407496 115902 407552
rect 115386 405592 115442 405648
rect 115754 405592 115810 405648
rect 115846 404504 115902 404560
rect 115846 403416 115902 403472
rect 115662 401240 115718 401296
rect 115846 399336 115902 399392
rect 115570 398248 115626 398304
rect 115846 396364 115902 396400
rect 115846 396344 115848 396364
rect 115848 396344 115900 396364
rect 115900 396344 115902 396364
rect 115846 395256 115902 395312
rect 115846 394168 115902 394224
rect 115846 393080 115902 393136
rect 115386 391992 115442 392048
rect 116122 418240 116178 418296
rect 116030 414840 116086 414896
rect 116122 411576 116178 411632
rect 119342 583752 119398 583808
rect 116766 451288 116822 451344
rect 116766 437280 116822 437336
rect 119434 455504 119490 455560
rect 116674 406272 116730 406328
rect 116582 397432 116638 397488
rect 117318 385600 117374 385656
rect 119342 397432 119398 397488
rect 118698 386280 118754 386336
rect 117226 371884 117282 371920
rect 117226 371864 117228 371884
rect 117228 371864 117280 371884
rect 117280 371864 117282 371884
rect 116030 320728 116086 320784
rect 115294 238040 115350 238096
rect 115202 224848 115258 224904
rect 115202 222808 115258 222864
rect 114466 217232 114522 217288
rect 113822 213152 113878 213208
rect 113086 208936 113142 208992
rect 111890 108296 111946 108352
rect 111154 79736 111210 79792
rect 113822 89664 113878 89720
rect 114374 89664 114430 89720
rect 110510 3440 110566 3496
rect 115938 181328 115994 181384
rect 115294 89664 115350 89720
rect 117962 283056 118018 283112
rect 120170 440272 120226 440328
rect 119986 387504 120042 387560
rect 119342 382200 119398 382256
rect 120722 364928 120778 364984
rect 120722 294480 120778 294536
rect 120170 289040 120226 289096
rect 119342 233960 119398 234016
rect 119986 225664 120042 225720
rect 119342 88168 119398 88224
rect 123482 462848 123538 462904
rect 122102 366968 122158 367024
rect 122746 310664 122802 310720
rect 121550 104080 121606 104136
rect 122930 304136 122986 304192
rect 122838 301416 122894 301472
rect 122838 143248 122894 143304
rect 122838 142704 122894 142760
rect 124310 380704 124366 380760
rect 124862 417424 124918 417480
rect 124862 400832 124918 400888
rect 124862 380704 124918 380760
rect 124402 379344 124458 379400
rect 125782 406272 125838 406328
rect 133142 582664 133198 582720
rect 128450 417424 128506 417480
rect 126886 386280 126942 386336
rect 127622 380840 127678 380896
rect 126334 370504 126390 370560
rect 126242 298696 126298 298752
rect 124954 153176 125010 153232
rect 133142 460944 133198 461000
rect 132498 434696 132554 434752
rect 129094 384920 129150 384976
rect 126334 233960 126390 234016
rect 129094 320184 129150 320240
rect 129094 287680 129150 287736
rect 129094 287136 129150 287192
rect 129002 276664 129058 276720
rect 126334 147736 126390 147792
rect 129186 270544 129242 270600
rect 131762 302368 131818 302424
rect 133142 300872 133198 300928
rect 136638 536016 136694 536072
rect 136546 387640 136602 387696
rect 142066 451832 142122 451888
rect 135902 328480 135958 328536
rect 134614 291760 134670 291816
rect 137466 326304 137522 326360
rect 137374 267144 137430 267200
rect 137282 261432 137338 261488
rect 137466 251096 137522 251152
rect 140042 268504 140098 268560
rect 141514 287680 141570 287736
rect 141514 273808 141570 273864
rect 147586 454144 147642 454200
rect 144182 380840 144238 380896
rect 146942 331200 146998 331256
rect 144182 316104 144238 316160
rect 142986 269728 143042 269784
rect 145562 317464 145618 317520
rect 144182 156168 144238 156224
rect 147034 164328 147090 164384
rect 155222 376488 155278 376544
rect 148414 301416 148470 301472
rect 149886 274760 149942 274816
rect 149794 153312 149850 153368
rect 152462 303864 152518 303920
rect 151174 280744 151230 280800
rect 151266 157528 151322 157584
rect 155406 327120 155462 327176
rect 152554 271088 152610 271144
rect 152554 154672 152610 154728
rect 152646 135904 152702 135960
rect 153106 94696 153162 94752
rect 153934 233960 153990 234016
rect 155314 293120 155370 293176
rect 156602 289040 156658 289096
rect 155958 267008 156014 267064
rect 156418 267028 156474 267064
rect 156418 267008 156420 267028
rect 156420 267008 156472 267028
rect 156472 267008 156474 267028
rect 155314 149368 155370 149424
rect 157246 287000 157302 287056
rect 157246 285776 157302 285832
rect 166262 453056 166318 453112
rect 158718 376624 158774 376680
rect 159454 376624 159510 376680
rect 159362 332560 159418 332616
rect 159546 321544 159602 321600
rect 158626 269728 158682 269784
rect 158074 235320 158130 235376
rect 156694 151136 156750 151192
rect 155958 144744 156014 144800
rect 156694 144744 156750 144800
rect 156694 143520 156750 143576
rect 157982 138624 158038 138680
rect 160926 285796 160982 285832
rect 160926 285776 160928 285796
rect 160928 285776 160980 285796
rect 160980 285776 160982 285796
rect 159546 268368 159602 268424
rect 159454 217912 159510 217968
rect 155314 93064 155370 93120
rect 155498 93064 155554 93120
rect 157982 82592 158038 82648
rect 159546 145696 159602 145752
rect 161938 322088 161994 322144
rect 166262 406272 166318 406328
rect 163502 318824 163558 318880
rect 162122 313384 162178 313440
rect 162766 313384 162822 313440
rect 161386 282784 161442 282840
rect 161110 272448 161166 272504
rect 162306 282784 162362 282840
rect 162306 281560 162362 281616
rect 162122 265104 162178 265160
rect 162214 106256 162270 106312
rect 163686 262792 163742 262848
rect 166354 388864 166410 388920
rect 166262 377304 166318 377360
rect 166446 290400 166502 290456
rect 166446 289856 166502 289912
rect 167642 322904 167698 322960
rect 169666 442992 169722 443048
rect 168378 381656 168434 381712
rect 169022 375264 169078 375320
rect 168286 322904 168342 322960
rect 166538 238040 166594 238096
rect 166538 237360 166594 237416
rect 166906 237360 166962 237416
rect 170494 364928 170550 364984
rect 168470 281560 168526 281616
rect 168286 152496 168342 152552
rect 167642 75112 167698 75168
rect 169114 179968 169170 180024
rect 169758 289040 169814 289096
rect 170678 314880 170734 314936
rect 170954 314880 171010 314936
rect 170770 260072 170826 260128
rect 175186 457000 175242 457056
rect 173254 384920 173310 384976
rect 173806 384920 173862 384976
rect 173254 368328 173310 368384
rect 172610 269728 172666 269784
rect 172610 235592 172666 235648
rect 172518 135224 172574 135280
rect 173254 240896 173310 240952
rect 174726 329840 174782 329896
rect 173254 220224 173310 220280
rect 173346 144200 173402 144256
rect 173806 135224 173862 135280
rect 173346 123392 173402 123448
rect 173254 95240 173310 95296
rect 176014 304952 176070 305008
rect 176566 304952 176622 305008
rect 175186 236680 175242 236736
rect 175186 209616 175242 209672
rect 176750 396616 176806 396672
rect 184202 463664 184258 463720
rect 180062 461080 180118 461136
rect 178682 454008 178738 454064
rect 177302 309304 177358 309360
rect 176658 293936 176714 293992
rect 177210 293936 177266 293992
rect 183466 456864 183522 456920
rect 180154 455776 180210 455832
rect 178682 291896 178738 291952
rect 177946 240080 178002 240136
rect 177946 235864 178002 235920
rect 177394 144880 177450 144936
rect 177946 92384 178002 92440
rect 178866 284280 178922 284336
rect 178866 239672 178922 239728
rect 179510 388456 179566 388512
rect 179510 387776 179566 387832
rect 179326 228928 179382 228984
rect 181534 447888 181590 447944
rect 180154 369688 180210 369744
rect 182086 317328 182142 317384
rect 182086 316648 182142 316704
rect 181534 300056 181590 300112
rect 181534 291760 181590 291816
rect 181442 285504 181498 285560
rect 180246 273808 180302 273864
rect 180062 228248 180118 228304
rect 180062 226208 180118 226264
rect 181442 264968 181498 265024
rect 180246 230424 180302 230480
rect 180614 226208 180670 226264
rect 180154 217232 180210 217288
rect 180062 215872 180118 215928
rect 178774 83952 178830 84008
rect 179418 92248 179474 92304
rect 180062 86672 180118 86728
rect 181534 246200 181590 246256
rect 182086 238584 182142 238640
rect 181534 231784 181590 231840
rect 181534 210296 181590 210352
rect 181534 143520 181590 143576
rect 182362 119992 182418 120048
rect 183466 318688 183522 318744
rect 183466 318008 183522 318064
rect 183466 291896 183522 291952
rect 184202 317328 184258 317384
rect 184202 308080 184258 308136
rect 185674 458360 185730 458416
rect 184938 320048 184994 320104
rect 184846 290400 184902 290456
rect 184202 280744 184258 280800
rect 182914 251776 182970 251832
rect 187054 450064 187110 450120
rect 187054 437416 187110 437472
rect 186962 431976 187018 432032
rect 186962 418240 187018 418296
rect 187054 400832 187110 400888
rect 187054 386144 187110 386200
rect 185674 320048 185730 320104
rect 185674 309440 185730 309496
rect 184294 236816 184350 236872
rect 184294 232600 184350 232656
rect 184478 234504 184534 234560
rect 184294 228928 184350 228984
rect 184294 227704 184350 227760
rect 183006 214512 183062 214568
rect 183006 147056 183062 147112
rect 183006 133864 183062 133920
rect 183006 119992 183062 120048
rect 182914 85312 182970 85368
rect 182822 77832 182878 77888
rect 184386 150456 184442 150512
rect 188066 452920 188122 452976
rect 188066 444896 188122 444952
rect 188802 432520 188858 432576
rect 188526 382336 188582 382392
rect 188526 373904 188582 373960
rect 189722 452784 189778 452840
rect 189722 438776 189778 438832
rect 190274 412664 190330 412720
rect 190182 394712 190238 394768
rect 190090 393352 190146 393408
rect 190090 382880 190146 382936
rect 190090 382336 190146 382392
rect 189078 381520 189134 381576
rect 187698 361528 187754 361584
rect 188618 318960 188674 319016
rect 188618 312432 188674 312488
rect 188434 312024 188490 312080
rect 187698 305088 187754 305144
rect 187698 298832 187754 298888
rect 185766 151136 185822 151192
rect 185674 148280 185730 148336
rect 185582 145016 185638 145072
rect 184294 81368 184350 81424
rect 184386 79872 184442 79928
rect 185766 122848 185822 122904
rect 188342 282920 188398 282976
rect 187606 265512 187662 265568
rect 187054 264968 187110 265024
rect 187054 241440 187110 241496
rect 187606 241440 187662 241496
rect 187698 240896 187754 240952
rect 187606 240760 187662 240816
rect 187146 233824 187202 233880
rect 186962 144064 187018 144120
rect 186870 135904 186926 135960
rect 185582 89528 185638 89584
rect 189078 367104 189134 367160
rect 188986 361528 189042 361584
rect 188342 239808 188398 239864
rect 188526 248376 188582 248432
rect 188434 237904 188490 237960
rect 190182 367104 190238 367160
rect 190458 447208 190514 447264
rect 191286 454280 191342 454336
rect 191194 446392 191250 446448
rect 191470 449112 191526 449168
rect 191654 449112 191710 449168
rect 208398 470600 208454 470656
rect 194598 465160 194654 465216
rect 191746 446392 191802 446448
rect 191746 445032 191802 445088
rect 191746 437960 191802 438016
rect 191746 435240 191802 435296
rect 191654 433608 191710 433664
rect 191194 429528 191250 429584
rect 191470 429528 191526 429584
rect 191010 425448 191066 425504
rect 190826 422456 190882 422512
rect 191010 415384 191066 415440
rect 191562 428168 191618 428224
rect 191562 426808 191618 426864
rect 191562 419736 191618 419792
rect 191562 418376 191618 418432
rect 191562 417016 191618 417072
rect 191562 414024 191618 414080
rect 191470 411304 191526 411360
rect 190826 409944 190882 410000
rect 191470 406952 191526 407008
rect 191378 405592 191434 405648
rect 191470 404232 191526 404288
rect 191378 402872 191434 402928
rect 190826 400152 190882 400208
rect 191102 398520 191158 398576
rect 191470 401512 191526 401568
rect 191470 397160 191526 397216
rect 191010 390904 191066 390960
rect 189722 272448 189778 272504
rect 189722 245792 189778 245848
rect 188986 241032 189042 241088
rect 188986 240080 189042 240136
rect 188526 235184 188582 235240
rect 187698 216008 187754 216064
rect 187698 215328 187754 215384
rect 188342 215328 188398 215384
rect 188894 201320 188950 201376
rect 189998 306448 190054 306504
rect 191102 301552 191158 301608
rect 191102 301028 191158 301064
rect 191102 301008 191104 301028
rect 191104 301008 191156 301028
rect 191156 301008 191158 301028
rect 190642 298968 190698 299024
rect 189998 294480 190054 294536
rect 190642 287408 190698 287464
rect 191010 286456 191066 286512
rect 191102 284280 191158 284336
rect 189814 232464 189870 232520
rect 189998 242936 190054 242992
rect 189998 236544 190054 236600
rect 189906 224712 189962 224768
rect 189722 162832 189778 162888
rect 188894 158752 188950 158808
rect 187698 147872 187754 147928
rect 188434 146376 188490 146432
rect 187698 145560 187754 145616
rect 189078 142160 189134 142216
rect 188894 128424 188950 128480
rect 187606 87896 187662 87952
rect 188342 85448 188398 85504
rect 187054 81096 187110 81152
rect 187698 71732 187754 71768
rect 187698 71712 187700 71732
rect 187700 71712 187752 71732
rect 187752 71712 187754 71732
rect 188526 93064 188582 93120
rect 189078 139304 189134 139360
rect 189814 135088 189870 135144
rect 189722 132504 189778 132560
rect 189722 124208 189778 124264
rect 188894 71712 188950 71768
rect 190826 270000 190882 270056
rect 190826 266056 190882 266112
rect 191010 263200 191066 263256
rect 190826 256400 190882 256456
rect 191010 255448 191066 255504
rect 190642 250688 190698 250744
rect 190826 249600 190882 249656
rect 190366 138488 190422 138544
rect 189906 133864 189962 133920
rect 191470 391720 191526 391776
rect 191470 298016 191526 298072
rect 191562 291216 191618 291272
rect 191562 289312 191618 289368
rect 193310 451424 193366 451480
rect 194598 450200 194654 450256
rect 197082 458260 197084 458280
rect 197084 458260 197136 458280
rect 197136 458260 197138 458280
rect 197082 458224 197138 458260
rect 197910 454144 197966 454200
rect 207478 457000 207534 457056
rect 202878 455640 202934 455696
rect 202142 452920 202198 452976
rect 201590 450336 201646 450392
rect 204442 451832 204498 451888
rect 207018 451424 207074 451480
rect 210698 452784 210754 452840
rect 210698 451424 210754 451480
rect 213918 465160 213974 465216
rect 215206 465160 215262 465216
rect 212538 462168 212594 462224
rect 213182 462168 213238 462224
rect 212538 461080 212594 461136
rect 215298 465024 215354 465080
rect 215942 465024 215998 465080
rect 215298 463664 215354 463720
rect 215390 456864 215446 456920
rect 216678 458632 216734 458688
rect 216678 458360 216734 458416
rect 220082 458632 220138 458688
rect 220818 458360 220874 458416
rect 219806 455776 219862 455832
rect 222566 454280 222622 454336
rect 222106 452920 222162 452976
rect 224958 455640 225014 455696
rect 225970 453056 226026 453112
rect 225602 452784 225658 452840
rect 230478 456864 230534 456920
rect 231122 456864 231178 456920
rect 228730 452784 228786 452840
rect 228086 450200 228142 450256
rect 220818 449928 220874 449984
rect 235354 451560 235410 451616
rect 233146 450064 233202 450120
rect 242162 455368 242218 455424
rect 243542 455368 243598 455424
rect 243542 454144 243598 454200
rect 246026 452920 246082 452976
rect 242438 450064 242494 450120
rect 237654 449928 237710 449984
rect 251546 452920 251602 452976
rect 249706 451288 249762 451344
rect 250258 449928 250314 449984
rect 193494 449656 193550 449712
rect 242990 449656 243046 449712
rect 252466 452648 252522 452704
rect 253846 452784 253902 452840
rect 193310 447888 193366 447944
rect 193126 442040 193182 442096
rect 192942 436600 192998 436656
rect 191838 425448 191894 425504
rect 192850 423816 192906 423872
rect 193034 408584 193090 408640
rect 192942 386960 192998 387016
rect 192850 385600 192906 385656
rect 254122 459584 254178 459640
rect 253938 440408 253994 440464
rect 253938 431976 253994 432032
rect 193310 391176 193366 391232
rect 253662 392808 253718 392864
rect 195978 390768 196034 390824
rect 193126 363568 193182 363624
rect 197358 383832 197414 383888
rect 197358 381656 197414 381712
rect 195978 355952 196034 356008
rect 196622 355952 196678 356008
rect 196622 355272 196678 355328
rect 193494 353912 193550 353968
rect 192574 306584 192630 306640
rect 191746 300872 191802 300928
rect 191746 299940 191802 299976
rect 191746 299920 191748 299940
rect 191748 299920 191800 299940
rect 191800 299920 191802 299940
rect 192206 299512 192262 299568
rect 192758 302268 192760 302288
rect 192760 302268 192812 302288
rect 192812 302268 192814 302288
rect 192758 302232 192814 302268
rect 192574 298152 192630 298208
rect 191746 297064 191802 297120
rect 192482 295160 192538 295216
rect 191746 294208 191802 294264
rect 191746 292596 191802 292632
rect 191746 292576 191748 292596
rect 191748 292576 191800 292596
rect 191800 292576 191802 292596
rect 191746 292168 191802 292224
rect 191746 290300 191748 290320
rect 191748 290300 191800 290320
rect 191800 290300 191802 290320
rect 191746 290264 191802 290300
rect 191746 288380 191802 288416
rect 191746 288360 191748 288380
rect 191748 288360 191800 288380
rect 191800 288360 191802 288380
rect 191654 285504 191710 285560
rect 191746 284416 191802 284472
rect 191654 284280 191710 284336
rect 191562 282512 191618 282568
rect 191746 281580 191802 281616
rect 191746 281560 191748 281580
rect 191748 281560 191800 281580
rect 191800 281560 191802 281580
rect 191286 280608 191342 280664
rect 191562 279656 191618 279712
rect 191194 274760 191250 274816
rect 191562 274760 191618 274816
rect 191470 269048 191526 269104
rect 191654 272856 191710 272912
rect 191746 271940 191748 271960
rect 191748 271940 191800 271960
rect 191800 271940 191802 271960
rect 191746 271904 191802 271940
rect 191746 270952 191802 271008
rect 191746 268096 191802 268152
rect 191562 261296 191618 261352
rect 191746 267008 191802 267064
rect 191746 264152 191802 264208
rect 191746 262268 191802 262304
rect 191746 262248 191748 262268
rect 191748 262248 191800 262268
rect 191800 262248 191802 262268
rect 191746 260344 191802 260400
rect 191746 258304 191802 258360
rect 191654 257352 191710 257408
rect 191654 254496 191710 254552
rect 191562 253544 191618 253600
rect 191654 252628 191656 252648
rect 191656 252628 191708 252648
rect 191708 252628 191710 252648
rect 191654 252592 191710 252628
rect 191654 247696 191710 247752
rect 191654 244840 191710 244896
rect 191654 243888 191710 243944
rect 191654 139848 191710 139904
rect 191654 136312 191710 136368
rect 191654 135496 191710 135552
rect 191194 131960 191250 132016
rect 190826 130056 190882 130112
rect 191010 125740 191012 125760
rect 191012 125740 191064 125760
rect 191064 125740 191066 125760
rect 191010 125704 191066 125740
rect 191654 129240 191710 129296
rect 191654 127608 191710 127664
rect 191562 122168 191618 122224
rect 190826 121352 190882 121408
rect 190274 110744 190330 110800
rect 189906 98232 189962 98288
rect 189814 92248 189870 92304
rect 190458 120264 190514 120320
rect 191562 119448 191618 119504
rect 191562 118632 191618 118688
rect 190826 117972 190882 118008
rect 190826 117952 190828 117972
rect 190828 117952 190880 117972
rect 190880 117952 190882 117972
rect 191562 116728 191618 116784
rect 191378 115912 191434 115968
rect 191010 115096 191066 115152
rect 190826 114008 190882 114064
rect 191562 113192 191618 113248
rect 191562 112376 191618 112432
rect 191194 110472 191250 110528
rect 191010 109656 191066 109712
rect 190642 106936 190698 106992
rect 191010 106120 191066 106176
rect 191562 105032 191618 105088
rect 191562 103400 191618 103456
rect 191470 102584 191526 102640
rect 190642 101496 190698 101552
rect 190642 97144 190698 97200
rect 191562 100680 191618 100736
rect 191102 84224 191158 84280
rect 191470 84224 191526 84280
rect 192942 302232 192998 302288
rect 193034 296112 193090 296168
rect 193310 295160 193366 295216
rect 193034 283464 193090 283520
rect 192942 280608 192998 280664
rect 192850 277752 192906 277808
rect 192022 246200 192078 246256
rect 192022 245656 192078 245712
rect 192482 237904 192538 237960
rect 195702 303728 195758 303784
rect 194138 301552 194194 301608
rect 198094 367104 198150 367160
rect 201130 388320 201186 388376
rect 200118 356632 200174 356688
rect 197450 312024 197506 312080
rect 198738 323060 198794 323096
rect 198738 323040 198740 323060
rect 198740 323040 198792 323060
rect 198792 323040 198794 323060
rect 204258 376624 204314 376680
rect 205546 376624 205602 376680
rect 202326 324400 202382 324456
rect 200302 316104 200358 316160
rect 200210 309168 200266 309224
rect 199474 306448 199530 306504
rect 198094 303456 198150 303512
rect 200118 302504 200174 302560
rect 202050 307808 202106 307864
rect 201406 303456 201462 303512
rect 203430 311888 203486 311944
rect 207754 384920 207810 384976
rect 205546 313928 205602 313984
rect 207018 317464 207074 317520
rect 205638 310528 205694 310584
rect 208490 385600 208546 385656
rect 208490 367648 208546 367704
rect 213458 388456 213514 388512
rect 212538 371864 212594 371920
rect 208398 337320 208454 337376
rect 216402 383968 216458 384024
rect 213918 334600 213974 334656
rect 211802 331744 211858 331800
rect 208398 328480 208454 328536
rect 207110 307672 207166 307728
rect 207110 306992 207166 307048
rect 207662 302368 207718 302424
rect 210238 306584 210294 306640
rect 209594 305224 209650 305280
rect 219438 361528 219494 361584
rect 215942 325760 215998 325816
rect 216218 318008 216274 318064
rect 211802 312432 211858 312488
rect 212722 308080 212778 308136
rect 214010 305088 214066 305144
rect 213366 303864 213422 303920
rect 216218 311208 216274 311264
rect 219990 310664 220046 310720
rect 218058 308352 218114 308408
rect 218058 303592 218114 303648
rect 220818 313248 220874 313304
rect 223486 326304 223542 326360
rect 223118 314744 223174 314800
rect 222198 307672 222254 307728
rect 221554 306720 221610 306776
rect 222566 301552 222622 301608
rect 228362 338680 228418 338736
rect 227810 331200 227866 331256
rect 227718 305088 227774 305144
rect 225050 301824 225106 301880
rect 226982 301552 227038 301608
rect 234066 389408 234122 389464
rect 231122 355408 231178 355464
rect 233882 384240 233938 384296
rect 232594 357992 232650 358048
rect 236274 386416 236330 386472
rect 238114 384376 238170 384432
rect 237378 370504 237434 370560
rect 232502 316648 232558 316704
rect 237378 369824 237434 369880
rect 238022 369824 238078 369880
rect 235262 314064 235318 314120
rect 240138 389272 240194 389328
rect 241058 389272 241114 389328
rect 238114 307128 238170 307184
rect 233882 305632 233938 305688
rect 229190 303728 229246 303784
rect 229834 302232 229890 302288
rect 236090 302232 236146 302288
rect 231306 301552 231362 301608
rect 235262 301552 235318 301608
rect 237746 301552 237802 301608
rect 240874 303592 240930 303648
rect 241150 302232 241206 302288
rect 240230 301688 240286 301744
rect 241058 301688 241114 301744
rect 242990 383560 243046 383616
rect 244002 383560 244058 383616
rect 244370 380160 244426 380216
rect 244278 353912 244334 353968
rect 242806 304136 242862 304192
rect 203062 301416 203118 301472
rect 204350 301416 204406 301472
rect 207018 301416 207074 301472
rect 210606 301416 210662 301472
rect 216770 301416 216826 301472
rect 222566 301416 222622 301472
rect 223854 301416 223910 301472
rect 225786 301416 225842 301472
rect 226706 301416 226762 301472
rect 228270 301416 228326 301472
rect 230110 301416 230166 301472
rect 230570 301416 230626 301472
rect 232134 301416 232190 301472
rect 232686 301416 232742 301472
rect 233330 301416 233386 301472
rect 233974 301416 234030 301472
rect 234802 301416 234858 301472
rect 236642 301416 236698 301472
rect 237654 301416 237710 301472
rect 239678 301416 239734 301472
rect 244370 329840 244426 329896
rect 244462 314880 244518 314936
rect 247038 388320 247094 388376
rect 247682 388320 247738 388376
rect 247038 387640 247094 387696
rect 245750 363568 245806 363624
rect 244554 308352 244610 308408
rect 245566 303592 245622 303648
rect 249706 390224 249762 390280
rect 248694 379344 248750 379400
rect 249062 379344 249118 379400
rect 249982 389136 250038 389192
rect 249982 377984 250038 378040
rect 249062 316648 249118 316704
rect 246302 308488 246358 308544
rect 245842 306448 245898 306504
rect 245750 301688 245806 301744
rect 246486 301552 246542 301608
rect 248786 302368 248842 302424
rect 243450 301416 243506 301472
rect 246578 301416 246634 301472
rect 247866 301416 247922 301472
rect 249706 336640 249762 336696
rect 249614 321680 249670 321736
rect 249338 307672 249394 307728
rect 249338 306448 249394 306504
rect 249706 307672 249762 307728
rect 251914 389136 251970 389192
rect 251270 360848 251326 360904
rect 252558 368364 252560 368384
rect 252560 368364 252612 368384
rect 252612 368364 252614 368384
rect 252558 368328 252614 368364
rect 255318 455504 255374 455560
rect 254674 451288 254730 451344
rect 254122 447480 254178 447536
rect 254582 447480 254638 447536
rect 255318 444760 255374 444816
rect 255134 442040 255190 442096
rect 255226 436736 255282 436792
rect 255226 424224 255282 424280
rect 254122 413752 254178 413808
rect 254030 391448 254086 391504
rect 253938 364928 253994 364984
rect 254214 402600 254270 402656
rect 250718 313384 250774 313440
rect 249614 302368 249670 302424
rect 252558 338000 252614 338056
rect 251914 308352 251970 308408
rect 251270 307128 251326 307184
rect 251914 303864 251970 303920
rect 251270 303592 251326 303648
rect 250718 302776 250774 302832
rect 252558 321680 252614 321736
rect 250258 301416 250314 301472
rect 252834 300192 252890 300248
rect 193586 298696 193642 298752
rect 252834 296928 252890 296984
rect 252834 296520 252890 296576
rect 193126 278704 193182 278760
rect 193402 278704 193458 278760
rect 193034 232464 193090 232520
rect 193218 276800 193274 276856
rect 193402 258848 193458 258904
rect 193678 242800 193734 242856
rect 193126 210296 193182 210352
rect 192482 153040 192538 153096
rect 192574 144880 192630 144936
rect 193218 178608 193274 178664
rect 192666 138216 192722 138272
rect 192942 138216 192998 138272
rect 192482 137264 192538 137320
rect 192482 134680 192538 134736
rect 191746 100816 191802 100872
rect 191746 99864 191802 99920
rect 191746 97996 191748 98016
rect 191748 97996 191800 98016
rect 191800 97996 191802 98016
rect 191746 97960 191802 97996
rect 192574 132096 192630 132152
rect 193126 126520 193182 126576
rect 193034 123800 193090 123856
rect 193034 96328 193090 96384
rect 192574 86128 192630 86184
rect 193034 78376 193090 78432
rect 193402 145696 193458 145752
rect 194598 140528 194654 140584
rect 201590 241440 201646 241496
rect 198002 239944 198058 240000
rect 195242 214648 195298 214704
rect 196622 235728 196678 235784
rect 195978 163376 196034 163432
rect 197358 181328 197414 181384
rect 196622 142160 196678 142216
rect 208398 241440 208454 241496
rect 204258 240080 204314 240136
rect 204258 239400 204314 239456
rect 202234 236816 202290 236872
rect 198646 228384 198702 228440
rect 198094 214512 198150 214568
rect 198094 161608 198150 161664
rect 198738 228248 198794 228304
rect 198646 143112 198702 143168
rect 202234 235728 202290 235784
rect 202786 235728 202842 235784
rect 200854 211928 200910 211984
rect 199382 161608 199438 161664
rect 200210 164192 200266 164248
rect 200854 164192 200910 164248
rect 200302 157392 200358 157448
rect 203522 184184 203578 184240
rect 200302 153040 200358 153096
rect 201590 152496 201646 152552
rect 202050 152360 202106 152416
rect 206374 229064 206430 229120
rect 203522 159296 203578 159352
rect 202142 144200 202198 144256
rect 204258 151000 204314 151056
rect 207662 206216 207718 206272
rect 207018 175208 207074 175264
rect 207662 175208 207718 175264
rect 207018 173984 207074 174040
rect 204994 142160 205050 142216
rect 206282 143384 206338 143440
rect 206834 143384 206890 143440
rect 206466 143248 206522 143304
rect 209778 240080 209834 240136
rect 215206 241476 215208 241496
rect 215208 241476 215260 241496
rect 215260 241476 215262 241496
rect 208122 144064 208178 144120
rect 208122 141344 208178 141400
rect 211158 221584 211214 221640
rect 211158 219272 211214 219328
rect 212446 219272 212502 219328
rect 209134 156032 209190 156088
rect 209226 154536 209282 154592
rect 213182 219136 213238 219192
rect 213182 218048 213238 218104
rect 212630 175888 212686 175944
rect 213182 175888 213238 175944
rect 211802 155896 211858 155952
rect 212446 155896 212502 155952
rect 211802 154536 211858 154592
rect 209226 151680 209282 151736
rect 209042 143792 209098 143848
rect 210054 146920 210110 146976
rect 209962 140936 210018 140992
rect 211158 149096 211214 149152
rect 211250 143656 211306 143712
rect 212446 149096 212502 149152
rect 213918 172488 213974 172544
rect 212630 143384 212686 143440
rect 213274 151000 213330 151056
rect 213458 143384 213514 143440
rect 215206 241440 215262 241476
rect 218610 241440 218666 241496
rect 218702 239672 218758 239728
rect 220910 241440 220966 241496
rect 221554 241440 221610 241496
rect 220082 228928 220138 228984
rect 220082 227704 220138 227760
rect 219714 177384 219770 177440
rect 215298 165688 215354 165744
rect 215390 160112 215446 160168
rect 218702 152632 218758 152688
rect 217230 145016 217286 145072
rect 222290 230288 222346 230344
rect 222106 222964 222162 223000
rect 222106 222944 222108 222964
rect 222108 222944 222160 222964
rect 222160 222944 222162 222964
rect 222290 221448 222346 221504
rect 223762 217232 223818 217288
rect 222198 169768 222254 169824
rect 222842 169768 222898 169824
rect 220818 168408 220874 168464
rect 219438 142160 219494 142216
rect 221922 142160 221978 142216
rect 225510 241440 225566 241496
rect 229098 240080 229154 240136
rect 228546 239400 228602 239456
rect 228454 236544 228510 236600
rect 223394 143520 223450 143576
rect 214286 140800 214342 140856
rect 196806 140392 196862 140448
rect 224222 157528 224278 157584
rect 224222 142296 224278 142352
rect 223394 140392 223450 140448
rect 193218 104216 193274 104272
rect 211710 93336 211766 93392
rect 224774 93336 224830 93392
rect 193310 75792 193366 75848
rect 193862 75792 193918 75848
rect 196162 92656 196218 92712
rect 196530 92384 196586 92440
rect 197358 92520 197414 92576
rect 197082 86536 197138 86592
rect 194598 66136 194654 66192
rect 195242 66136 195298 66192
rect 198738 92520 198794 92576
rect 199474 92520 199530 92576
rect 199290 92384 199346 92440
rect 197450 78512 197506 78568
rect 200762 86672 200818 86728
rect 201590 92792 201646 92848
rect 202602 92248 202658 92304
rect 203522 90480 203578 90536
rect 201866 90208 201922 90264
rect 202786 90208 202842 90264
rect 200394 85312 200450 85368
rect 201314 85312 201370 85368
rect 204442 90616 204498 90672
rect 203706 90344 203762 90400
rect 204350 90208 204406 90264
rect 204166 80008 204222 80064
rect 205454 92792 205510 92848
rect 205546 90208 205602 90264
rect 206098 89528 206154 89584
rect 204994 88032 205050 88088
rect 204442 86808 204498 86864
rect 204350 79736 204406 79792
rect 203522 79600 203578 79656
rect 204166 79600 204222 79656
rect 204350 79464 204406 79520
rect 204902 79464 204958 79520
rect 208398 92792 208454 92848
rect 208674 90208 208730 90264
rect 209686 90208 209742 90264
rect 209226 89664 209282 89720
rect 210054 92792 210110 92848
rect 212170 91840 212226 91896
rect 209778 82728 209834 82784
rect 214562 91704 214618 91760
rect 214562 89392 214618 89448
rect 214838 89664 214894 89720
rect 216034 92656 216090 92712
rect 215850 90888 215906 90944
rect 219530 89936 219586 89992
rect 220266 92792 220322 92848
rect 219714 90888 219770 90944
rect 213274 79872 213330 79928
rect 219438 84088 219494 84144
rect 220082 89936 220138 89992
rect 220726 90888 220782 90944
rect 220634 89528 220690 89584
rect 222658 92928 222714 92984
rect 221922 88168 221978 88224
rect 220082 77152 220138 77208
rect 223946 92792 224002 92848
rect 225050 129512 225106 129568
rect 225050 104896 225106 104952
rect 224314 90888 224370 90944
rect 226338 147056 226394 147112
rect 226338 139848 226394 139904
rect 226338 131960 226394 132016
rect 225602 130872 225658 130928
rect 226338 130056 226394 130112
rect 225326 129240 225382 129296
rect 225234 116728 225290 116784
rect 225142 100680 225198 100736
rect 226614 138216 226670 138272
rect 226614 137128 226670 137184
rect 226614 133592 226670 133648
rect 226522 132776 226578 132832
rect 226522 126520 226578 126576
rect 226614 125704 226670 125760
rect 226614 122984 226670 123040
rect 226614 122168 226670 122224
rect 226614 120264 226670 120320
rect 226614 119448 226670 119504
rect 226614 117544 226670 117600
rect 226614 115948 226616 115968
rect 226616 115948 226668 115968
rect 226668 115948 226670 115968
rect 226614 115912 226670 115948
rect 226522 113192 226578 113248
rect 226798 140392 226854 140448
rect 226798 134680 226854 134736
rect 227074 128424 227130 128480
rect 226798 127336 226854 127392
rect 226798 124616 226854 124672
rect 226798 118360 226854 118416
rect 226614 112104 226670 112160
rect 226706 110472 226762 110528
rect 226430 109656 226486 109712
rect 226614 108568 226670 108624
rect 226706 106936 226762 106992
rect 226706 105848 226762 105904
rect 226522 104216 226578 104272
rect 226614 103400 226670 103456
rect 226430 99592 226486 99648
rect 226430 98776 226486 98832
rect 226338 95240 226394 95296
rect 226706 97996 226708 98016
rect 226708 97996 226760 98016
rect 226760 97996 226762 98016
rect 226706 97960 226762 97996
rect 226522 97144 226578 97200
rect 226982 111288 227038 111344
rect 227442 101496 227498 101552
rect 226982 96056 227038 96112
rect 226798 94424 226854 94480
rect 226890 93608 226946 93664
rect 226522 92384 226578 92440
rect 226430 89392 226486 89448
rect 227994 114824 228050 114880
rect 227810 114008 227866 114064
rect 227902 102312 227958 102368
rect 227718 89936 227774 89992
rect 227718 88984 227774 89040
rect 234618 240080 234674 240136
rect 233882 238720 233938 238776
rect 231766 235184 231822 235240
rect 229834 233960 229890 234016
rect 229834 233144 229890 233200
rect 229098 208936 229154 208992
rect 229098 153176 229154 153232
rect 229190 147872 229246 147928
rect 231858 160248 231914 160304
rect 230478 150456 230534 150512
rect 229834 147872 229890 147928
rect 229834 142160 229890 142216
rect 227994 81368 228050 81424
rect 231950 143656 232006 143712
rect 230478 83952 230534 84008
rect 235446 241440 235502 241496
rect 238666 241440 238722 241496
rect 238758 241032 238814 241088
rect 238758 235864 238814 235920
rect 237378 227060 237380 227080
rect 237380 227060 237432 227080
rect 237432 227060 237434 227080
rect 237378 227024 237434 227060
rect 237378 222844 237380 222864
rect 237380 222844 237432 222864
rect 237432 222844 237434 222864
rect 237378 222808 237434 222844
rect 238666 222808 238722 222864
rect 236090 161472 236146 161528
rect 237378 154400 237434 154456
rect 236642 140936 236698 140992
rect 236090 138488 236146 138544
rect 234618 72392 234674 72448
rect 238022 154672 238078 154728
rect 237562 154400 237618 154456
rect 237562 153312 237618 153368
rect 240046 228404 240102 228440
rect 240046 228384 240048 228404
rect 240048 228384 240100 228404
rect 240100 228384 240102 228404
rect 240230 224848 240286 224904
rect 238850 164328 238906 164384
rect 238758 152360 238814 152416
rect 242254 241440 242310 241496
rect 244278 240796 244280 240816
rect 244280 240796 244332 240816
rect 244332 240796 244334 240816
rect 244278 240760 244334 240796
rect 241610 240080 241666 240136
rect 240230 149368 240286 149424
rect 240230 120264 240286 120320
rect 238114 78376 238170 78432
rect 245658 241440 245714 241496
rect 243542 89528 243598 89584
rect 241610 80008 241666 80064
rect 248418 239672 248474 239728
rect 246394 237904 246450 237960
rect 246302 226208 246358 226264
rect 245658 146104 245714 146160
rect 248418 226888 248474 226944
rect 246486 146104 246542 146160
rect 246486 144880 246542 144936
rect 250442 240080 250498 240136
rect 250350 232600 250406 232656
rect 251270 239808 251326 239864
rect 250442 228928 250498 228984
rect 251914 230424 251970 230480
rect 254582 318008 254638 318064
rect 254582 314064 254638 314120
rect 253938 313928 253994 313984
rect 253662 301280 253718 301336
rect 253110 298968 253166 299024
rect 253202 296928 253258 296984
rect 253018 296520 253074 296576
rect 253202 289856 253258 289912
rect 253846 289584 253902 289640
rect 252834 285368 252890 285424
rect 253662 283872 253718 283928
rect 252926 266328 252982 266384
rect 252834 253136 252890 253192
rect 254214 308488 254270 308544
rect 254122 263200 254178 263256
rect 253938 253680 253994 253736
rect 253938 249464 253994 249520
rect 252834 242800 252890 242856
rect 252742 239944 252798 240000
rect 252926 242392 252982 242448
rect 252650 229880 252706 229936
rect 252742 182824 252798 182880
rect 258078 467880 258134 467936
rect 255962 454008 256018 454064
rect 255962 448840 256018 448896
rect 255686 446120 255742 446176
rect 255410 443400 255466 443456
rect 255410 439048 255466 439104
rect 255502 437688 255558 437744
rect 255502 436736 255558 436792
rect 255410 434968 255466 435024
rect 255410 433608 255466 433664
rect 256054 446120 256110 446176
rect 255594 430616 255650 430672
rect 255410 427896 255466 427952
rect 255502 426536 255558 426592
rect 256606 429256 256662 429312
rect 256606 425176 256662 425232
rect 258170 452648 258226 452704
rect 255502 423544 255558 423600
rect 255502 422184 255558 422240
rect 255594 420824 255650 420880
rect 255502 419464 255558 419520
rect 255594 418104 255650 418160
rect 255502 416780 255504 416800
rect 255504 416780 255556 416800
rect 255556 416780 255558 416800
rect 255502 416744 255558 416780
rect 256606 415112 256662 415168
rect 255502 412392 255558 412448
rect 255502 411032 255558 411088
rect 255502 409672 255558 409728
rect 255502 408312 255558 408368
rect 255502 406952 255558 407008
rect 255502 403960 255558 404016
rect 255502 401240 255558 401296
rect 255502 399880 255558 399936
rect 255502 398520 255558 398576
rect 255502 396888 255558 396944
rect 255594 394168 255650 394224
rect 256698 377304 256754 377360
rect 258078 386416 258134 386472
rect 255502 328344 255558 328400
rect 254766 313928 254822 313984
rect 255594 295024 255650 295080
rect 255502 293800 255558 293856
rect 255410 292576 255466 292632
rect 255410 292204 255412 292224
rect 255412 292204 255464 292224
rect 255464 292204 255466 292224
rect 255410 292168 255466 292204
rect 255410 290808 255466 290864
rect 256606 300736 256662 300792
rect 256514 300328 256570 300384
rect 256606 298288 256662 298344
rect 256606 297880 256662 297936
rect 256514 297472 256570 297528
rect 255870 297064 255926 297120
rect 256606 296928 256662 296984
rect 256606 295432 256662 295488
rect 256606 295044 256662 295080
rect 256606 295024 256608 295044
rect 256608 295024 256660 295044
rect 256660 295024 256662 295044
rect 256606 294208 256662 294264
rect 255686 293392 255742 293448
rect 256606 292984 256662 293040
rect 255318 287544 255374 287600
rect 255502 288768 255558 288824
rect 255502 287136 255558 287192
rect 255042 263236 255044 263256
rect 255044 263236 255096 263256
rect 255096 263236 255098 263256
rect 255042 263200 255098 263236
rect 254582 259528 254638 259584
rect 254582 258440 254638 258496
rect 255226 254768 255282 254824
rect 255226 254360 255282 254416
rect 254950 249464 255006 249520
rect 254582 248648 254638 248704
rect 254214 247424 254270 247480
rect 255502 286320 255558 286376
rect 255410 285912 255466 285968
rect 255410 285504 255466 285560
rect 255410 284280 255466 284336
rect 255502 283056 255558 283112
rect 255502 282648 255558 282704
rect 255410 281868 255412 281888
rect 255412 281868 255464 281888
rect 255464 281868 255466 281888
rect 255410 281832 255466 281868
rect 255410 281324 255412 281344
rect 255412 281324 255464 281344
rect 255464 281324 255466 281344
rect 255410 281288 255466 281324
rect 255410 280472 255466 280528
rect 255410 280100 255412 280120
rect 255412 280100 255464 280120
rect 255464 280100 255466 280120
rect 255410 280064 255466 280100
rect 256790 325760 256846 325816
rect 256790 289992 256846 290048
rect 256974 298696 257030 298752
rect 258722 403552 258778 403608
rect 258354 382200 258410 382256
rect 258262 375264 258318 375320
rect 260930 460944 260986 461000
rect 259458 316512 259514 316568
rect 257066 291760 257122 291816
rect 256882 284688 256938 284744
rect 256698 279248 256754 279304
rect 255502 278840 255558 278896
rect 255410 277616 255466 277672
rect 255410 276392 255466 276448
rect 255502 275984 255558 276040
rect 255410 275168 255466 275224
rect 255410 274760 255466 274816
rect 255410 274352 255466 274408
rect 255502 273944 255558 274000
rect 255410 273148 255466 273184
rect 255410 273128 255412 273148
rect 255412 273128 255464 273148
rect 255464 273128 255466 273148
rect 255502 272720 255558 272776
rect 256882 271904 256938 271960
rect 255410 271360 255466 271416
rect 255410 270564 255466 270600
rect 255410 270544 255412 270564
rect 255412 270544 255464 270564
rect 255464 270544 255466 270564
rect 255502 270136 255558 270192
rect 255410 269728 255466 269784
rect 256698 269320 256754 269376
rect 255410 268948 255412 268968
rect 255412 268948 255464 268968
rect 255464 268948 255466 268968
rect 255410 268912 255466 268948
rect 255502 268096 255558 268152
rect 255502 267688 255558 267744
rect 255410 266872 255466 266928
rect 255502 266056 255558 266112
rect 255410 265240 255466 265296
rect 255594 264832 255650 264888
rect 255410 264424 255466 264480
rect 255410 264016 255466 264072
rect 255502 263744 255558 263800
rect 255502 262384 255558 262440
rect 255410 260616 255466 260672
rect 255594 260208 255650 260264
rect 255410 259412 255466 259448
rect 255410 259392 255412 259412
rect 255412 259392 255464 259412
rect 255464 259392 255466 259412
rect 255594 258712 255650 258768
rect 255502 258576 255558 258632
rect 255410 257388 255412 257408
rect 255412 257388 255464 257408
rect 255464 257388 255466 257408
rect 255410 257352 255466 257388
rect 255410 256944 255466 257000
rect 255410 256536 255466 256592
rect 255594 256128 255650 256184
rect 255502 255312 255558 255368
rect 255410 254496 255466 254552
rect 255594 254496 255650 254552
rect 255502 254088 255558 254144
rect 255410 252864 255466 252920
rect 255410 252456 255466 252512
rect 255502 252048 255558 252104
rect 255502 251096 255558 251152
rect 255870 249908 255872 249928
rect 255872 249908 255924 249928
rect 255924 249908 255926 249928
rect 255870 249872 255926 249908
rect 255410 249076 255466 249112
rect 255410 249056 255412 249076
rect 255412 249056 255464 249076
rect 255464 249056 255466 249076
rect 255502 247016 255558 247072
rect 255410 246608 255466 246664
rect 255686 246200 255742 246256
rect 255410 245812 255466 245848
rect 255410 245792 255412 245812
rect 255412 245792 255464 245812
rect 255464 245792 255466 245812
rect 255410 245384 255466 245440
rect 255594 244976 255650 245032
rect 255502 244568 255558 244624
rect 255410 244196 255412 244216
rect 255412 244196 255464 244216
rect 255464 244196 255466 244216
rect 255410 244160 255466 244196
rect 255502 243752 255558 243808
rect 255410 240896 255466 240952
rect 255594 242256 255650 242312
rect 255594 240780 255650 240816
rect 256054 242120 256110 242176
rect 255594 240760 255596 240780
rect 255596 240760 255648 240780
rect 255648 240760 255650 240780
rect 255410 236544 255466 236600
rect 255962 214512 256018 214568
rect 253294 139984 253350 140040
rect 251270 91840 251326 91896
rect 251270 91160 251326 91216
rect 251822 91160 251878 91216
rect 256054 207576 256110 207632
rect 255318 204992 255374 205048
rect 255962 204992 256018 205048
rect 255318 90888 255374 90944
rect 258170 283464 258226 283520
rect 258262 280744 258318 280800
rect 263598 450200 263654 450256
rect 260930 376488 260986 376544
rect 261482 376488 261538 376544
rect 261482 363024 261538 363080
rect 260102 305768 260158 305824
rect 259734 302776 259790 302832
rect 258814 280880 258870 280936
rect 258722 279656 258778 279712
rect 258078 276800 258134 276856
rect 257342 269728 257398 269784
rect 257342 240760 257398 240816
rect 257250 239672 257306 239728
rect 256790 235184 256846 235240
rect 256054 153040 256110 153096
rect 258262 270564 258318 270600
rect 258262 270544 258264 270564
rect 258264 270544 258316 270564
rect 258316 270544 258318 270564
rect 258538 251504 258594 251560
rect 258262 241032 258318 241088
rect 258078 213152 258134 213208
rect 259550 277208 259606 277264
rect 259458 273148 259514 273184
rect 259458 273128 259460 273148
rect 259460 273128 259512 273148
rect 259512 273128 259514 273148
rect 259274 265512 259330 265568
rect 258722 212472 258778 212528
rect 256698 89664 256754 89720
rect 259734 265648 259790 265704
rect 260746 259412 260802 259448
rect 260746 259392 260748 259412
rect 260748 259392 260800 259412
rect 260800 259392 260802 259412
rect 259734 240896 259790 240952
rect 261114 312432 261170 312488
rect 263598 320048 263654 320104
rect 263782 386280 263838 386336
rect 263782 320048 263838 320104
rect 263782 318960 263838 319016
rect 263690 318824 263746 318880
rect 262862 313928 262918 313984
rect 262310 277208 262366 277264
rect 260930 273808 260986 273864
rect 259550 86128 259606 86184
rect 263598 290672 263654 290728
rect 262310 207576 262366 207632
rect 262678 247832 262734 247888
rect 262218 94696 262274 94752
rect 262218 76472 262274 76528
rect 263690 285504 263746 285560
rect 263690 277888 263746 277944
rect 265070 305632 265126 305688
rect 264886 296928 264942 296984
rect 263874 288224 263930 288280
rect 263782 270816 263838 270872
rect 263874 263744 263930 263800
rect 266450 387640 266506 387696
rect 266450 339516 266506 339552
rect 266450 339496 266452 339516
rect 266452 339496 266504 339516
rect 266504 339496 266506 339516
rect 266358 298016 266414 298072
rect 265346 285368 265402 285424
rect 265346 284280 265402 284336
rect 266358 284280 266414 284336
rect 265070 258848 265126 258904
rect 265070 258576 265126 258632
rect 265622 242800 265678 242856
rect 265070 189624 265126 189680
rect 266450 283464 266506 283520
rect 267738 309304 267794 309360
rect 266634 278296 266690 278352
rect 267922 308352 267978 308408
rect 267922 291760 267978 291816
rect 267738 272176 267794 272232
rect 266818 267028 266874 267064
rect 266818 267008 266820 267028
rect 266820 267008 266872 267028
rect 266872 267008 266874 267028
rect 267186 264832 267242 264888
rect 266910 255176 266966 255232
rect 266634 227024 266690 227080
rect 269118 309032 269174 309088
rect 269118 304952 269174 305008
rect 269118 295296 269174 295352
rect 268014 267960 268070 268016
rect 269026 248412 269028 248432
rect 269028 248412 269080 248432
rect 269080 248412 269082 248432
rect 269026 248376 269082 248412
rect 270590 321544 270646 321600
rect 269394 309032 269450 309088
rect 269394 307808 269450 307864
rect 270590 287408 270646 287464
rect 270498 287000 270554 287056
rect 270590 273808 270646 273864
rect 270498 272176 270554 272232
rect 269854 263608 269910 263664
rect 269394 252592 269450 252648
rect 271878 320592 271934 320648
rect 270774 289040 270830 289096
rect 270682 259528 270738 259584
rect 270682 254360 270738 254416
rect 270498 151680 270554 151736
rect 272154 320592 272210 320648
rect 272154 320184 272210 320240
rect 272062 298016 272118 298072
rect 271970 251096 272026 251152
rect 271970 250552 272026 250608
rect 273258 299512 273314 299568
rect 272522 299412 272524 299432
rect 272524 299412 272576 299432
rect 272576 299412 272578 299432
rect 272522 299376 272578 299412
rect 272154 265512 272210 265568
rect 272154 250688 272210 250744
rect 270590 97416 270646 97472
rect 269210 92520 269266 92576
rect 269118 75792 269174 75848
rect 273534 255584 273590 255640
rect 273350 234504 273406 234560
rect 274914 280744 274970 280800
rect 273534 220224 273590 220280
rect 276202 380840 276258 380896
rect 276202 379480 276258 379536
rect 276202 277888 276258 277944
rect 276018 135904 276074 135960
rect 273350 78512 273406 78568
rect 277674 306448 277730 306504
rect 277582 282104 277638 282160
rect 277398 268368 277454 268424
rect 277398 266736 277454 266792
rect 278778 302368 278834 302424
rect 278134 258712 278190 258768
rect 278870 295160 278926 295216
rect 278870 293936 278926 293992
rect 278870 287408 278926 287464
rect 278962 254496 279018 254552
rect 280250 311208 280306 311264
rect 280342 311072 280398 311128
rect 281446 311208 281502 311264
rect 280802 311072 280858 311128
rect 280434 296656 280490 296712
rect 280434 295296 280490 295352
rect 278870 146240 278926 146296
rect 559654 702480 559710 702536
rect 580906 697176 580962 697232
rect 582378 683848 582434 683904
rect 580170 577632 580226 577688
rect 580170 484608 580226 484664
rect 284390 458360 284446 458416
rect 282182 388320 282238 388376
rect 282918 382916 282920 382936
rect 282920 382916 282972 382936
rect 282972 382916 282974 382936
rect 282918 382880 282974 382916
rect 281722 271088 281778 271144
rect 282918 303592 282974 303648
rect 281538 82728 281594 82784
rect 283102 255584 283158 255640
rect 283010 247696 283066 247752
rect 285678 386280 285734 386336
rect 284574 367648 284630 367704
rect 284482 295296 284538 295352
rect 284390 242800 284446 242856
rect 284390 242120 284446 242176
rect 285678 293936 285734 293992
rect 284574 242800 284630 242856
rect 284666 233144 284722 233200
rect 284482 163376 284538 163432
rect 284390 88032 284446 88088
rect 287058 456864 287114 456920
rect 288346 456864 288402 456920
rect 288438 453056 288494 453112
rect 287150 451288 287206 451344
rect 285954 146920 286010 146976
rect 288438 219136 288494 219192
rect 289818 366968 289874 367024
rect 288622 86808 288678 86864
rect 288438 71032 288494 71088
rect 285678 60560 285734 60616
rect 286414 60560 286470 60616
rect 289726 86808 289782 86864
rect 289726 85584 289782 85640
rect 580170 458088 580226 458144
rect 582654 670656 582710 670712
rect 582470 644000 582526 644056
rect 582378 431568 582434 431624
rect 582562 630808 582618 630864
rect 582838 617480 582894 617536
rect 582746 590960 582802 591016
rect 582654 458768 582710 458824
rect 582562 390496 582618 390552
rect 582470 383832 582526 383888
rect 582470 378392 582526 378448
rect 582378 376624 582434 376680
rect 582378 365064 582434 365120
rect 291658 269728 291714 269784
rect 580262 325216 580318 325272
rect 580170 298696 580226 298752
rect 580170 272176 580226 272232
rect 580170 258848 580226 258904
rect 582930 564304 582986 564360
rect 582838 524456 582894 524512
rect 583022 537784 583078 537840
rect 583206 511264 583262 511320
rect 583114 471416 583170 471472
rect 582930 418240 582986 418296
rect 583206 451288 583262 451344
rect 583206 404912 583262 404968
rect 582654 351872 582710 351928
rect 582562 312024 582618 312080
rect 582470 302232 582526 302288
rect 582378 245520 582434 245576
rect 580170 232328 580226 232384
rect 579894 219000 579950 219056
rect 582378 215872 582434 215928
rect 580262 205672 580318 205728
rect 295430 144064 295486 144120
rect 303618 163376 303674 163432
rect 302238 144064 302294 144120
rect 301962 7520 302018 7576
rect 305642 6160 305698 6216
rect 309782 84224 309838 84280
rect 335358 155216 335414 155272
rect 319718 6160 319774 6216
rect 327078 80688 327134 80744
rect 348054 3440 348110 3496
rect 353298 3440 353354 3496
rect 580170 192480 580226 192536
rect 580170 179152 580226 179208
rect 580262 88984 580318 89040
rect 580262 72936 580318 72992
rect 580170 46280 580226 46336
rect 582562 250416 582618 250472
rect 582562 152632 582618 152688
rect 582838 165824 582894 165880
rect 582746 139304 582802 139360
rect 583022 140800 583078 140856
rect 582930 125976 582986 126032
rect 582654 112784 582710 112840
rect 582654 99456 582710 99512
rect 582930 87488 582986 87544
rect 582654 78512 582710 78568
rect 582838 33088 582894 33144
rect 582562 19760 582618 19816
rect 583022 59608 583078 59664
rect 582930 6568 582986 6624
<< metal3 >>
rect 258574 702476 258580 702540
rect 258644 702538 258650 702540
rect 559649 702538 559715 702541
rect 258644 702536 559715 702538
rect 258644 702480 559654 702536
rect 559710 702480 559715 702536
rect 258644 702478 559715 702480
rect 258644 702476 258650 702478
rect 559649 702475 559715 702478
rect -960 697220 480 697460
rect 580901 697234 580967 697237
rect 583520 697234 584960 697324
rect 580901 697232 584960 697234
rect 580901 697176 580906 697232
rect 580962 697176 584960 697232
rect 580901 697174 584960 697176
rect 580901 697171 580967 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 582373 683906 582439 683909
rect 583520 683906 584960 683996
rect 582373 683904 584960 683906
rect 582373 683848 582378 683904
rect 582434 683848 584960 683904
rect 582373 683846 584960 683848
rect 582373 683843 582439 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 582649 670714 582715 670717
rect 583520 670714 584960 670804
rect 582649 670712 584960 670714
rect 582649 670656 582654 670712
rect 582710 670656 584960 670712
rect 582649 670654 584960 670656
rect 582649 670651 582715 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 582465 644058 582531 644061
rect 583520 644058 584960 644148
rect 582465 644056 584960 644058
rect 582465 644000 582470 644056
rect 582526 644000 584960 644056
rect 582465 643998 584960 644000
rect 582465 643995 582531 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 582557 630866 582623 630869
rect 583520 630866 584960 630956
rect 582557 630864 584960 630866
rect 582557 630808 582562 630864
rect 582618 630808 584960 630864
rect 582557 630806 584960 630808
rect 582557 630803 582623 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3509 619170 3575 619173
rect -960 619168 3575 619170
rect -960 619112 3514 619168
rect 3570 619112 3575 619168
rect -960 619110 3575 619112
rect -960 619020 480 619110
rect 3509 619107 3575 619110
rect 582833 617538 582899 617541
rect 583520 617538 584960 617628
rect 582833 617536 584960 617538
rect 582833 617480 582838 617536
rect 582894 617480 584960 617536
rect 582833 617478 584960 617480
rect 582833 617475 582899 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 2773 606114 2839 606117
rect -960 606112 2839 606114
rect -960 606056 2778 606112
rect 2834 606056 2839 606112
rect -960 606054 2839 606056
rect -960 605964 480 606054
rect 2773 606051 2839 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 582741 591018 582807 591021
rect 583520 591018 584960 591108
rect 582741 591016 584960 591018
rect 582741 590960 582746 591016
rect 582802 590960 584960 591016
rect 582741 590958 584960 590960
rect 582741 590955 582807 590958
rect 583520 590868 584960 590958
rect 71773 585170 71839 585173
rect 75862 585170 75868 585172
rect 71773 585168 75868 585170
rect 71773 585112 71778 585168
rect 71834 585112 75868 585168
rect 71773 585110 75868 585112
rect 71773 585107 71839 585110
rect 75862 585108 75868 585110
rect 75932 585108 75938 585172
rect 92105 583810 92171 583813
rect 119337 583810 119403 583813
rect 92105 583808 119403 583810
rect 92105 583752 92110 583808
rect 92166 583752 119342 583808
rect 119398 583752 119403 583808
rect 92105 583750 119403 583752
rect 92105 583747 92171 583750
rect 119337 583747 119403 583750
rect 85481 582722 85547 582725
rect 133137 582722 133203 582725
rect 85481 582720 133203 582722
rect 85481 582664 85486 582720
rect 85542 582664 133142 582720
rect 133198 582664 133203 582720
rect 85481 582662 133203 582664
rect 85481 582659 85547 582662
rect 133137 582659 133203 582662
rect 73521 582586 73587 582589
rect 107009 582586 107075 582589
rect 73521 582584 107075 582586
rect 73521 582528 73526 582584
rect 73582 582528 107014 582584
rect 107070 582528 107075 582584
rect 73521 582526 107075 582528
rect 73521 582523 73587 582526
rect 107009 582523 107075 582526
rect 80237 581226 80303 581229
rect 80646 581226 80652 581228
rect 64830 581224 80652 581226
rect 64830 581168 80242 581224
rect 80298 581168 80652 581224
rect 64830 581166 80652 581168
rect 8109 581090 8175 581093
rect 64830 581090 64890 581166
rect 80237 581163 80303 581166
rect 80646 581164 80652 581166
rect 80716 581164 80722 581228
rect 8109 581088 64890 581090
rect 8109 581032 8114 581088
rect 8170 581032 64890 581088
rect 8109 581030 64890 581032
rect 75361 581090 75427 581093
rect 75678 581090 75684 581092
rect 75361 581088 75684 581090
rect 75361 581032 75366 581088
rect 75422 581032 75684 581088
rect 75361 581030 75684 581032
rect 8109 581027 8175 581030
rect 75361 581027 75427 581030
rect 75678 581028 75684 581030
rect 75748 581028 75754 581092
rect 82721 581090 82787 581093
rect 101254 581090 101260 581092
rect 82721 581088 101260 581090
rect 82721 581032 82726 581088
rect 82782 581032 101260 581088
rect 82721 581030 101260 581032
rect 82721 581027 82787 581030
rect 101254 581028 101260 581030
rect 101324 581028 101330 581092
rect 70342 580756 70348 580820
rect 70412 580818 70418 580820
rect 70853 580818 70919 580821
rect 70412 580816 70919 580818
rect 70412 580760 70858 580816
rect 70914 580760 70919 580816
rect 70412 580758 70919 580760
rect 70412 580756 70418 580758
rect 70853 580755 70919 580758
rect 79869 580820 79935 580821
rect 79869 580816 79916 580820
rect 79980 580818 79986 580820
rect 79869 580760 79874 580816
rect 79869 580756 79916 580760
rect 79980 580758 80026 580818
rect 79980 580756 79986 580758
rect 83958 580756 83964 580820
rect 84028 580818 84034 580820
rect 84193 580818 84259 580821
rect 84028 580816 84259 580818
rect 84028 580760 84198 580816
rect 84254 580760 84259 580816
rect 84028 580758 84259 580760
rect 84028 580756 84034 580758
rect 79869 580755 79935 580756
rect 84193 580755 84259 580758
rect 88885 580820 88951 580821
rect 92565 580820 92631 580821
rect 88885 580816 88932 580820
rect 88996 580818 89002 580820
rect 88885 580760 88890 580816
rect 88885 580756 88932 580760
rect 88996 580758 89042 580818
rect 92565 580816 92612 580820
rect 92676 580818 92682 580820
rect 92565 580760 92570 580816
rect 88996 580756 89002 580758
rect 92565 580756 92612 580760
rect 92676 580758 92722 580818
rect 92676 580756 92682 580758
rect 88885 580755 88951 580756
rect 92565 580755 92631 580756
rect -960 580002 480 580092
rect 3509 580002 3575 580005
rect -960 580000 3575 580002
rect -960 579944 3514 580000
rect 3570 579944 3575 580000
rect -960 579942 3575 579944
rect -960 579852 480 579942
rect 3509 579939 3575 579942
rect 66529 580002 66595 580005
rect 68878 580002 68938 580584
rect 66529 580000 68938 580002
rect 66529 579944 66534 580000
rect 66590 579944 68938 580000
rect 66529 579942 68938 579944
rect 66529 579939 66595 579942
rect 67541 578642 67607 578645
rect 68878 578642 68938 579224
rect 94638 578914 94698 579496
rect 97165 578914 97231 578917
rect 94638 578912 97231 578914
rect 94638 578856 97170 578912
rect 97226 578856 97231 578912
rect 94638 578854 97231 578856
rect 97165 578851 97231 578854
rect 67541 578640 68938 578642
rect 67541 578584 67546 578640
rect 67602 578584 68938 578640
rect 67541 578582 68938 578584
rect 67541 578579 67607 578582
rect 67449 577282 67515 577285
rect 68878 577282 68938 577864
rect 94638 577554 94698 578136
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 97165 577554 97231 577557
rect 94638 577552 97231 577554
rect 94638 577496 97170 577552
rect 97226 577496 97231 577552
rect 583520 577540 584960 577630
rect 94638 577494 97231 577496
rect 97165 577491 97231 577494
rect 67449 577280 68938 577282
rect 67449 577224 67454 577280
rect 67510 577224 68938 577280
rect 67449 577222 68938 577224
rect 67449 577219 67515 577222
rect 67633 575922 67699 575925
rect 68878 575922 68938 576504
rect 94638 576466 94698 576776
rect 97901 576466 97967 576469
rect 94638 576464 97967 576466
rect 94638 576408 97906 576464
rect 97962 576408 97967 576464
rect 94638 576406 97967 576408
rect 97901 576403 97967 576406
rect 67633 575920 68938 575922
rect 67633 575864 67638 575920
rect 67694 575864 68938 575920
rect 67633 575862 68938 575864
rect 67633 575859 67699 575862
rect 67725 575378 67791 575381
rect 67725 575376 68938 575378
rect 67725 575320 67730 575376
rect 67786 575320 68938 575376
rect 67725 575318 68938 575320
rect 67725 575315 67791 575318
rect 68878 575144 68938 575318
rect 94638 574834 94698 575416
rect 95233 574834 95299 574837
rect 94638 574832 95299 574834
rect 94638 574776 95238 574832
rect 95294 574776 95299 574832
rect 94638 574774 95299 574776
rect 95233 574771 95299 574774
rect 66529 573202 66595 573205
rect 68878 573202 68938 573784
rect 94638 573474 94698 574056
rect 97901 573474 97967 573477
rect 94638 573472 97967 573474
rect 94638 573416 97906 573472
rect 97962 573416 97967 573472
rect 94638 573414 97967 573416
rect 97901 573411 97967 573414
rect 66529 573200 68938 573202
rect 66529 573144 66534 573200
rect 66590 573144 68938 573200
rect 66529 573142 68938 573144
rect 66529 573139 66595 573142
rect 66529 571842 66595 571845
rect 68878 571842 68938 572424
rect 94638 572114 94698 572696
rect 96797 572114 96863 572117
rect 94638 572112 96863 572114
rect 94638 572056 96802 572112
rect 96858 572056 96863 572112
rect 94638 572054 96863 572056
rect 96797 572051 96863 572054
rect 66529 571840 68938 571842
rect 66529 571784 66534 571840
rect 66590 571784 68938 571840
rect 66529 571782 68938 571784
rect 66529 571779 66595 571782
rect 97257 571434 97323 571437
rect 94638 571432 97323 571434
rect 94638 571376 97262 571432
rect 97318 571376 97323 571432
rect 94638 571374 97323 571376
rect 94638 571336 94698 571374
rect 97257 571371 97323 571374
rect 66897 570210 66963 570213
rect 68878 570210 68938 570792
rect 66897 570208 68938 570210
rect 66897 570152 66902 570208
rect 66958 570152 68938 570208
rect 66897 570150 68938 570152
rect 66897 570147 66963 570150
rect 97901 570074 97967 570077
rect 94638 570072 97967 570074
rect 94638 570016 97906 570072
rect 97962 570016 97967 570072
rect 94638 570014 97967 570016
rect 94638 569976 94698 570014
rect 97901 570011 97967 570014
rect 67357 568850 67423 568853
rect 68878 568850 68938 569432
rect 67357 568848 68938 568850
rect 67357 568792 67362 568848
rect 67418 568792 68938 568848
rect 67357 568790 68938 568792
rect 67357 568787 67423 568790
rect 96705 568714 96771 568717
rect 97901 568714 97967 568717
rect 94638 568712 97967 568714
rect 94638 568656 96710 568712
rect 96766 568656 97906 568712
rect 97962 568656 97967 568712
rect 94638 568654 97967 568656
rect 94638 568616 94698 568654
rect 96705 568651 96771 568654
rect 97901 568651 97967 568654
rect 65977 567626 66043 567629
rect 68878 567626 68938 568072
rect 65977 567624 68938 567626
rect 65977 567568 65982 567624
rect 66038 567568 68938 567624
rect 65977 567566 68938 567568
rect 65977 567563 66043 567566
rect 94638 567218 94698 567256
rect 95601 567218 95667 567221
rect 94638 567216 95667 567218
rect 94638 567160 95606 567216
rect 95662 567160 95667 567216
rect 94638 567158 95667 567160
rect 95601 567155 95667 567158
rect -960 566946 480 567036
rect 3417 566946 3483 566949
rect -960 566944 3483 566946
rect -960 566888 3422 566944
rect 3478 566888 3483 566944
rect -960 566886 3483 566888
rect -960 566796 480 566886
rect 3417 566883 3483 566886
rect 66161 566810 66227 566813
rect 66161 566808 68938 566810
rect 66161 566752 66166 566808
rect 66222 566752 68938 566808
rect 66161 566750 68938 566752
rect 66161 566747 66227 566750
rect 68878 566712 68938 566750
rect 94638 565858 94698 565896
rect 96705 565858 96771 565861
rect 94638 565856 96771 565858
rect 94638 565800 96710 565856
rect 96766 565800 96771 565856
rect 94638 565798 96771 565800
rect 96705 565795 96771 565798
rect 97257 565858 97323 565861
rect 104934 565858 104940 565860
rect 97257 565856 104940 565858
rect 97257 565800 97262 565856
rect 97318 565800 104940 565856
rect 97257 565798 104940 565800
rect 97257 565795 97323 565798
rect 104934 565796 104940 565798
rect 105004 565796 105010 565860
rect 66529 564770 66595 564773
rect 68878 564770 68938 565352
rect 66529 564768 68938 564770
rect 66529 564712 66534 564768
rect 66590 564712 68938 564768
rect 66529 564710 68938 564712
rect 66529 564707 66595 564710
rect 582925 564362 582991 564365
rect 583520 564362 584960 564452
rect 582925 564360 584960 564362
rect 582925 564304 582930 564360
rect 582986 564304 584960 564360
rect 582925 564302 584960 564304
rect 582925 564299 582991 564302
rect 66529 563410 66595 563413
rect 68878 563410 68938 563992
rect 94638 563682 94698 564264
rect 583520 564212 584960 564302
rect 95417 563682 95483 563685
rect 94638 563680 95483 563682
rect 94638 563624 95422 563680
rect 95478 563624 95483 563680
rect 94638 563622 95483 563624
rect 95417 563619 95483 563622
rect 66529 563408 68938 563410
rect 66529 563352 66534 563408
rect 66590 563352 68938 563408
rect 66529 563350 68938 563352
rect 66529 563347 66595 563350
rect 67766 561988 67772 562052
rect 67836 562050 67842 562052
rect 68878 562050 68938 562632
rect 94638 562322 94698 562904
rect 96797 562322 96863 562325
rect 94638 562320 96863 562322
rect 94638 562264 96802 562320
rect 96858 562264 96863 562320
rect 94638 562262 96863 562264
rect 96797 562259 96863 562262
rect 67836 561990 68938 562050
rect 67836 561988 67842 561990
rect 66713 560690 66779 560693
rect 68878 560690 68938 561272
rect 94638 560962 94698 561544
rect 96889 560962 96955 560965
rect 94638 560960 96955 560962
rect 94638 560904 96894 560960
rect 96950 560904 96955 560960
rect 94638 560902 96955 560904
rect 96889 560899 96955 560902
rect 66713 560688 68938 560690
rect 66713 560632 66718 560688
rect 66774 560632 68938 560688
rect 66713 560630 68938 560632
rect 66713 560627 66779 560630
rect 66713 559330 66779 559333
rect 68878 559330 68938 559912
rect 94638 559602 94698 560184
rect 96797 559602 96863 559605
rect 94638 559600 96863 559602
rect 94638 559544 96802 559600
rect 96858 559544 96863 559600
rect 94638 559542 96863 559544
rect 96797 559539 96863 559542
rect 66713 559328 68938 559330
rect 66713 559272 66718 559328
rect 66774 559272 68938 559328
rect 66713 559270 68938 559272
rect 66713 559267 66779 559270
rect 94638 558653 94698 558824
rect 94638 558650 94747 558653
rect 95509 558650 95575 558653
rect 94638 558648 95575 558650
rect 94638 558592 94686 558648
rect 94742 558592 95514 558648
rect 95570 558592 95575 558648
rect 94638 558590 95575 558592
rect 94681 558587 94747 558590
rect 95509 558587 95575 558590
rect 66713 557970 66779 557973
rect 68878 557970 68938 558552
rect 66713 557968 68938 557970
rect 66713 557912 66718 557968
rect 66774 557912 68938 557968
rect 66713 557910 68938 557912
rect 66713 557907 66779 557910
rect 67725 556610 67791 556613
rect 68878 556610 68938 557192
rect 94638 556882 94698 557464
rect 96797 556882 96863 556885
rect 94638 556880 96863 556882
rect 94638 556824 96802 556880
rect 96858 556824 96863 556880
rect 94638 556822 96863 556824
rect 96797 556819 96863 556822
rect 67725 556608 68938 556610
rect 67725 556552 67730 556608
rect 67786 556552 68938 556608
rect 67725 556550 68938 556552
rect 67725 556547 67791 556550
rect 66069 555250 66135 555253
rect 68878 555250 68938 555832
rect 94638 555522 94698 556104
rect 96981 555522 97047 555525
rect 94638 555520 97047 555522
rect 94638 555464 96986 555520
rect 97042 555464 97047 555520
rect 94638 555462 97047 555464
rect 96981 555459 97047 555462
rect 66069 555248 68938 555250
rect 66069 555192 66074 555248
rect 66130 555192 68938 555248
rect 66069 555190 68938 555192
rect 66069 555187 66135 555190
rect -960 553890 480 553980
rect 3325 553890 3391 553893
rect -960 553888 3391 553890
rect -960 553832 3330 553888
rect 3386 553832 3391 553888
rect -960 553830 3391 553832
rect -960 553740 480 553830
rect 3325 553827 3391 553830
rect 66529 553754 66595 553757
rect 68878 553754 68938 554200
rect 94638 554162 94698 554744
rect 96654 554162 96660 554164
rect 94638 554102 96660 554162
rect 96654 554100 96660 554102
rect 96724 554100 96730 554164
rect 66529 553752 68938 553754
rect 66529 553696 66534 553752
rect 66590 553696 68938 553752
rect 66529 553694 68938 553696
rect 66529 553691 66595 553694
rect 67817 552258 67883 552261
rect 68878 552258 68938 552840
rect 94638 552802 94698 553384
rect 96981 552802 97047 552805
rect 94638 552800 97047 552802
rect 94638 552744 96986 552800
rect 97042 552744 97047 552800
rect 94638 552742 97047 552744
rect 96981 552739 97047 552742
rect 96613 552530 96679 552533
rect 67817 552256 68938 552258
rect 67817 552200 67822 552256
rect 67878 552200 68938 552256
rect 67817 552198 68938 552200
rect 94638 552528 96679 552530
rect 94638 552472 96618 552528
rect 96674 552472 96679 552528
rect 94638 552470 96679 552472
rect 94638 552261 94698 552470
rect 96613 552467 96679 552470
rect 94638 552258 94747 552261
rect 94638 552256 94828 552258
rect 94638 552200 94686 552256
rect 94742 552200 94828 552256
rect 94638 552198 94828 552200
rect 67817 552195 67883 552198
rect 94638 552195 94747 552198
rect 94638 552024 94698 552195
rect 65885 550898 65951 550901
rect 68878 550898 68938 551480
rect 583520 551020 584960 551260
rect 65885 550896 68938 550898
rect 65885 550840 65890 550896
rect 65946 550840 68938 550896
rect 65885 550838 68938 550840
rect 65885 550835 65951 550838
rect 97901 550762 97967 550765
rect 94638 550760 97967 550762
rect 94638 550704 97906 550760
rect 97962 550704 97967 550760
rect 94638 550702 97967 550704
rect 94638 550664 94698 550702
rect 97901 550699 97967 550702
rect 66529 549674 66595 549677
rect 68878 549674 68938 550120
rect 66529 549672 68938 549674
rect 66529 549616 66534 549672
rect 66590 549616 68938 549672
rect 66529 549614 68938 549616
rect 66529 549611 66595 549614
rect 100702 549402 100708 549404
rect 94638 549342 100708 549402
rect 94638 549304 94698 549342
rect 100702 549340 100708 549342
rect 100772 549340 100778 549404
rect 66805 548178 66871 548181
rect 68878 548178 68938 548760
rect 66805 548176 68938 548178
rect 66805 548120 66810 548176
rect 66866 548120 68938 548176
rect 66805 548118 68938 548120
rect 66805 548115 66871 548118
rect 69062 546820 69122 547400
rect 94638 547090 94698 547672
rect 96838 547090 96844 547092
rect 94638 547030 96844 547090
rect 96838 547028 96844 547030
rect 96908 547028 96914 547092
rect 69054 546756 69060 546820
rect 69124 546756 69130 546820
rect 66713 545458 66779 545461
rect 68878 545458 68938 546040
rect 94638 545730 94698 546312
rect 96981 545730 97047 545733
rect 94638 545728 97047 545730
rect 94638 545672 96986 545728
rect 97042 545672 97047 545728
rect 94638 545670 97047 545672
rect 96981 545667 97047 545670
rect 66713 545456 68938 545458
rect 66713 545400 66718 545456
rect 66774 545400 68938 545456
rect 66713 545398 68938 545400
rect 66713 545395 66779 545398
rect 65793 544098 65859 544101
rect 68878 544098 68938 544680
rect 94638 544370 94698 544952
rect 97073 544370 97139 544373
rect 94638 544368 97139 544370
rect 94638 544312 97078 544368
rect 97134 544312 97139 544368
rect 94638 544310 97139 544312
rect 97073 544307 97139 544310
rect 65793 544096 68938 544098
rect 65793 544040 65798 544096
rect 65854 544040 68938 544096
rect 65793 544038 68938 544040
rect 65793 544035 65859 544038
rect 67265 543418 67331 543421
rect 67950 543418 67956 543420
rect 67265 543416 67956 543418
rect 67265 543360 67270 543416
rect 67326 543360 67956 543416
rect 67265 543358 67956 543360
rect 67265 543355 67331 543358
rect 67950 543356 67956 543358
rect 68020 543418 68026 543420
rect 68020 543358 68938 543418
rect 68020 543356 68026 543358
rect 68878 543320 68938 543358
rect 94638 543010 94698 543592
rect 94773 543010 94839 543013
rect 94638 543008 94839 543010
rect 94638 542952 94778 543008
rect 94834 542952 94839 543008
rect 94638 542950 94839 542952
rect 94773 542947 94839 542950
rect 69246 541652 69306 541960
rect 69238 541588 69244 541652
rect 69308 541588 69314 541652
rect 94638 541650 94698 542232
rect 97165 541650 97231 541653
rect 94638 541648 97231 541650
rect 94638 541592 97170 541648
rect 97226 541592 97231 541648
rect 94638 541590 97231 541592
rect 14457 541106 14523 541109
rect 69246 541106 69306 541588
rect 97165 541587 97231 541590
rect 14457 541104 69306 541106
rect 14457 541048 14462 541104
rect 14518 541048 69306 541104
rect 14457 541046 69306 541048
rect 14457 541043 14523 541046
rect -960 540684 480 540924
rect 66437 540154 66503 540157
rect 68878 540154 68938 540600
rect 66437 540152 68938 540154
rect 66437 540096 66442 540152
rect 66498 540096 68938 540152
rect 66437 540094 68938 540096
rect 66437 540091 66503 540094
rect 94270 539749 94330 540872
rect 94270 539744 94379 539749
rect 94270 539688 94318 539744
rect 94374 539688 94379 539744
rect 94270 539686 94379 539688
rect 94313 539683 94379 539686
rect 75862 539548 75868 539612
rect 75932 539610 75938 539612
rect 76741 539610 76807 539613
rect 75932 539608 76807 539610
rect 75932 539552 76746 539608
rect 76802 539552 76807 539608
rect 75932 539550 76807 539552
rect 75932 539548 75938 539550
rect 76741 539547 76807 539550
rect 93945 538930 94011 538933
rect 94086 538930 94146 539512
rect 93945 538928 94146 538930
rect 93945 538872 93950 538928
rect 94006 538872 94146 538928
rect 93945 538870 94146 538872
rect 93945 538867 94011 538870
rect 583017 537842 583083 537845
rect 583520 537842 584960 537932
rect 583017 537840 584960 537842
rect 583017 537784 583022 537840
rect 583078 537784 584960 537840
rect 583017 537782 584960 537784
rect 583017 537779 583083 537782
rect 583520 537692 584960 537782
rect 60549 537434 60615 537437
rect 96838 537434 96844 537436
rect 60549 537432 96844 537434
rect 60549 537376 60554 537432
rect 60610 537376 96844 537432
rect 60549 537374 96844 537376
rect 60549 537371 60615 537374
rect 96838 537372 96844 537374
rect 96908 537372 96914 537436
rect 84009 536210 84075 536213
rect 104249 536210 104315 536213
rect 84009 536208 104315 536210
rect 84009 536152 84014 536208
rect 84070 536152 104254 536208
rect 104310 536152 104315 536208
rect 84009 536150 104315 536152
rect 84009 536147 84075 536150
rect 104249 536147 104315 536150
rect 80053 536074 80119 536077
rect 87597 536074 87663 536077
rect 80053 536072 87663 536074
rect 80053 536016 80058 536072
rect 80114 536016 87602 536072
rect 87658 536016 87663 536072
rect 80053 536014 87663 536016
rect 80053 536011 80119 536014
rect 87597 536011 87663 536014
rect 93393 536074 93459 536077
rect 136633 536074 136699 536077
rect 93393 536072 136699 536074
rect 93393 536016 93398 536072
rect 93454 536016 136638 536072
rect 136694 536016 136699 536072
rect 93393 536014 136699 536016
rect 93393 536011 93459 536014
rect 136633 536011 136699 536014
rect 68921 535530 68987 535533
rect 73797 535530 73863 535533
rect 68921 535528 73863 535530
rect 68921 535472 68926 535528
rect 68982 535472 73802 535528
rect 73858 535472 73863 535528
rect 68921 535470 73863 535472
rect 68921 535467 68987 535470
rect 73797 535467 73863 535470
rect 104433 535530 104499 535533
rect 105118 535530 105124 535532
rect 104433 535528 105124 535530
rect 104433 535472 104438 535528
rect 104494 535472 105124 535528
rect 104433 535470 105124 535472
rect 104433 535467 104499 535470
rect 105118 535468 105124 535470
rect 105188 535468 105194 535532
rect 79726 534652 79732 534716
rect 79796 534714 79802 534716
rect 95601 534714 95667 534717
rect 79796 534712 95667 534714
rect 79796 534656 95606 534712
rect 95662 534656 95667 534712
rect 79796 534654 95667 534656
rect 79796 534652 79802 534654
rect 95601 534651 95667 534654
rect -960 527914 480 528004
rect 3509 527914 3575 527917
rect -960 527912 3575 527914
rect -960 527856 3514 527912
rect 3570 527856 3575 527912
rect -960 527854 3575 527856
rect -960 527764 480 527854
rect 3509 527851 3575 527854
rect 582833 524514 582899 524517
rect 583520 524514 584960 524604
rect 582833 524512 584960 524514
rect 582833 524456 582838 524512
rect 582894 524456 584960 524512
rect 582833 524454 584960 524456
rect 582833 524451 582899 524454
rect 583520 524364 584960 524454
rect 72734 523636 72740 523700
rect 72804 523698 72810 523700
rect 95417 523698 95483 523701
rect 72804 523696 95483 523698
rect 72804 523640 95422 523696
rect 95478 523640 95483 523696
rect 72804 523638 95483 523640
rect 72804 523636 72810 523638
rect 95417 523635 95483 523638
rect 65977 522338 66043 522341
rect 114502 522338 114508 522340
rect 65977 522336 114508 522338
rect 65977 522280 65982 522336
rect 66038 522280 114508 522336
rect 65977 522278 114508 522280
rect 65977 522275 66043 522278
rect 114502 522276 114508 522278
rect 114572 522276 114578 522340
rect 69790 520916 69796 520980
rect 69860 520978 69866 520980
rect 88742 520978 88748 520980
rect 69860 520918 88748 520978
rect 69860 520916 69866 520918
rect 88742 520916 88748 520918
rect 88812 520916 88818 520980
rect -960 514858 480 514948
rect 3509 514858 3575 514861
rect -960 514856 3575 514858
rect -960 514800 3514 514856
rect 3570 514800 3575 514856
rect -960 514798 3575 514800
rect -960 514708 480 514798
rect 3509 514795 3575 514798
rect 583201 511322 583267 511325
rect 583520 511322 584960 511412
rect 583201 511320 584960 511322
rect 583201 511264 583206 511320
rect 583262 511264 584960 511320
rect 583201 511262 584960 511264
rect 583201 511259 583267 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3417 501802 3483 501805
rect -960 501800 3483 501802
rect -960 501744 3422 501800
rect 3478 501744 3483 501800
rect -960 501742 3483 501744
rect -960 501652 480 501742
rect 3417 501739 3483 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect 67766 482156 67772 482220
rect 67836 482218 67842 482220
rect 91318 482218 91324 482220
rect 67836 482158 91324 482218
rect 67836 482156 67842 482158
rect 91318 482156 91324 482158
rect 91388 482156 91394 482220
rect 73286 478076 73292 478140
rect 73356 478138 73362 478140
rect 92606 478138 92612 478140
rect 73356 478078 92612 478138
rect 73356 478076 73362 478078
rect 92606 478076 92612 478078
rect 92676 478076 92682 478140
rect 69606 476716 69612 476780
rect 69676 476778 69682 476780
rect 104198 476778 104204 476780
rect 69676 476718 104204 476778
rect 69676 476716 69682 476718
rect 104198 476716 104204 476718
rect 104268 476716 104274 476780
rect -960 475690 480 475780
rect 2773 475690 2839 475693
rect -960 475688 2839 475690
rect -960 475632 2778 475688
rect 2834 475632 2839 475688
rect -960 475630 2839 475632
rect -960 475540 480 475630
rect 2773 475627 2839 475630
rect 65977 475418 66043 475421
rect 75862 475418 75868 475420
rect 65977 475416 75868 475418
rect 65977 475360 65982 475416
rect 66038 475360 75868 475416
rect 65977 475358 75868 475360
rect 65977 475355 66043 475358
rect 75862 475356 75868 475358
rect 75932 475356 75938 475420
rect 67633 474058 67699 474061
rect 96838 474058 96844 474060
rect 67633 474056 96844 474058
rect 67633 474000 67638 474056
rect 67694 474000 96844 474056
rect 67633 473998 96844 474000
rect 67633 473995 67699 473998
rect 96838 473996 96844 473998
rect 96908 473996 96914 474060
rect 73153 472562 73219 472565
rect 111926 472562 111932 472564
rect 73153 472560 111932 472562
rect 73153 472504 73158 472560
rect 73214 472504 111932 472560
rect 73153 472502 111932 472504
rect 73153 472499 73219 472502
rect 111926 472500 111932 472502
rect 111996 472500 112002 472564
rect 67950 471820 67956 471884
rect 68020 471882 68026 471884
rect 68921 471882 68987 471885
rect 68020 471880 68987 471882
rect 68020 471824 68926 471880
rect 68982 471824 68987 471880
rect 68020 471822 68987 471824
rect 68020 471820 68026 471822
rect 68921 471819 68987 471822
rect 583109 471474 583175 471477
rect 583520 471474 584960 471564
rect 583109 471472 584960 471474
rect 583109 471416 583114 471472
rect 583170 471416 584960 471472
rect 583109 471414 584960 471416
rect 583109 471411 583175 471414
rect 583520 471324 584960 471414
rect 68921 470658 68987 470661
rect 208393 470658 208459 470661
rect 68921 470656 208459 470658
rect 68921 470600 68926 470656
rect 68982 470600 208398 470656
rect 208454 470600 208459 470656
rect 68921 470598 208459 470600
rect 68921 470595 68987 470598
rect 208393 470595 208459 470598
rect 67766 467876 67772 467940
rect 67836 467938 67842 467940
rect 70342 467938 70348 467940
rect 67836 467878 70348 467938
rect 67836 467876 67842 467878
rect 70342 467876 70348 467878
rect 70412 467876 70418 467940
rect 107009 467938 107075 467941
rect 107561 467938 107627 467941
rect 258073 467938 258139 467941
rect 107009 467936 258139 467938
rect 107009 467880 107014 467936
rect 107070 467880 107566 467936
rect 107622 467880 258078 467936
rect 258134 467880 258139 467936
rect 107009 467878 258139 467880
rect 107009 467875 107075 467878
rect 107561 467875 107627 467878
rect 258073 467875 258139 467878
rect 69657 465218 69723 465221
rect 194593 465218 194659 465221
rect 69657 465216 194659 465218
rect 69657 465160 69662 465216
rect 69718 465160 194598 465216
rect 194654 465160 194659 465216
rect 69657 465158 194659 465160
rect 69657 465155 69723 465158
rect 194593 465155 194659 465158
rect 213913 465218 213979 465221
rect 215201 465218 215267 465221
rect 269062 465218 269068 465220
rect 213913 465216 269068 465218
rect 213913 465160 213918 465216
rect 213974 465160 215206 465216
rect 215262 465160 269068 465216
rect 213913 465158 269068 465160
rect 213913 465155 213979 465158
rect 215201 465155 215267 465158
rect 269062 465156 269068 465158
rect 269132 465156 269138 465220
rect 215293 465082 215359 465085
rect 215937 465082 216003 465085
rect 215293 465080 216003 465082
rect 215293 465024 215298 465080
rect 215354 465024 215942 465080
rect 215998 465024 216003 465080
rect 215293 465022 216003 465024
rect 215293 465019 215359 465022
rect 215937 465019 216003 465022
rect 75678 464340 75684 464404
rect 75748 464402 75754 464404
rect 92381 464402 92447 464405
rect 75748 464400 92447 464402
rect 75748 464344 92386 464400
rect 92442 464344 92447 464400
rect 75748 464342 92447 464344
rect 75748 464340 75754 464342
rect 92381 464339 92447 464342
rect 184197 463722 184263 463725
rect 215293 463722 215359 463725
rect 184197 463720 215359 463722
rect 184197 463664 184202 463720
rect 184258 463664 215298 463720
rect 215354 463664 215359 463720
rect 184197 463662 215359 463664
rect 184197 463659 184263 463662
rect 215293 463659 215359 463662
rect 123477 462906 123543 462909
rect 258574 462906 258580 462908
rect 123477 462904 258580 462906
rect 123477 462848 123482 462904
rect 123538 462848 258580 462904
rect 123477 462846 258580 462848
rect 123477 462843 123543 462846
rect 258574 462844 258580 462846
rect 258644 462844 258650 462908
rect -960 462634 480 462724
rect 3509 462634 3575 462637
rect -960 462632 3575 462634
rect -960 462576 3514 462632
rect 3570 462576 3575 462632
rect -960 462574 3575 462576
rect -960 462484 480 462574
rect 3509 462571 3575 462574
rect 212533 462226 212599 462229
rect 213177 462226 213243 462229
rect 212533 462224 213243 462226
rect 212533 462168 212538 462224
rect 212594 462168 213182 462224
rect 213238 462168 213243 462224
rect 212533 462166 213243 462168
rect 212533 462163 212599 462166
rect 213177 462163 213243 462166
rect 180057 461138 180123 461141
rect 212533 461138 212599 461141
rect 180057 461136 212599 461138
rect 180057 461080 180062 461136
rect 180118 461080 212538 461136
rect 212594 461080 212599 461136
rect 180057 461078 212599 461080
rect 180057 461075 180123 461078
rect 212533 461075 212599 461078
rect 133137 461002 133203 461005
rect 260925 461002 260991 461005
rect 133137 461000 260991 461002
rect 133137 460944 133142 461000
rect 133198 460944 260930 461000
rect 260986 460944 260991 461000
rect 133137 460942 260991 460944
rect 133137 460939 133203 460942
rect 260925 460939 260991 460942
rect 71773 460186 71839 460189
rect 114318 460186 114324 460188
rect 71773 460184 114324 460186
rect 71773 460128 71778 460184
rect 71834 460128 114324 460184
rect 71773 460126 114324 460128
rect 71773 460123 71839 460126
rect 114318 460124 114324 460126
rect 114388 460124 114394 460188
rect 101990 459580 101996 459644
rect 102060 459642 102066 459644
rect 254117 459642 254183 459645
rect 102060 459640 254183 459642
rect 102060 459584 254122 459640
rect 254178 459584 254183 459640
rect 102060 459582 254183 459584
rect 102060 459580 102066 459582
rect 254117 459579 254183 459582
rect 582649 458826 582715 458829
rect 287010 458824 582715 458826
rect 287010 458768 582654 458824
rect 582710 458768 582715 458824
rect 287010 458766 582715 458768
rect 216673 458690 216739 458693
rect 220077 458690 220143 458693
rect 216673 458688 220143 458690
rect 216673 458632 216678 458688
rect 216734 458632 220082 458688
rect 220138 458632 220143 458688
rect 216673 458630 220143 458632
rect 216673 458627 216739 458630
rect 220077 458627 220143 458630
rect 115289 458554 115355 458557
rect 253054 458554 253060 458556
rect 115289 458552 253060 458554
rect 115289 458496 115294 458552
rect 115350 458496 253060 458552
rect 115289 458494 253060 458496
rect 115289 458491 115355 458494
rect 253054 458492 253060 458494
rect 253124 458492 253130 458556
rect 185669 458418 185735 458421
rect 216673 458418 216739 458421
rect 185669 458416 216739 458418
rect 185669 458360 185674 458416
rect 185730 458360 216678 458416
rect 216734 458360 216739 458416
rect 185669 458358 216739 458360
rect 185669 458355 185735 458358
rect 216673 458355 216739 458358
rect 220813 458418 220879 458421
rect 284385 458418 284451 458421
rect 287010 458418 287070 458766
rect 582649 458763 582715 458766
rect 220813 458416 287070 458418
rect 220813 458360 220818 458416
rect 220874 458360 284390 458416
rect 284446 458360 287070 458416
rect 220813 458358 287070 458360
rect 220813 458355 220879 458358
rect 284385 458355 284451 458358
rect 197077 458284 197143 458285
rect 197077 458280 197124 458284
rect 197188 458282 197194 458284
rect 197077 458224 197082 458280
rect 197077 458220 197124 458224
rect 197188 458222 197234 458282
rect 197188 458220 197194 458222
rect 197077 458219 197143 458220
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect 175181 457058 175247 457061
rect 207473 457058 207539 457061
rect 175181 457056 207539 457058
rect 175181 457000 175186 457056
rect 175242 457000 207478 457056
rect 207534 457000 207539 457056
rect 175181 456998 207539 457000
rect 175181 456995 175247 456998
rect 207473 456995 207539 456998
rect 183461 456922 183527 456925
rect 215385 456922 215451 456925
rect 183461 456920 215451 456922
rect 183461 456864 183466 456920
rect 183522 456864 215390 456920
rect 215446 456864 215451 456920
rect 183461 456862 215451 456864
rect 183461 456859 183527 456862
rect 215385 456859 215451 456862
rect 230473 456922 230539 456925
rect 231117 456922 231183 456925
rect 287053 456922 287119 456925
rect 288341 456922 288407 456925
rect 230473 456920 288407 456922
rect 230473 456864 230478 456920
rect 230534 456864 231122 456920
rect 231178 456864 287058 456920
rect 287114 456864 288346 456920
rect 288402 456864 288407 456920
rect 230473 456862 288407 456864
rect 230473 456859 230539 456862
rect 231117 456859 231183 456862
rect 287053 456859 287119 456862
rect 288341 456859 288407 456862
rect 96613 456108 96679 456109
rect 80646 456044 80652 456108
rect 80716 456106 80722 456108
rect 96613 456106 96660 456108
rect 80716 456046 84210 456106
rect 96568 456104 96660 456106
rect 96568 456048 96618 456104
rect 96568 456046 96660 456048
rect 80716 456044 80722 456046
rect 84150 455970 84210 456046
rect 96613 456044 96660 456046
rect 96724 456044 96730 456108
rect 96613 456043 96679 456044
rect 96654 455970 96660 455972
rect 84150 455910 96660 455970
rect 96654 455908 96660 455910
rect 96724 455908 96730 455972
rect 180149 455834 180215 455837
rect 219801 455834 219867 455837
rect 180149 455832 219867 455834
rect 180149 455776 180154 455832
rect 180210 455776 219806 455832
rect 219862 455776 219867 455832
rect 180149 455774 219867 455776
rect 180149 455771 180215 455774
rect 219801 455771 219867 455774
rect 78029 455698 78095 455701
rect 202873 455698 202939 455701
rect 78029 455696 202939 455698
rect 78029 455640 78034 455696
rect 78090 455640 202878 455696
rect 202934 455640 202939 455696
rect 78029 455638 202939 455640
rect 78029 455635 78095 455638
rect 202873 455635 202939 455638
rect 224953 455698 225019 455701
rect 267774 455698 267780 455700
rect 224953 455696 267780 455698
rect 224953 455640 224958 455696
rect 225014 455640 267780 455696
rect 224953 455638 267780 455640
rect 224953 455635 225019 455638
rect 267774 455636 267780 455638
rect 267844 455636 267850 455700
rect 119429 455562 119495 455565
rect 255313 455562 255379 455565
rect 119429 455560 255379 455562
rect 119429 455504 119434 455560
rect 119490 455504 255318 455560
rect 255374 455504 255379 455560
rect 119429 455502 255379 455504
rect 119429 455499 119495 455502
rect 255313 455499 255379 455502
rect 242157 455426 242223 455429
rect 243537 455426 243603 455429
rect 242157 455424 243603 455426
rect 242157 455368 242162 455424
rect 242218 455368 243542 455424
rect 243598 455368 243603 455424
rect 242157 455366 243603 455368
rect 242157 455363 242223 455366
rect 243537 455363 243603 455366
rect 191281 454338 191347 454341
rect 222561 454338 222627 454341
rect 191281 454336 222627 454338
rect 191281 454280 191286 454336
rect 191342 454280 222566 454336
rect 222622 454280 222627 454336
rect 191281 454278 222627 454280
rect 191281 454275 191347 454278
rect 222561 454275 222627 454278
rect 147581 454202 147647 454205
rect 197905 454202 197971 454205
rect 147581 454200 197971 454202
rect 147581 454144 147586 454200
rect 147642 454144 197910 454200
rect 197966 454144 197971 454200
rect 147581 454142 197971 454144
rect 147581 454139 147647 454142
rect 197905 454139 197971 454142
rect 243537 454202 243603 454205
rect 266486 454202 266492 454204
rect 243537 454200 266492 454202
rect 243537 454144 243542 454200
rect 243598 454144 266492 454200
rect 243537 454142 266492 454144
rect 243537 454139 243603 454142
rect 266486 454140 266492 454142
rect 266556 454140 266562 454204
rect 178677 454066 178743 454069
rect 255957 454066 256023 454069
rect 178677 454064 256023 454066
rect 178677 454008 178682 454064
rect 178738 454008 255962 454064
rect 256018 454008 256023 454064
rect 178677 454006 256023 454008
rect 178677 454003 178743 454006
rect 255957 454003 256023 454006
rect 44081 453250 44147 453253
rect 85757 453250 85823 453253
rect 44081 453248 85823 453250
rect 44081 453192 44086 453248
rect 44142 453192 85762 453248
rect 85818 453192 85823 453248
rect 44081 453190 85823 453192
rect 44081 453187 44147 453190
rect 85757 453187 85823 453190
rect 166257 453114 166323 453117
rect 194542 453114 194548 453116
rect 166257 453112 194548 453114
rect 166257 453056 166262 453112
rect 166318 453056 194548 453112
rect 166257 453054 194548 453056
rect 166257 453051 166323 453054
rect 194542 453052 194548 453054
rect 194612 453052 194618 453116
rect 225965 453114 226031 453117
rect 288433 453114 288499 453117
rect 225965 453112 288499 453114
rect 225965 453056 225970 453112
rect 226026 453056 288438 453112
rect 288494 453056 288499 453112
rect 225965 453054 288499 453056
rect 225965 453051 226031 453054
rect 288433 453051 288499 453054
rect 188061 452978 188127 452981
rect 202137 452978 202203 452981
rect 188061 452976 202203 452978
rect 188061 452920 188066 452976
rect 188122 452920 202142 452976
rect 202198 452920 202203 452976
rect 188061 452918 202203 452920
rect 188061 452915 188127 452918
rect 202137 452915 202203 452918
rect 222101 452978 222167 452981
rect 241646 452978 241652 452980
rect 222101 452976 241652 452978
rect 222101 452920 222106 452976
rect 222162 452920 241652 452976
rect 222101 452918 241652 452920
rect 222101 452915 222167 452918
rect 241646 452916 241652 452918
rect 241716 452916 241722 452980
rect 246021 452978 246087 452981
rect 251541 452978 251607 452981
rect 246021 452976 251607 452978
rect 246021 452920 246026 452976
rect 246082 452920 251546 452976
rect 251602 452920 251607 452976
rect 246021 452918 251607 452920
rect 246021 452915 246087 452918
rect 251541 452915 251607 452918
rect 189717 452842 189783 452845
rect 210693 452842 210759 452845
rect 189717 452840 210759 452842
rect 189717 452784 189722 452840
rect 189778 452784 210698 452840
rect 210754 452784 210759 452840
rect 189717 452782 210759 452784
rect 189717 452779 189783 452782
rect 210693 452779 210759 452782
rect 225597 452842 225663 452845
rect 228725 452842 228791 452845
rect 253841 452842 253907 452845
rect 225597 452840 253907 452842
rect 225597 452784 225602 452840
rect 225658 452784 228730 452840
rect 228786 452784 253846 452840
rect 253902 452784 253907 452840
rect 225597 452782 253907 452784
rect 225597 452779 225663 452782
rect 228725 452779 228791 452782
rect 253841 452779 253907 452782
rect 252461 452706 252527 452709
rect 258165 452706 258231 452709
rect 252461 452704 258231 452706
rect 252461 452648 252466 452704
rect 252522 452648 258170 452704
rect 258226 452648 258231 452704
rect 252461 452646 258231 452648
rect 252461 452643 252527 452646
rect 258165 452643 258231 452646
rect 142061 451890 142127 451893
rect 204437 451890 204503 451893
rect 142061 451888 204503 451890
rect 142061 451832 142066 451888
rect 142122 451832 204442 451888
rect 204498 451832 204503 451888
rect 142061 451830 204503 451832
rect 142061 451827 142127 451830
rect 204437 451827 204503 451830
rect 235349 451618 235415 451621
rect 247718 451618 247724 451620
rect 235349 451616 247724 451618
rect 235349 451560 235354 451616
rect 235410 451560 247724 451616
rect 235349 451558 247724 451560
rect 235349 451555 235415 451558
rect 247718 451556 247724 451558
rect 247788 451556 247794 451620
rect 193305 451482 193371 451485
rect 207013 451482 207079 451485
rect 193305 451480 207079 451482
rect 193305 451424 193310 451480
rect 193366 451424 207018 451480
rect 207074 451424 207079 451480
rect 193305 451422 207079 451424
rect 193305 451419 193371 451422
rect 207013 451419 207079 451422
rect 210693 451482 210759 451485
rect 210693 451480 277410 451482
rect 210693 451424 210698 451480
rect 210754 451424 277410 451480
rect 210693 451422 277410 451424
rect 210693 451419 210759 451422
rect 116761 451346 116827 451349
rect 249701 451346 249767 451349
rect 254669 451346 254735 451349
rect 116761 451344 254735 451346
rect 116761 451288 116766 451344
rect 116822 451288 249706 451344
rect 249762 451288 254674 451344
rect 254730 451288 254735 451344
rect 116761 451286 254735 451288
rect 277350 451346 277410 451422
rect 287145 451346 287211 451349
rect 583201 451346 583267 451349
rect 277350 451344 583267 451346
rect 277350 451288 287150 451344
rect 287206 451288 583206 451344
rect 583262 451288 583267 451344
rect 277350 451286 583267 451288
rect 116761 451283 116827 451286
rect 249701 451283 249767 451286
rect 254669 451283 254735 451286
rect 287145 451283 287211 451286
rect 583201 451283 583267 451286
rect 193806 450332 193812 450396
rect 193876 450394 193882 450396
rect 201585 450394 201651 450397
rect 193876 450392 201651 450394
rect 193876 450336 201590 450392
rect 201646 450336 201651 450392
rect 193876 450334 201651 450336
rect 193876 450332 193882 450334
rect 201585 450331 201651 450334
rect 194593 450260 194659 450261
rect 194542 450196 194548 450260
rect 194612 450258 194659 450260
rect 228081 450258 228147 450261
rect 263593 450258 263659 450261
rect 194612 450256 194704 450258
rect 194654 450200 194704 450256
rect 194612 450198 194704 450200
rect 228081 450256 263659 450258
rect 228081 450200 228086 450256
rect 228142 450200 263598 450256
rect 263654 450200 263659 450256
rect 228081 450198 263659 450200
rect 194612 450196 194659 450198
rect 194593 450195 194659 450196
rect 228081 450195 228147 450198
rect 263593 450195 263659 450198
rect 187049 450122 187115 450125
rect 233141 450122 233207 450125
rect 187049 450120 233207 450122
rect 187049 450064 187054 450120
rect 187110 450064 233146 450120
rect 233202 450064 233207 450120
rect 187049 450062 233207 450064
rect 187049 450059 187115 450062
rect 233141 450059 233207 450062
rect 242433 450122 242499 450125
rect 256734 450122 256740 450124
rect 242433 450120 256740 450122
rect 242433 450064 242438 450120
rect 242494 450064 256740 450120
rect 242433 450062 256740 450064
rect 242433 450059 242499 450062
rect 256734 450060 256740 450062
rect 256804 450060 256810 450124
rect 92565 449986 92631 449989
rect 220813 449986 220879 449989
rect 92565 449984 220879 449986
rect 92565 449928 92570 449984
rect 92626 449928 220818 449984
rect 220874 449928 220879 449984
rect 92565 449926 220879 449928
rect 92565 449923 92631 449926
rect 220813 449923 220879 449926
rect 237649 449986 237715 449989
rect 244406 449986 244412 449988
rect 237649 449984 244412 449986
rect 237649 449928 237654 449984
rect 237710 449928 244412 449984
rect 237649 449926 244412 449928
rect 237649 449923 237715 449926
rect 244406 449924 244412 449926
rect 244476 449924 244482 449988
rect 249742 449924 249748 449988
rect 249812 449986 249818 449988
rect 250253 449986 250319 449989
rect 249812 449984 250319 449986
rect 249812 449928 250258 449984
rect 250314 449928 250319 449984
rect 249812 449926 250319 449928
rect 249812 449924 249818 449926
rect 250253 449923 250319 449926
rect 193489 449716 193555 449717
rect 242985 449716 243051 449717
rect 193438 449714 193444 449716
rect -960 449578 480 449668
rect 193398 449654 193444 449714
rect 193508 449712 193555 449716
rect 242934 449714 242940 449716
rect 193550 449656 193555 449712
rect 193438 449652 193444 449654
rect 193508 449652 193555 449656
rect 242894 449654 242940 449714
rect 243004 449712 243051 449716
rect 243046 449656 243051 449712
rect 242934 449652 242940 449654
rect 243004 449652 243051 449656
rect 193489 449651 193555 449652
rect 242985 449651 243051 449652
rect 3141 449578 3207 449581
rect -960 449576 3207 449578
rect -960 449520 3146 449576
rect 3202 449520 3207 449576
rect -960 449518 3207 449520
rect -960 449428 480 449518
rect 3141 449515 3207 449518
rect 111057 449170 111123 449173
rect 191465 449170 191531 449173
rect 111057 449168 191531 449170
rect 111057 449112 111062 449168
rect 111118 449112 191470 449168
rect 191526 449112 191531 449168
rect 111057 449110 191531 449112
rect 111057 449107 111123 449110
rect 191465 449107 191531 449110
rect 191649 449170 191715 449173
rect 191649 449168 193660 449170
rect 191649 449112 191654 449168
rect 191710 449112 193660 449168
rect 191649 449110 193660 449112
rect 191649 449107 191715 449110
rect 255957 448898 256023 448901
rect 253460 448896 256023 448898
rect 253460 448840 255962 448896
rect 256018 448840 256023 448896
rect 253460 448838 256023 448840
rect 255957 448835 256023 448838
rect 110413 448626 110479 448629
rect 111057 448626 111123 448629
rect 110413 448624 111123 448626
rect 110413 448568 110418 448624
rect 110474 448568 111062 448624
rect 111118 448568 111123 448624
rect 110413 448566 111123 448568
rect 110413 448563 110479 448566
rect 111057 448563 111123 448566
rect 181529 447946 181595 447949
rect 193305 447946 193371 447949
rect 181529 447944 193371 447946
rect 181529 447888 181534 447944
rect 181590 447888 193310 447944
rect 193366 447888 193371 447944
rect 181529 447886 193371 447888
rect 181529 447883 181595 447886
rect 193305 447883 193371 447886
rect 190453 447266 190519 447269
rect 193630 447266 193690 447780
rect 254117 447538 254183 447541
rect 254577 447538 254643 447541
rect 253460 447536 254643 447538
rect 253460 447480 254122 447536
rect 254178 447480 254582 447536
rect 254638 447480 254643 447536
rect 253460 447478 254643 447480
rect 254117 447475 254183 447478
rect 254577 447475 254643 447478
rect 190453 447264 193690 447266
rect 190453 447208 190458 447264
rect 190514 447208 193690 447264
rect 190453 447206 193690 447208
rect 190453 447203 190519 447206
rect 95141 446450 95207 446453
rect 96470 446450 96476 446452
rect 95141 446448 96476 446450
rect 95141 446392 95146 446448
rect 95202 446392 96476 446448
rect 95141 446390 96476 446392
rect 95141 446387 95207 446390
rect 96470 446388 96476 446390
rect 96540 446450 96546 446452
rect 191189 446450 191255 446453
rect 96540 446448 191255 446450
rect 96540 446392 191194 446448
rect 191250 446392 191255 446448
rect 96540 446390 191255 446392
rect 96540 446388 96546 446390
rect 191189 446387 191255 446390
rect 191741 446450 191807 446453
rect 191741 446448 193660 446450
rect 191741 446392 191746 446448
rect 191802 446392 193660 446448
rect 191741 446390 193660 446392
rect 191741 446387 191807 446390
rect 255681 446178 255747 446181
rect 256049 446178 256115 446181
rect 253460 446176 256115 446178
rect 253460 446120 255686 446176
rect 255742 446120 256054 446176
rect 256110 446120 256115 446176
rect 253460 446118 256115 446120
rect 255681 446115 255747 446118
rect 256049 446115 256115 446118
rect 191741 445090 191807 445093
rect 191741 445088 193660 445090
rect 191741 445032 191746 445088
rect 191802 445032 193660 445088
rect 191741 445030 193660 445032
rect 191741 445027 191807 445030
rect 75361 444954 75427 444957
rect 188061 444954 188127 444957
rect 75361 444952 188127 444954
rect 75361 444896 75366 444952
rect 75422 444896 188066 444952
rect 188122 444896 188127 444952
rect 75361 444894 188127 444896
rect 75361 444891 75427 444894
rect 188061 444891 188127 444894
rect 255313 444818 255379 444821
rect 253460 444816 255379 444818
rect 253460 444760 255318 444816
rect 255374 444760 255379 444816
rect 253460 444758 255379 444760
rect 255313 444755 255379 444758
rect 583520 444668 584960 444908
rect 66069 443050 66135 443053
rect 70485 443050 70551 443053
rect 66069 443048 70551 443050
rect 66069 442992 66074 443048
rect 66130 442992 70490 443048
rect 70546 442992 70551 443048
rect 66069 442990 70551 442992
rect 66069 442987 66135 442990
rect 70485 442987 70551 442990
rect 71129 443050 71195 443053
rect 169661 443050 169727 443053
rect 193630 443050 193690 443700
rect 255405 443458 255471 443461
rect 253460 443456 255471 443458
rect 253460 443400 255410 443456
rect 255466 443400 255471 443456
rect 253460 443398 255471 443400
rect 255405 443395 255471 443398
rect 71129 443048 193690 443050
rect 71129 442992 71134 443048
rect 71190 442992 169666 443048
rect 169722 442992 193690 443048
rect 71129 442990 193690 442992
rect 71129 442987 71195 442990
rect 169661 442987 169727 442990
rect 71681 442914 71747 442917
rect 193438 442914 193444 442916
rect 71681 442912 193444 442914
rect 71681 442856 71686 442912
rect 71742 442856 193444 442912
rect 71681 442854 193444 442856
rect 71681 442851 71747 442854
rect 193438 442852 193444 442854
rect 193508 442852 193514 442916
rect 193121 442098 193187 442101
rect 255129 442098 255195 442101
rect 258390 442098 258396 442100
rect 193121 442096 193660 442098
rect 193121 442040 193126 442096
rect 193182 442040 193660 442096
rect 193121 442038 193660 442040
rect 253460 442096 258396 442098
rect 253460 442040 255134 442096
rect 255190 442040 258396 442096
rect 253460 442038 258396 442040
rect 193121 442035 193187 442038
rect 255129 442035 255195 442038
rect 258390 442036 258396 442038
rect 258460 442036 258466 442100
rect 95325 440874 95391 440877
rect 107694 440874 107700 440876
rect 95325 440872 107700 440874
rect 95325 440816 95330 440872
rect 95386 440816 107700 440872
rect 95325 440814 107700 440816
rect 95325 440811 95391 440814
rect 107694 440812 107700 440814
rect 107764 440812 107770 440876
rect 192702 440676 192708 440740
rect 192772 440738 192778 440740
rect 192772 440678 193660 440738
rect 192772 440676 192778 440678
rect 253933 440466 253999 440469
rect 252908 440464 253999 440466
rect 252908 440436 253938 440464
rect 252878 440408 253938 440436
rect 253994 440408 253999 440464
rect 252878 440406 253999 440408
rect 67950 440268 67956 440332
rect 68020 440330 68026 440332
rect 69013 440330 69079 440333
rect 68020 440328 69079 440330
rect 68020 440272 69018 440328
rect 69074 440272 69079 440328
rect 68020 440270 69079 440272
rect 68020 440268 68026 440270
rect 69013 440267 69079 440270
rect 88517 440330 88583 440333
rect 120165 440330 120231 440333
rect 252878 440332 252938 440406
rect 253933 440403 253999 440406
rect 88517 440328 120231 440330
rect 88517 440272 88522 440328
rect 88578 440272 120170 440328
rect 120226 440272 120231 440328
rect 88517 440270 120231 440272
rect 88517 440267 88583 440270
rect 120165 440267 120231 440270
rect 252870 440268 252876 440332
rect 252940 440268 252946 440332
rect 61745 439514 61811 439517
rect 75913 439514 75979 439517
rect 82905 439514 82971 439517
rect 61745 439512 82971 439514
rect 61745 439456 61750 439512
rect 61806 439456 75918 439512
rect 75974 439456 82910 439512
rect 82966 439456 82971 439512
rect 61745 439454 82971 439456
rect 61745 439451 61811 439454
rect 75913 439451 75979 439454
rect 82905 439451 82971 439454
rect 69422 438908 69428 438972
rect 69492 438970 69498 438972
rect 193630 438970 193690 439348
rect 255405 439106 255471 439109
rect 253460 439104 255471 439106
rect 253460 439048 255410 439104
rect 255466 439048 255471 439104
rect 253460 439046 255471 439048
rect 255405 439043 255471 439046
rect 69492 438910 193690 438970
rect 69492 438908 69498 438910
rect 88926 438772 88932 438836
rect 88996 438834 89002 438836
rect 189717 438834 189783 438837
rect 88996 438832 189783 438834
rect 88996 438776 189722 438832
rect 189778 438776 189783 438832
rect 88996 438774 189783 438776
rect 88996 438772 89002 438774
rect 189717 438771 189783 438774
rect 81341 438290 81407 438293
rect 88926 438290 88932 438292
rect 81341 438288 88932 438290
rect 81341 438232 81346 438288
rect 81402 438232 88932 438288
rect 81341 438230 88932 438232
rect 81341 438227 81407 438230
rect 88926 438228 88932 438230
rect 88996 438228 89002 438292
rect 62757 438154 62823 438157
rect 65793 438154 65859 438157
rect 82813 438154 82879 438157
rect 62757 438152 82879 438154
rect 62757 438096 62762 438152
rect 62818 438096 65798 438152
rect 65854 438096 82818 438152
rect 82874 438096 82879 438152
rect 62757 438094 82879 438096
rect 62757 438091 62823 438094
rect 65793 438091 65859 438094
rect 82813 438091 82879 438094
rect 101990 438092 101996 438156
rect 102060 438154 102066 438156
rect 112110 438154 112116 438156
rect 102060 438094 112116 438154
rect 102060 438092 102066 438094
rect 112110 438092 112116 438094
rect 112180 438092 112186 438156
rect 191741 438018 191807 438021
rect 191741 438016 193660 438018
rect 191741 437960 191746 438016
rect 191802 437960 193660 438016
rect 191741 437958 193660 437960
rect 191741 437955 191807 437958
rect 255497 437746 255563 437749
rect 253460 437744 255563 437746
rect 253460 437688 255502 437744
rect 255558 437688 255563 437744
rect 253460 437686 255563 437688
rect 255497 437683 255563 437686
rect 82118 437412 82124 437476
rect 82188 437474 82194 437476
rect 83958 437474 83964 437476
rect 82188 437414 83964 437474
rect 82188 437412 82194 437414
rect 83958 437412 83964 437414
rect 84028 437412 84034 437476
rect 187049 437474 187115 437477
rect 122790 437472 187115 437474
rect 122790 437416 187054 437472
rect 187110 437416 187115 437472
rect 122790 437414 187115 437416
rect 109677 437338 109743 437341
rect 116761 437338 116827 437341
rect 109677 437336 116827 437338
rect 109677 437280 109682 437336
rect 109738 437280 116766 437336
rect 116822 437280 116827 437336
rect 109677 437278 116827 437280
rect 109677 437275 109743 437278
rect 116761 437275 116827 437278
rect 68921 437202 68987 437205
rect 71589 437202 71655 437205
rect 122790 437202 122850 437414
rect 187049 437411 187115 437414
rect 68921 437200 71655 437202
rect 68921 437144 68926 437200
rect 68982 437144 71594 437200
rect 71650 437144 71655 437200
rect 68921 437142 71655 437144
rect 68921 437139 68987 437142
rect 71589 437139 71655 437142
rect 113130 437142 122850 437202
rect 106641 437066 106707 437069
rect 113130 437066 113190 437142
rect 106641 437064 113190 437066
rect 106641 437008 106646 437064
rect 106702 437008 113190 437064
rect 106641 437006 113190 437008
rect 106641 437003 106707 437006
rect 113265 436796 113331 436797
rect 113214 436794 113220 436796
rect -960 436508 480 436748
rect 113174 436734 113220 436794
rect 113284 436792 113331 436796
rect 113326 436736 113331 436792
rect 113214 436732 113220 436734
rect 113284 436732 113331 436736
rect 253054 436732 253060 436796
rect 253124 436794 253130 436796
rect 255221 436794 255287 436797
rect 255497 436794 255563 436797
rect 253124 436792 255563 436794
rect 253124 436736 255226 436792
rect 255282 436736 255502 436792
rect 255558 436736 255563 436792
rect 253124 436734 255563 436736
rect 253124 436732 253130 436734
rect 113265 436731 113331 436732
rect 192937 436658 193003 436661
rect 192937 436656 193660 436658
rect 192937 436600 192942 436656
rect 192998 436600 193660 436656
rect 192937 436598 193660 436600
rect 192937 436595 193003 436598
rect 94998 436460 95004 436524
rect 95068 436522 95074 436524
rect 99373 436522 99439 436525
rect 99741 436522 99807 436525
rect 95068 436520 99807 436522
rect 95068 436464 99378 436520
rect 99434 436464 99746 436520
rect 99802 436464 99807 436520
rect 95068 436462 99807 436464
rect 95068 436460 95074 436462
rect 99373 436459 99439 436462
rect 99741 436459 99807 436462
rect 96286 436324 96292 436388
rect 96356 436386 96362 436388
rect 101213 436386 101279 436389
rect 96356 436384 101279 436386
rect 96356 436328 101218 436384
rect 101274 436328 101279 436384
rect 253062 436356 253122 436732
rect 255221 436731 255287 436734
rect 255497 436731 255563 436734
rect 96356 436326 101279 436328
rect 96356 436324 96362 436326
rect 101213 436323 101279 436326
rect 68553 436250 68619 436253
rect 68553 436248 70410 436250
rect 68553 436192 68558 436248
rect 68614 436192 70410 436248
rect 68553 436190 70410 436192
rect 68553 436187 68619 436190
rect 61837 436114 61903 436117
rect 68921 436114 68987 436117
rect 61837 436112 68987 436114
rect 61837 436056 61842 436112
rect 61898 436056 68926 436112
rect 68982 436056 68987 436112
rect 61837 436054 68987 436056
rect 70350 436114 70410 436190
rect 73654 436188 73660 436252
rect 73724 436250 73730 436252
rect 80329 436250 80395 436253
rect 73724 436248 80395 436250
rect 73724 436192 80334 436248
rect 80390 436192 80395 436248
rect 73724 436190 80395 436192
rect 73724 436188 73730 436190
rect 80329 436187 80395 436190
rect 83958 436188 83964 436252
rect 84028 436250 84034 436252
rect 89713 436250 89779 436253
rect 84028 436248 89779 436250
rect 84028 436192 89718 436248
rect 89774 436192 89779 436248
rect 84028 436190 89779 436192
rect 84028 436188 84034 436190
rect 89713 436187 89779 436190
rect 71865 436114 71931 436117
rect 72693 436114 72759 436117
rect 70350 436112 72759 436114
rect 70350 436056 71870 436112
rect 71926 436056 72698 436112
rect 72754 436056 72759 436112
rect 70350 436054 72759 436056
rect 61837 436051 61903 436054
rect 68921 436051 68987 436054
rect 71865 436051 71931 436054
rect 72693 436051 72759 436054
rect 102726 436052 102732 436116
rect 102796 436114 102802 436116
rect 107653 436114 107719 436117
rect 108389 436114 108455 436117
rect 102796 436112 108455 436114
rect 102796 436056 107658 436112
rect 107714 436056 108394 436112
rect 108450 436056 108455 436112
rect 102796 436054 108455 436056
rect 102796 436052 102802 436054
rect 107653 436051 107719 436054
rect 108389 436051 108455 436054
rect 85849 435298 85915 435301
rect 86861 435298 86927 435301
rect 85849 435296 86927 435298
rect 85849 435240 85854 435296
rect 85910 435240 86866 435296
rect 86922 435240 86927 435296
rect 85849 435238 86927 435240
rect 85849 435235 85915 435238
rect 86861 435235 86927 435238
rect 191741 435298 191807 435301
rect 191741 435296 193660 435298
rect 191741 435240 191746 435296
rect 191802 435240 193660 435296
rect 191741 435238 193660 435240
rect 191741 435235 191807 435238
rect 72601 435026 72667 435029
rect 255405 435026 255471 435029
rect 72601 435024 84946 435026
rect 72601 434968 72606 435024
rect 72662 434968 84946 435024
rect 72601 434966 84946 434968
rect 253460 435024 255471 435026
rect 253460 434968 255410 435024
rect 255466 434968 255471 435024
rect 253460 434966 255471 434968
rect 72601 434963 72667 434966
rect 45461 434890 45527 434893
rect 81341 434890 81407 434893
rect 45461 434888 81407 434890
rect 45461 434832 45466 434888
rect 45522 434832 81346 434888
rect 81402 434832 81407 434888
rect 45461 434830 81407 434832
rect 45461 434827 45527 434830
rect 81341 434827 81407 434830
rect 84886 434754 84946 434966
rect 255405 434963 255471 434966
rect 86861 434890 86927 434893
rect 118734 434890 118740 434892
rect 86861 434888 118740 434890
rect 86861 434832 86866 434888
rect 86922 434832 118740 434888
rect 86861 434830 118740 434832
rect 86861 434827 86927 434830
rect 118734 434828 118740 434830
rect 118804 434828 118810 434892
rect 132493 434754 132559 434757
rect 84886 434752 132559 434754
rect 84886 434696 132498 434752
rect 132554 434696 132559 434752
rect 84886 434694 132559 434696
rect 132493 434691 132559 434694
rect 70158 434556 70164 434620
rect 70228 434618 70234 434620
rect 75637 434618 75703 434621
rect 70228 434616 75703 434618
rect 70228 434560 75642 434616
rect 75698 434560 75703 434616
rect 70228 434558 75703 434560
rect 70228 434556 70234 434558
rect 75637 434555 75703 434558
rect 92473 434618 92539 434621
rect 92974 434618 92980 434620
rect 92473 434616 92980 434618
rect 92473 434560 92478 434616
rect 92534 434560 92980 434616
rect 92473 434558 92980 434560
rect 92473 434555 92539 434558
rect 92974 434556 92980 434558
rect 93044 434556 93050 434620
rect 71630 434420 71636 434484
rect 71700 434482 71706 434484
rect 72509 434482 72575 434485
rect 71700 434480 72575 434482
rect 71700 434424 72514 434480
rect 72570 434424 72575 434480
rect 71700 434422 72575 434424
rect 71700 434420 71706 434422
rect 72509 434419 72575 434422
rect 72550 433740 72556 433804
rect 72620 433802 72626 433804
rect 79869 433802 79935 433805
rect 72620 433800 79935 433802
rect 72620 433744 79874 433800
rect 79930 433744 79935 433800
rect 72620 433742 79935 433744
rect 72620 433740 72626 433742
rect 79869 433739 79935 433742
rect 90214 433740 90220 433804
rect 90284 433802 90290 433804
rect 91461 433802 91527 433805
rect 90284 433800 91527 433802
rect 90284 433744 91466 433800
rect 91522 433744 91527 433800
rect 90284 433742 91527 433744
rect 90284 433740 90290 433742
rect 91461 433739 91527 433742
rect 94446 433740 94452 433804
rect 94516 433802 94522 433804
rect 96705 433802 96771 433805
rect 94516 433800 96771 433802
rect 94516 433744 96710 433800
rect 96766 433744 96771 433800
rect 94516 433742 96771 433744
rect 94516 433740 94522 433742
rect 96705 433739 96771 433742
rect 99966 433740 99972 433804
rect 100036 433802 100042 433804
rect 100477 433802 100543 433805
rect 100036 433800 100543 433802
rect 100036 433744 100482 433800
rect 100538 433744 100543 433800
rect 100036 433742 100543 433744
rect 100036 433740 100042 433742
rect 100477 433739 100543 433742
rect 67817 433666 67883 433669
rect 71129 433666 71195 433669
rect 67817 433664 71195 433666
rect 67817 433608 67822 433664
rect 67878 433608 71134 433664
rect 71190 433608 71195 433664
rect 67817 433606 71195 433608
rect 67817 433603 67883 433606
rect 71129 433603 71195 433606
rect 74574 433604 74580 433668
rect 74644 433666 74650 433668
rect 74717 433666 74783 433669
rect 76373 433668 76439 433669
rect 76373 433666 76420 433668
rect 74644 433664 74783 433666
rect 74644 433608 74722 433664
rect 74778 433608 74783 433664
rect 74644 433606 74783 433608
rect 76328 433664 76420 433666
rect 76328 433608 76378 433664
rect 76328 433606 76420 433608
rect 74644 433604 74650 433606
rect 74717 433603 74783 433606
rect 76373 433604 76420 433606
rect 76484 433604 76490 433668
rect 77334 433604 77340 433668
rect 77404 433666 77410 433668
rect 78213 433666 78279 433669
rect 81893 433668 81959 433669
rect 84653 433668 84719 433669
rect 81893 433666 81940 433668
rect 77404 433664 78279 433666
rect 77404 433608 78218 433664
rect 78274 433608 78279 433664
rect 77404 433606 78279 433608
rect 81848 433664 81940 433666
rect 81848 433608 81898 433664
rect 81848 433606 81940 433608
rect 77404 433604 77410 433606
rect 76373 433603 76439 433604
rect 78213 433603 78279 433606
rect 81893 433604 81940 433606
rect 82004 433604 82010 433668
rect 84653 433666 84700 433668
rect 84608 433664 84700 433666
rect 84608 433608 84658 433664
rect 84608 433606 84700 433608
rect 84653 433604 84700 433606
rect 84764 433604 84770 433668
rect 85798 433604 85804 433668
rect 85868 433666 85874 433668
rect 85941 433666 86007 433669
rect 85868 433664 86007 433666
rect 85868 433608 85946 433664
rect 86002 433608 86007 433664
rect 85868 433606 86007 433608
rect 85868 433604 85874 433606
rect 81893 433603 81959 433604
rect 84653 433603 84719 433604
rect 85941 433603 86007 433606
rect 87086 433604 87092 433668
rect 87156 433666 87162 433668
rect 87229 433666 87295 433669
rect 87156 433664 87295 433666
rect 87156 433608 87234 433664
rect 87290 433608 87295 433664
rect 87156 433606 87295 433608
rect 87156 433604 87162 433606
rect 87229 433603 87295 433606
rect 87454 433604 87460 433668
rect 87524 433666 87530 433668
rect 89989 433666 90055 433669
rect 91185 433668 91251 433669
rect 91134 433666 91140 433668
rect 87524 433664 90055 433666
rect 87524 433608 89994 433664
rect 90050 433608 90055 433664
rect 87524 433606 90055 433608
rect 91094 433606 91140 433666
rect 91204 433664 91251 433668
rect 91246 433608 91251 433664
rect 87524 433604 87530 433606
rect 89989 433603 90055 433606
rect 91134 433604 91140 433606
rect 91204 433604 91251 433608
rect 92606 433604 92612 433668
rect 92676 433666 92682 433668
rect 92933 433666 92999 433669
rect 92676 433664 92999 433666
rect 92676 433608 92938 433664
rect 92994 433608 92999 433664
rect 92676 433606 92999 433608
rect 92676 433604 92682 433606
rect 91185 433603 91251 433604
rect 92933 433603 92999 433606
rect 96337 433666 96403 433669
rect 98177 433668 98243 433669
rect 96470 433666 96476 433668
rect 96337 433664 96476 433666
rect 96337 433608 96342 433664
rect 96398 433608 96476 433664
rect 96337 433606 96476 433608
rect 96337 433603 96403 433606
rect 96470 433604 96476 433606
rect 96540 433604 96546 433668
rect 98126 433666 98132 433668
rect 98086 433606 98132 433666
rect 98196 433664 98243 433668
rect 98238 433608 98243 433664
rect 98126 433604 98132 433606
rect 98196 433604 98243 433608
rect 98310 433604 98316 433668
rect 98380 433666 98386 433668
rect 98453 433666 98519 433669
rect 98380 433664 98519 433666
rect 98380 433608 98458 433664
rect 98514 433608 98519 433664
rect 98380 433606 98519 433608
rect 98380 433604 98386 433606
rect 98177 433603 98243 433604
rect 98453 433603 98519 433606
rect 99833 433666 99899 433669
rect 100150 433666 100156 433668
rect 99833 433664 100156 433666
rect 99833 433608 99838 433664
rect 99894 433608 100156 433664
rect 99833 433606 100156 433608
rect 99833 433603 99899 433606
rect 100150 433604 100156 433606
rect 100220 433604 100226 433668
rect 102542 433604 102548 433668
rect 102612 433666 102618 433668
rect 104709 433666 104775 433669
rect 102612 433664 104775 433666
rect 102612 433608 104714 433664
rect 104770 433608 104775 433664
rect 102612 433606 104775 433608
rect 102612 433604 102618 433606
rect 104709 433603 104775 433606
rect 106406 433604 106412 433668
rect 106476 433666 106482 433668
rect 106733 433666 106799 433669
rect 109033 433668 109099 433669
rect 110689 433668 110755 433669
rect 111793 433668 111859 433669
rect 108982 433666 108988 433668
rect 106476 433664 106799 433666
rect 106476 433608 106738 433664
rect 106794 433608 106799 433664
rect 106476 433606 106799 433608
rect 108906 433606 108988 433666
rect 109052 433664 109099 433668
rect 110638 433666 110644 433668
rect 109094 433608 109099 433664
rect 106476 433604 106482 433606
rect 106733 433603 106799 433606
rect 108982 433604 108988 433606
rect 109052 433604 109099 433608
rect 110598 433606 110644 433666
rect 110708 433664 110755 433668
rect 111742 433666 111748 433668
rect 110750 433608 110755 433664
rect 110638 433604 110644 433606
rect 110708 433604 110755 433608
rect 111702 433606 111748 433666
rect 111812 433664 111859 433668
rect 111854 433608 111859 433664
rect 111742 433604 111748 433606
rect 111812 433604 111859 433608
rect 109033 433603 109099 433604
rect 110689 433603 110755 433604
rect 111793 433603 111859 433604
rect 191649 433666 191715 433669
rect 255405 433666 255471 433669
rect 191649 433664 193660 433666
rect 191649 433608 191654 433664
rect 191710 433608 193660 433664
rect 191649 433606 193660 433608
rect 253460 433664 255471 433666
rect 253460 433608 255410 433664
rect 255466 433608 255471 433664
rect 253460 433606 255471 433608
rect 191649 433603 191715 433606
rect 255405 433603 255471 433606
rect 53557 433394 53623 433397
rect 65793 433394 65859 433397
rect 115013 433394 115079 433397
rect 53557 433392 68908 433394
rect 53557 433336 53562 433392
rect 53618 433336 65798 433392
rect 65854 433336 68908 433392
rect 53557 433334 68908 433336
rect 112700 433392 115079 433394
rect 112700 433336 115018 433392
rect 115074 433336 115079 433392
rect 112700 433334 115079 433336
rect 53557 433331 53623 433334
rect 65793 433331 65859 433334
rect 115013 433331 115079 433334
rect 68645 433122 68711 433125
rect 68645 433120 68938 433122
rect 68645 433064 68650 433120
rect 68706 433064 68938 433120
rect 68645 433062 68938 433064
rect 68645 433059 68711 433062
rect 68878 432548 68938 433062
rect 112110 432788 112116 432852
rect 112180 432788 112186 432852
rect 112118 432276 112178 432788
rect 188797 432578 188863 432581
rect 193438 432578 193444 432580
rect 188797 432576 193444 432578
rect 188797 432520 188802 432576
rect 188858 432520 193444 432576
rect 188797 432518 193444 432520
rect 188797 432515 188863 432518
rect 193438 432516 193444 432518
rect 193508 432516 193514 432580
rect 186957 432034 187023 432037
rect 193630 432034 193690 432276
rect 253933 432034 253999 432037
rect 186957 432032 193690 432034
rect 186957 431976 186962 432032
rect 187018 431976 193690 432032
rect 186957 431974 193690 431976
rect 253460 432032 253999 432034
rect 253460 431976 253938 432032
rect 253994 431976 253999 432032
rect 253460 431974 253999 431976
rect 186957 431971 187023 431974
rect 253933 431971 253999 431974
rect 582373 431626 582439 431629
rect 583520 431626 584960 431716
rect 582373 431624 584960 431626
rect 582373 431568 582378 431624
rect 582434 431568 584960 431624
rect 582373 431566 584960 431568
rect 582373 431563 582439 431566
rect 66253 431490 66319 431493
rect 66253 431488 68908 431490
rect 66253 431432 66258 431488
rect 66314 431432 68908 431488
rect 583520 431476 584960 431566
rect 66253 431430 68908 431432
rect 66253 431427 66319 431430
rect 115289 431218 115355 431221
rect 112700 431216 115355 431218
rect 112700 431160 115294 431216
rect 115350 431160 115355 431216
rect 112700 431158 115355 431160
rect 115289 431155 115355 431158
rect 193254 430884 193260 430948
rect 193324 430946 193330 430948
rect 193324 430886 193660 430946
rect 193324 430884 193330 430886
rect 255589 430674 255655 430677
rect 253460 430672 255655 430674
rect 253460 430616 255594 430672
rect 255650 430616 255655 430672
rect 253460 430614 255655 430616
rect 255589 430611 255655 430614
rect 67173 430402 67239 430405
rect 67173 430400 68908 430402
rect 67173 430344 67178 430400
rect 67234 430344 68908 430400
rect 67173 430342 68908 430344
rect 67173 430339 67239 430342
rect 115841 430130 115907 430133
rect 112700 430128 115907 430130
rect 112700 430072 115846 430128
rect 115902 430072 115907 430128
rect 112700 430070 115907 430072
rect 115841 430067 115907 430070
rect 67817 429858 67883 429861
rect 67817 429856 68938 429858
rect 67817 429800 67822 429856
rect 67878 429800 68938 429856
rect 67817 429798 68938 429800
rect 67817 429795 67883 429798
rect 68878 429284 68938 429798
rect 191189 429586 191255 429589
rect 191465 429586 191531 429589
rect 191189 429584 193660 429586
rect 191189 429528 191194 429584
rect 191250 429528 191470 429584
rect 191526 429528 193660 429584
rect 191189 429526 193660 429528
rect 191189 429523 191255 429526
rect 191465 429523 191531 429526
rect 114645 429314 114711 429317
rect 256601 429314 256667 429317
rect 112700 429312 114711 429314
rect 112700 429256 114650 429312
rect 114706 429256 114711 429312
rect 112700 429254 114711 429256
rect 253460 429312 256667 429314
rect 253460 429256 256606 429312
rect 256662 429256 256667 429312
rect 253460 429254 256667 429256
rect 114645 429251 114711 429254
rect 256601 429251 256667 429254
rect 66253 428226 66319 428229
rect 115841 428226 115907 428229
rect 66253 428224 68908 428226
rect 66253 428168 66258 428224
rect 66314 428168 68908 428224
rect 66253 428166 68908 428168
rect 112700 428224 115907 428226
rect 112700 428168 115846 428224
rect 115902 428168 115907 428224
rect 112700 428166 115907 428168
rect 66253 428163 66319 428166
rect 115841 428163 115907 428166
rect 191557 428226 191623 428229
rect 191557 428224 193660 428226
rect 191557 428168 191562 428224
rect 191618 428168 193660 428224
rect 191557 428166 193660 428168
rect 191557 428163 191623 428166
rect 255405 427954 255471 427957
rect 253460 427952 255471 427954
rect 253460 427896 255410 427952
rect 255466 427896 255471 427952
rect 253460 427894 255471 427896
rect 255405 427891 255471 427894
rect 66897 427410 66963 427413
rect 66897 427408 68908 427410
rect 66897 427352 66902 427408
rect 66958 427352 68908 427408
rect 66897 427350 68908 427352
rect 66897 427347 66963 427350
rect 115841 427138 115907 427141
rect 112700 427136 115907 427138
rect 112700 427080 115846 427136
rect 115902 427080 115907 427136
rect 112700 427078 115907 427080
rect 115841 427075 115907 427078
rect 191557 426866 191623 426869
rect 191557 426864 193660 426866
rect 191557 426808 191562 426864
rect 191618 426808 193660 426864
rect 191557 426806 193660 426808
rect 191557 426803 191623 426806
rect 255497 426594 255563 426597
rect 253460 426592 255563 426594
rect 253460 426536 255502 426592
rect 255558 426536 255563 426592
rect 253460 426534 255563 426536
rect 255497 426531 255563 426534
rect 69430 426188 69490 426292
rect 69422 426124 69428 426188
rect 69492 426124 69498 426188
rect 69430 425642 69490 426124
rect 113449 426050 113515 426053
rect 115289 426050 115355 426053
rect 112700 426048 115355 426050
rect 112700 425992 113454 426048
rect 113510 425992 115294 426048
rect 115350 425992 115355 426048
rect 112700 425990 115355 425992
rect 113449 425987 113515 425990
rect 115289 425987 115355 425990
rect 64830 425582 69490 425642
rect 60641 425098 60707 425101
rect 64830 425098 64890 425582
rect 191005 425506 191071 425509
rect 191833 425506 191899 425509
rect 191005 425504 193660 425506
rect 191005 425448 191010 425504
rect 191066 425448 191838 425504
rect 191894 425448 193660 425504
rect 191005 425446 193660 425448
rect 191005 425443 191071 425446
rect 191833 425443 191899 425446
rect 66621 425234 66687 425237
rect 256601 425234 256667 425237
rect 66621 425232 68908 425234
rect 66621 425176 66626 425232
rect 66682 425176 68908 425232
rect 66621 425174 68908 425176
rect 253460 425232 256667 425234
rect 253460 425176 256606 425232
rect 256662 425176 256667 425232
rect 253460 425174 256667 425176
rect 66621 425171 66687 425174
rect 256601 425171 256667 425174
rect 60641 425096 64890 425098
rect 60641 425040 60646 425096
rect 60702 425040 64890 425096
rect 60641 425038 64890 425040
rect 60641 425035 60707 425038
rect 115289 424962 115355 424965
rect 112700 424960 115355 424962
rect 112700 424904 115294 424960
rect 115350 424904 115355 424960
rect 112700 424902 115355 424904
rect 115289 424899 115355 424902
rect 255221 424282 255287 424285
rect 262254 424282 262260 424284
rect 255221 424280 262260 424282
rect 255221 424224 255226 424280
rect 255282 424224 262260 424280
rect 255221 424222 262260 424224
rect 255221 424219 255287 424222
rect 262254 424220 262260 424222
rect 262324 424220 262330 424284
rect 66805 424146 66871 424149
rect 115105 424146 115171 424149
rect 66805 424144 68908 424146
rect 66805 424088 66810 424144
rect 66866 424088 68908 424144
rect 66805 424086 68908 424088
rect 112700 424144 115171 424146
rect 112700 424088 115110 424144
rect 115166 424088 115171 424144
rect 112700 424086 115171 424088
rect 66805 424083 66871 424086
rect 115105 424083 115171 424086
rect 192845 423874 192911 423877
rect 192845 423872 193660 423874
rect 192845 423816 192850 423872
rect 192906 423816 193660 423872
rect 192845 423814 193660 423816
rect 192845 423811 192911 423814
rect -960 423602 480 423692
rect 3509 423602 3575 423605
rect 255497 423602 255563 423605
rect -960 423600 3575 423602
rect -960 423544 3514 423600
rect 3570 423544 3575 423600
rect -960 423542 3575 423544
rect 253460 423600 255563 423602
rect 253460 423544 255502 423600
rect 255558 423544 255563 423600
rect 253460 423542 255563 423544
rect -960 423452 480 423542
rect 3509 423539 3575 423542
rect 255497 423539 255563 423542
rect 66621 423330 66687 423333
rect 66621 423328 68908 423330
rect 66621 423272 66626 423328
rect 66682 423272 68908 423328
rect 66621 423270 68908 423272
rect 66621 423267 66687 423270
rect 115841 423058 115907 423061
rect 112700 423056 115907 423058
rect 112700 423000 115846 423056
rect 115902 423000 115907 423056
rect 112700 422998 115907 423000
rect 115841 422995 115907 422998
rect 190821 422514 190887 422517
rect 190821 422512 193660 422514
rect 190821 422456 190826 422512
rect 190882 422456 193660 422512
rect 190821 422454 193660 422456
rect 190821 422451 190887 422454
rect 57697 422242 57763 422245
rect 66805 422242 66871 422245
rect 255497 422242 255563 422245
rect 57697 422240 64890 422242
rect 57697 422184 57702 422240
rect 57758 422184 64890 422240
rect 57697 422182 64890 422184
rect 57697 422179 57763 422182
rect 64830 421834 64890 422182
rect 66805 422240 68908 422242
rect 66805 422184 66810 422240
rect 66866 422184 68908 422240
rect 66805 422182 68908 422184
rect 253460 422240 255563 422242
rect 253460 422184 255502 422240
rect 255558 422184 255563 422240
rect 253460 422182 255563 422184
rect 66805 422179 66871 422182
rect 255497 422179 255563 422182
rect 114645 421970 114711 421973
rect 112700 421968 114711 421970
rect 112700 421912 114650 421968
rect 114706 421912 114711 421968
rect 112700 421910 114711 421912
rect 114645 421907 114711 421910
rect 64830 421774 68938 421834
rect 68878 421124 68938 421774
rect 188838 420956 188844 421020
rect 188908 421018 188914 421020
rect 193630 421018 193690 421124
rect 188908 420958 193690 421018
rect 188908 420956 188914 420958
rect 114553 420882 114619 420885
rect 255589 420882 255655 420885
rect 112700 420880 114619 420882
rect 112700 420824 114558 420880
rect 114614 420824 114619 420880
rect 112700 420822 114619 420824
rect 253460 420880 255655 420882
rect 253460 420824 255594 420880
rect 255650 420824 255655 420880
rect 253460 420822 255655 420824
rect 114553 420819 114619 420822
rect 255589 420819 255655 420822
rect 66897 420066 66963 420069
rect 115841 420066 115907 420069
rect 66897 420064 68908 420066
rect 66897 420008 66902 420064
rect 66958 420008 68908 420064
rect 66897 420006 68908 420008
rect 112700 420064 115907 420066
rect 112700 420008 115846 420064
rect 115902 420008 115907 420064
rect 112700 420006 115907 420008
rect 66897 420003 66963 420006
rect 115841 420003 115907 420006
rect 191557 419794 191623 419797
rect 191557 419792 193660 419794
rect 191557 419736 191562 419792
rect 191618 419736 193660 419792
rect 191557 419734 193660 419736
rect 191557 419731 191623 419734
rect 255497 419522 255563 419525
rect 253460 419520 255563 419522
rect 253460 419464 255502 419520
rect 255558 419464 255563 419520
rect 253460 419462 255563 419464
rect 255497 419459 255563 419462
rect 66805 418978 66871 418981
rect 115197 418978 115263 418981
rect 66805 418976 68908 418978
rect 66805 418920 66810 418976
rect 66866 418920 68908 418976
rect 66805 418918 68908 418920
rect 112700 418976 115263 418978
rect 112700 418920 115202 418976
rect 115258 418920 115263 418976
rect 112700 418918 115263 418920
rect 66805 418915 66871 418918
rect 115197 418915 115263 418918
rect 191557 418434 191623 418437
rect 191557 418432 193660 418434
rect 191557 418376 191562 418432
rect 191618 418376 193660 418432
rect 191557 418374 193660 418376
rect 191557 418371 191623 418374
rect 114318 418236 114324 418300
rect 114388 418298 114394 418300
rect 116117 418298 116183 418301
rect 186957 418298 187023 418301
rect 114388 418296 187023 418298
rect 114388 418240 116122 418296
rect 116178 418240 186962 418296
rect 187018 418240 187023 418296
rect 114388 418238 187023 418240
rect 114388 418236 114394 418238
rect 116117 418235 116183 418238
rect 186957 418235 187023 418238
rect 582925 418298 582991 418301
rect 583520 418298 584960 418388
rect 582925 418296 584960 418298
rect 582925 418240 582930 418296
rect 582986 418240 584960 418296
rect 582925 418238 584960 418240
rect 582925 418235 582991 418238
rect 67449 418162 67515 418165
rect 67633 418162 67699 418165
rect 255589 418162 255655 418165
rect 67449 418160 68908 418162
rect 67449 418104 67454 418160
rect 67510 418104 67638 418160
rect 67694 418104 68908 418160
rect 67449 418102 68908 418104
rect 253460 418160 255655 418162
rect 253460 418104 255594 418160
rect 255650 418104 255655 418160
rect 583520 418148 584960 418238
rect 253460 418102 255655 418104
rect 67449 418099 67515 418102
rect 67633 418099 67699 418102
rect 255589 418099 255655 418102
rect 114686 417890 114692 417892
rect 112700 417830 114692 417890
rect 114686 417828 114692 417830
rect 114756 417828 114762 417892
rect 124857 417482 124923 417485
rect 128445 417482 128511 417485
rect 124857 417480 128511 417482
rect 124857 417424 124862 417480
rect 124918 417424 128450 417480
rect 128506 417424 128511 417480
rect 124857 417422 128511 417424
rect 124857 417419 124923 417422
rect 128445 417419 128511 417422
rect 66989 417074 67055 417077
rect 191557 417074 191623 417077
rect 66989 417072 68908 417074
rect 66989 417016 66994 417072
rect 67050 417016 68908 417072
rect 66989 417014 68908 417016
rect 191557 417072 193660 417074
rect 191557 417016 191562 417072
rect 191618 417016 193660 417072
rect 191557 417014 193660 417016
rect 66989 417011 67055 417014
rect 191557 417011 191623 417014
rect 113265 416802 113331 416805
rect 115841 416802 115907 416805
rect 255497 416802 255563 416805
rect 112700 416800 115907 416802
rect 112700 416744 113270 416800
rect 113326 416744 115846 416800
rect 115902 416744 115907 416800
rect 112700 416742 115907 416744
rect 253460 416800 255563 416802
rect 253460 416744 255502 416800
rect 255558 416744 255563 416800
rect 253460 416742 255563 416744
rect 113265 416739 113331 416742
rect 115841 416739 115907 416742
rect 255497 416739 255563 416742
rect 66897 415986 66963 415989
rect 66897 415984 68908 415986
rect 66897 415928 66902 415984
rect 66958 415928 68908 415984
rect 66897 415926 68908 415928
rect 66897 415923 66963 415926
rect 115841 415714 115907 415717
rect 112700 415712 115907 415714
rect 112700 415656 115846 415712
rect 115902 415656 115907 415712
rect 112700 415654 115907 415656
rect 115841 415651 115907 415654
rect 191005 415442 191071 415445
rect 191005 415440 193660 415442
rect 191005 415384 191010 415440
rect 191066 415384 193660 415440
rect 191005 415382 193660 415384
rect 191005 415379 191071 415382
rect 256601 415170 256667 415173
rect 253460 415168 256667 415170
rect 253460 415112 256606 415168
rect 256662 415112 256667 415168
rect 253460 415110 256667 415112
rect 256601 415107 256667 415110
rect 66713 414898 66779 414901
rect 113173 414898 113239 414901
rect 116025 414898 116091 414901
rect 66713 414896 68908 414898
rect 66713 414840 66718 414896
rect 66774 414840 68908 414896
rect 66713 414838 68908 414840
rect 112700 414896 116091 414898
rect 112700 414840 113178 414896
rect 113234 414840 116030 414896
rect 116086 414840 116091 414896
rect 112700 414838 116091 414840
rect 66713 414835 66779 414838
rect 113173 414835 113239 414838
rect 116025 414835 116091 414838
rect 67265 414082 67331 414085
rect 115013 414082 115079 414085
rect 188286 414082 188292 414084
rect 67265 414080 68908 414082
rect 67265 414024 67270 414080
rect 67326 414024 68908 414080
rect 67265 414022 68908 414024
rect 115013 414080 188292 414082
rect 115013 414024 115018 414080
rect 115074 414024 188292 414080
rect 115013 414022 188292 414024
rect 67265 414019 67331 414022
rect 115013 414019 115079 414022
rect 188286 414020 188292 414022
rect 188356 414020 188362 414084
rect 191557 414082 191623 414085
rect 191557 414080 193660 414082
rect 191557 414024 191562 414080
rect 191618 414024 193660 414080
rect 191557 414022 193660 414024
rect 191557 414019 191623 414022
rect 115841 413810 115907 413813
rect 254117 413810 254183 413813
rect 112700 413808 115907 413810
rect 112700 413752 115846 413808
rect 115902 413752 115907 413808
rect 112700 413750 115907 413752
rect 253460 413808 254183 413810
rect 253460 413752 254122 413808
rect 254178 413752 254183 413808
rect 253460 413750 254183 413752
rect 115841 413747 115907 413750
rect 254117 413747 254183 413750
rect 66253 412994 66319 412997
rect 66253 412992 68908 412994
rect 66253 412936 66258 412992
rect 66314 412936 68908 412992
rect 66253 412934 68908 412936
rect 66253 412931 66319 412934
rect 115013 412722 115079 412725
rect 112700 412720 115079 412722
rect 112700 412664 115018 412720
rect 115074 412664 115079 412720
rect 112700 412662 115079 412664
rect 115013 412659 115079 412662
rect 190269 412722 190335 412725
rect 190269 412720 193660 412722
rect 190269 412664 190274 412720
rect 190330 412664 193660 412720
rect 190269 412662 193660 412664
rect 190269 412659 190335 412662
rect 255497 412450 255563 412453
rect 253460 412448 255563 412450
rect 253460 412392 255502 412448
rect 255558 412392 255563 412448
rect 253460 412390 255563 412392
rect 255497 412387 255563 412390
rect 66805 411906 66871 411909
rect 66805 411904 68908 411906
rect 66805 411848 66810 411904
rect 66866 411848 68908 411904
rect 66805 411846 68908 411848
rect 66805 411843 66871 411846
rect 116117 411634 116183 411637
rect 112700 411632 116183 411634
rect 112700 411576 116122 411632
rect 116178 411576 116183 411632
rect 112700 411574 116183 411576
rect 116117 411571 116183 411574
rect 191465 411362 191531 411365
rect 191465 411360 193660 411362
rect 191465 411304 191470 411360
rect 191526 411304 193660 411360
rect 191465 411302 193660 411304
rect 191465 411299 191531 411302
rect 255497 411090 255563 411093
rect 253460 411088 255563 411090
rect 253460 411032 255502 411088
rect 255558 411032 255563 411088
rect 253460 411030 255563 411032
rect 255497 411027 255563 411030
rect 66897 410818 66963 410821
rect 66897 410816 68908 410818
rect 66897 410760 66902 410816
rect 66958 410760 68908 410816
rect 66897 410758 68908 410760
rect 66897 410755 66963 410758
rect -960 410546 480 410636
rect 2957 410546 3023 410549
rect 114502 410546 114508 410548
rect -960 410544 3023 410546
rect -960 410488 2962 410544
rect 3018 410488 3023 410544
rect -960 410486 3023 410488
rect 112700 410486 114508 410546
rect -960 410396 480 410486
rect 2957 410483 3023 410486
rect 114502 410484 114508 410486
rect 114572 410546 114578 410548
rect 115841 410546 115907 410549
rect 114572 410544 115907 410546
rect 114572 410488 115846 410544
rect 115902 410488 115907 410544
rect 114572 410486 115907 410488
rect 114572 410484 114578 410486
rect 115841 410483 115907 410486
rect 190821 410002 190887 410005
rect 190821 410000 193660 410002
rect 190821 409944 190826 410000
rect 190882 409944 193660 410000
rect 190821 409942 193660 409944
rect 190821 409939 190887 409942
rect 67766 409668 67772 409732
rect 67836 409730 67842 409732
rect 115841 409730 115907 409733
rect 255497 409730 255563 409733
rect 67836 409670 68908 409730
rect 112700 409728 115907 409730
rect 112700 409672 115846 409728
rect 115902 409672 115907 409728
rect 112700 409670 115907 409672
rect 253460 409728 255563 409730
rect 253460 409672 255502 409728
rect 255558 409672 255563 409728
rect 253460 409670 255563 409672
rect 67836 409668 67842 409670
rect 115841 409667 115907 409670
rect 255497 409667 255563 409670
rect 66805 408914 66871 408917
rect 66805 408912 68908 408914
rect 66805 408856 66810 408912
rect 66866 408856 68908 408912
rect 66805 408854 68908 408856
rect 66805 408851 66871 408854
rect 115841 408642 115907 408645
rect 112700 408640 115907 408642
rect 112700 408584 115846 408640
rect 115902 408584 115907 408640
rect 112700 408582 115907 408584
rect 115841 408579 115907 408582
rect 193029 408642 193095 408645
rect 193029 408640 193660 408642
rect 193029 408584 193034 408640
rect 193090 408584 193660 408640
rect 193029 408582 193660 408584
rect 193029 408579 193095 408582
rect 255497 408370 255563 408373
rect 253460 408368 255563 408370
rect 253460 408312 255502 408368
rect 255558 408312 255563 408368
rect 253460 408310 255563 408312
rect 255497 408307 255563 408310
rect 66805 407826 66871 407829
rect 66805 407824 68908 407826
rect 66805 407768 66810 407824
rect 66866 407768 68908 407824
rect 66805 407766 68908 407768
rect 66805 407763 66871 407766
rect 115841 407554 115907 407557
rect 112700 407552 115907 407554
rect 112700 407496 115846 407552
rect 115902 407496 115907 407552
rect 112700 407494 115907 407496
rect 115841 407491 115907 407494
rect 112713 407010 112779 407013
rect 112670 407008 112779 407010
rect 112670 406952 112718 407008
rect 112774 406952 112779 407008
rect 112670 406947 112779 406952
rect 191465 407010 191531 407013
rect 255497 407010 255563 407013
rect 191465 407008 193660 407010
rect 191465 406952 191470 407008
rect 191526 406952 193660 407008
rect 191465 406950 193660 406952
rect 253460 407008 255563 407010
rect 253460 406952 255502 407008
rect 255558 406952 255563 407008
rect 253460 406950 255563 406952
rect 191465 406947 191531 406950
rect 255497 406947 255563 406950
rect 68878 406058 68938 406708
rect 112670 406466 112730 406947
rect 115197 406466 115263 406469
rect 112670 406464 115263 406466
rect 112670 406436 115202 406464
rect 112700 406408 115202 406436
rect 115258 406408 115263 406464
rect 112700 406406 115263 406408
rect 115197 406403 115263 406406
rect 116669 406330 116735 406333
rect 125777 406330 125843 406333
rect 166257 406330 166323 406333
rect 116669 406328 166323 406330
rect 116669 406272 116674 406328
rect 116730 406272 125782 406328
rect 125838 406272 166262 406328
rect 166318 406272 166323 406328
rect 116669 406270 166323 406272
rect 116669 406267 116735 406270
rect 125777 406267 125843 406270
rect 166257 406267 166323 406270
rect 64830 405998 68938 406058
rect 59118 405724 59124 405788
rect 59188 405786 59194 405788
rect 63401 405786 63467 405789
rect 64830 405786 64890 405998
rect 59188 405784 64890 405786
rect 59188 405728 63406 405784
rect 63462 405728 64890 405784
rect 59188 405726 64890 405728
rect 59188 405724 59194 405726
rect 63401 405723 63467 405726
rect 67357 405650 67423 405653
rect 115381 405650 115447 405653
rect 115749 405650 115815 405653
rect 67357 405648 68908 405650
rect 67357 405592 67362 405648
rect 67418 405592 68908 405648
rect 67357 405590 68908 405592
rect 112700 405648 115815 405650
rect 112700 405592 115386 405648
rect 115442 405592 115754 405648
rect 115810 405592 115815 405648
rect 112700 405590 115815 405592
rect 67357 405587 67423 405590
rect 115381 405587 115447 405590
rect 115749 405587 115815 405590
rect 191373 405650 191439 405653
rect 191373 405648 193660 405650
rect 191373 405592 191378 405648
rect 191434 405592 193660 405648
rect 191373 405590 193660 405592
rect 191373 405587 191439 405590
rect 252878 404836 252938 405348
rect 583201 404970 583267 404973
rect 583520 404970 584960 405060
rect 583201 404968 584960 404970
rect 583201 404912 583206 404968
rect 583262 404912 584960 404968
rect 583201 404910 584960 404912
rect 583201 404907 583267 404910
rect 252870 404772 252876 404836
rect 252940 404772 252946 404836
rect 583520 404820 584960 404910
rect 66897 404562 66963 404565
rect 115841 404562 115907 404565
rect 66897 404560 68908 404562
rect 66897 404504 66902 404560
rect 66958 404504 68908 404560
rect 66897 404502 68908 404504
rect 112700 404560 115907 404562
rect 112700 404504 115846 404560
rect 115902 404504 115907 404560
rect 112700 404502 115907 404504
rect 66897 404499 66963 404502
rect 115841 404499 115907 404502
rect 191465 404290 191531 404293
rect 191465 404288 193660 404290
rect 191465 404232 191470 404288
rect 191526 404232 193660 404288
rect 191465 404230 193660 404232
rect 191465 404227 191531 404230
rect 255497 404018 255563 404021
rect 253460 404016 255563 404018
rect 253460 403960 255502 404016
rect 255558 403960 255563 404016
rect 253460 403958 255563 403960
rect 255497 403955 255563 403958
rect 66805 403746 66871 403749
rect 66805 403744 68908 403746
rect 66805 403688 66810 403744
rect 66866 403688 68908 403744
rect 66805 403686 68908 403688
rect 66805 403683 66871 403686
rect 258717 403610 258783 403613
rect 270534 403610 270540 403612
rect 258717 403608 270540 403610
rect 258717 403552 258722 403608
rect 258778 403552 270540 403608
rect 258717 403550 270540 403552
rect 258717 403547 258783 403550
rect 270534 403548 270540 403550
rect 270604 403548 270610 403612
rect 115841 403474 115907 403477
rect 112700 403472 115907 403474
rect 112700 403416 115846 403472
rect 115902 403416 115907 403472
rect 112700 403414 115907 403416
rect 115841 403411 115907 403414
rect 191373 402930 191439 402933
rect 191373 402928 193660 402930
rect 191373 402872 191378 402928
rect 191434 402872 193660 402928
rect 191373 402870 193660 402872
rect 191373 402867 191439 402870
rect 67541 402658 67607 402661
rect 254209 402658 254275 402661
rect 67541 402656 68908 402658
rect 67541 402600 67546 402656
rect 67602 402600 68908 402656
rect 67541 402598 68908 402600
rect 253460 402656 254275 402658
rect 253460 402600 254214 402656
rect 254270 402600 254275 402656
rect 253460 402598 254275 402600
rect 67541 402595 67607 402598
rect 254209 402595 254275 402598
rect 113357 402386 113423 402389
rect 112700 402384 113423 402386
rect 112700 402356 113362 402384
rect 112670 402328 113362 402356
rect 113418 402328 113423 402384
rect 112670 402326 113423 402328
rect 112670 401845 112730 402326
rect 113357 402323 113423 402326
rect 112670 401840 112779 401845
rect 112670 401784 112718 401840
rect 112774 401784 112779 401840
rect 112670 401782 112779 401784
rect 112713 401779 112779 401782
rect 67265 401706 67331 401709
rect 67541 401706 67607 401709
rect 67265 401704 67607 401706
rect 67265 401648 67270 401704
rect 67326 401648 67546 401704
rect 67602 401648 67607 401704
rect 67265 401646 67607 401648
rect 67265 401643 67331 401646
rect 67541 401643 67607 401646
rect 66713 401570 66779 401573
rect 191465 401570 191531 401573
rect 66713 401568 68908 401570
rect 66713 401512 66718 401568
rect 66774 401512 68908 401568
rect 66713 401510 68908 401512
rect 191465 401568 193660 401570
rect 191465 401512 191470 401568
rect 191526 401512 193660 401568
rect 191465 401510 193660 401512
rect 66713 401507 66779 401510
rect 191465 401507 191531 401510
rect 115657 401298 115723 401301
rect 255497 401298 255563 401301
rect 112700 401296 115723 401298
rect 112700 401240 115662 401296
rect 115718 401240 115723 401296
rect 112700 401238 115723 401240
rect 253460 401296 255563 401298
rect 253460 401240 255502 401296
rect 255558 401240 255563 401296
rect 253460 401238 255563 401240
rect 115657 401235 115723 401238
rect 255497 401235 255563 401238
rect 124857 400890 124923 400893
rect 187049 400890 187115 400893
rect 124857 400888 187115 400890
rect 124857 400832 124862 400888
rect 124918 400832 187054 400888
rect 187110 400832 187115 400888
rect 124857 400830 187115 400832
rect 124857 400827 124923 400830
rect 187049 400827 187115 400830
rect 67357 400482 67423 400485
rect 114737 400482 114803 400485
rect 67357 400480 68908 400482
rect 67357 400424 67362 400480
rect 67418 400424 68908 400480
rect 67357 400422 68908 400424
rect 112700 400480 114803 400482
rect 112700 400424 114742 400480
rect 114798 400424 114803 400480
rect 112700 400422 114803 400424
rect 67357 400419 67423 400422
rect 114737 400419 114803 400422
rect 190821 400210 190887 400213
rect 190821 400208 193660 400210
rect 190821 400152 190826 400208
rect 190882 400152 193660 400208
rect 190821 400150 193660 400152
rect 190821 400147 190887 400150
rect 255497 399938 255563 399941
rect 253460 399936 255563 399938
rect 253460 399880 255502 399936
rect 255558 399880 255563 399936
rect 253460 399878 255563 399880
rect 255497 399875 255563 399878
rect 67541 399666 67607 399669
rect 67541 399664 68908 399666
rect 67541 399608 67546 399664
rect 67602 399608 68908 399664
rect 67541 399606 68908 399608
rect 67541 399603 67607 399606
rect 48221 399530 48287 399533
rect 48221 399528 64890 399530
rect 48221 399472 48226 399528
rect 48282 399472 64890 399528
rect 48221 399470 64890 399472
rect 48221 399467 48287 399470
rect 64830 398850 64890 399470
rect 115841 399394 115907 399397
rect 112700 399392 115907 399394
rect 112700 399336 115846 399392
rect 115902 399336 115907 399392
rect 112700 399334 115907 399336
rect 115841 399331 115907 399334
rect 66662 398850 66668 398852
rect 64830 398790 66668 398850
rect 66662 398788 66668 398790
rect 66732 398850 66738 398852
rect 66732 398790 68938 398850
rect 66732 398788 66738 398790
rect 68878 398548 68938 398790
rect 191097 398578 191163 398581
rect 255497 398578 255563 398581
rect 191097 398576 193660 398578
rect 191097 398520 191102 398576
rect 191158 398520 193660 398576
rect 191097 398518 193660 398520
rect 253460 398576 255563 398578
rect 253460 398520 255502 398576
rect 255558 398520 255563 398576
rect 253460 398518 255563 398520
rect 191097 398515 191163 398518
rect 255497 398515 255563 398518
rect 115565 398306 115631 398309
rect 112700 398304 115631 398306
rect 112700 398248 115570 398304
rect 115626 398248 115631 398304
rect 112700 398246 115631 398248
rect 115565 398243 115631 398246
rect -960 397490 480 397580
rect 3509 397490 3575 397493
rect -960 397488 3575 397490
rect -960 397432 3514 397488
rect 3570 397432 3575 397488
rect -960 397430 3575 397432
rect -960 397340 480 397430
rect 3509 397427 3575 397430
rect 67725 397490 67791 397493
rect 116577 397490 116643 397493
rect 119337 397490 119403 397493
rect 67725 397488 68908 397490
rect 67725 397432 67730 397488
rect 67786 397432 68908 397488
rect 67725 397430 68908 397432
rect 115844 397488 119403 397490
rect 115844 397432 116582 397488
rect 116638 397432 119342 397488
rect 119398 397432 119403 397488
rect 115844 397430 119403 397432
rect 67725 397427 67791 397430
rect 115844 397218 115904 397430
rect 116577 397427 116643 397430
rect 119337 397427 119403 397430
rect 112700 397158 115904 397218
rect 191465 397218 191531 397221
rect 191465 397216 193660 397218
rect 191465 397160 191470 397216
rect 191526 397160 193660 397216
rect 191465 397158 193660 397160
rect 191465 397155 191531 397158
rect 255497 396946 255563 396949
rect 253460 396944 255563 396946
rect 253460 396888 255502 396944
rect 255558 396888 255563 396944
rect 253460 396886 255563 396888
rect 255497 396883 255563 396886
rect 160686 396612 160692 396676
rect 160756 396674 160762 396676
rect 176745 396674 176811 396677
rect 160756 396672 176811 396674
rect 160756 396616 176750 396672
rect 176806 396616 176811 396672
rect 160756 396614 176811 396616
rect 160756 396612 160762 396614
rect 176745 396611 176811 396614
rect 67725 396402 67791 396405
rect 67950 396402 67956 396404
rect 67725 396400 67956 396402
rect 67725 396344 67730 396400
rect 67786 396344 67956 396400
rect 67725 396342 67956 396344
rect 67725 396339 67791 396342
rect 67950 396340 67956 396342
rect 68020 396402 68026 396404
rect 113214 396402 113220 396404
rect 68020 396342 68908 396402
rect 112700 396342 113220 396402
rect 68020 396340 68026 396342
rect 113214 396340 113220 396342
rect 113284 396402 113290 396404
rect 115841 396402 115907 396405
rect 113284 396400 115907 396402
rect 113284 396344 115846 396400
rect 115902 396344 115907 396400
rect 113284 396342 115907 396344
rect 113284 396340 113290 396342
rect 115841 396339 115907 396342
rect 67173 395314 67239 395317
rect 115841 395314 115907 395317
rect 67173 395312 68908 395314
rect 67173 395256 67178 395312
rect 67234 395256 68908 395312
rect 67173 395254 68908 395256
rect 112700 395312 115907 395314
rect 112700 395256 115846 395312
rect 115902 395256 115907 395312
rect 112700 395254 115907 395256
rect 67173 395251 67239 395254
rect 115841 395251 115907 395254
rect 190177 394770 190243 394773
rect 193630 394770 193690 395828
rect 253974 395586 253980 395588
rect 253460 395526 253980 395586
rect 253974 395524 253980 395526
rect 254044 395524 254050 395588
rect 190177 394768 193690 394770
rect 190177 394712 190182 394768
rect 190238 394712 193690 394768
rect 190177 394710 193690 394712
rect 190177 394707 190243 394710
rect 66805 394498 66871 394501
rect 66805 394496 68908 394498
rect 66805 394440 66810 394496
rect 66866 394440 68908 394496
rect 66805 394438 68908 394440
rect 66805 394435 66871 394438
rect 115841 394226 115907 394229
rect 112700 394224 115907 394226
rect 112700 394168 115846 394224
rect 115902 394168 115907 394224
rect 112700 394166 115907 394168
rect 115841 394163 115907 394166
rect 65885 393410 65951 393413
rect 190085 393410 190151 393413
rect 193630 393410 193690 394468
rect 255589 394226 255655 394229
rect 253460 394224 255655 394226
rect 253460 394168 255594 394224
rect 255650 394168 255655 394224
rect 253460 394166 255655 394168
rect 255589 394163 255655 394166
rect 65885 393408 68908 393410
rect 65885 393352 65890 393408
rect 65946 393352 68908 393408
rect 65885 393350 68908 393352
rect 190085 393408 193690 393410
rect 190085 393352 190090 393408
rect 190146 393352 193690 393408
rect 190085 393350 193690 393352
rect 65885 393347 65951 393350
rect 190085 393347 190151 393350
rect 115841 393138 115907 393141
rect 112700 393136 115907 393138
rect 112700 393080 115846 393136
rect 115902 393080 115907 393136
rect 112700 393078 115907 393080
rect 115841 393075 115907 393078
rect 193814 392596 193874 393108
rect 253657 392866 253723 392869
rect 253460 392864 253723 392866
rect 253460 392808 253662 392864
rect 253718 392808 253723 392864
rect 253460 392806 253723 392808
rect 253657 392803 253723 392806
rect 193806 392532 193812 392596
rect 193876 392532 193882 392596
rect 66253 392322 66319 392325
rect 66253 392320 68908 392322
rect 66253 392264 66258 392320
rect 66314 392264 68908 392320
rect 66253 392262 68908 392264
rect 66253 392259 66319 392262
rect 67541 392050 67607 392053
rect 69606 392050 69612 392052
rect 67541 392048 69612 392050
rect 67541 391992 67546 392048
rect 67602 391992 69612 392048
rect 67541 391990 69612 391992
rect 67541 391987 67607 391990
rect 69606 391988 69612 391990
rect 69676 391988 69682 392052
rect 115381 392050 115447 392053
rect 112700 392048 115447 392050
rect 112700 391992 115386 392048
rect 115442 391992 115447 392048
rect 112700 391990 115447 391992
rect 115381 391987 115447 391990
rect 191465 391778 191531 391781
rect 191465 391776 193660 391778
rect 191465 391720 191470 391776
rect 191526 391720 193660 391776
rect 191465 391718 193660 391720
rect 191465 391715 191531 391718
rect 583520 391628 584960 391868
rect 55121 391506 55187 391509
rect 254025 391506 254091 391509
rect 55121 391504 64890 391506
rect 55121 391448 55126 391504
rect 55182 391448 64890 391504
rect 55121 391446 64890 391448
rect 253460 391504 254091 391506
rect 253460 391448 254030 391504
rect 254086 391448 254091 391504
rect 253460 391446 254091 391448
rect 55121 391443 55187 391446
rect 64830 390962 64890 391446
rect 254025 391443 254091 391446
rect 67541 391234 67607 391237
rect 114829 391234 114895 391237
rect 193305 391236 193371 391237
rect 193254 391234 193260 391236
rect 67541 391232 68908 391234
rect 67541 391176 67546 391232
rect 67602 391176 68908 391232
rect 67541 391174 68908 391176
rect 112700 391232 114895 391234
rect 112700 391176 114834 391232
rect 114890 391176 114895 391232
rect 112700 391174 114895 391176
rect 193214 391174 193260 391234
rect 193324 391232 193371 391236
rect 193366 391176 193371 391232
rect 67541 391171 67607 391174
rect 114829 391171 114895 391174
rect 193254 391172 193260 391174
rect 193324 391172 193371 391176
rect 193305 391171 193371 391172
rect 72509 390962 72575 390965
rect 64830 390960 72575 390962
rect 64830 390904 72514 390960
rect 72570 390904 72575 390960
rect 64830 390902 72575 390904
rect 72509 390899 72575 390902
rect 73470 390900 73476 390964
rect 73540 390962 73546 390964
rect 73981 390962 74047 390965
rect 73540 390960 74047 390962
rect 73540 390904 73986 390960
rect 74042 390904 74047 390960
rect 73540 390902 74047 390904
rect 73540 390900 73546 390902
rect 73981 390899 74047 390902
rect 76649 390962 76715 390965
rect 191005 390962 191071 390965
rect 76649 390960 191071 390962
rect 76649 390904 76654 390960
rect 76710 390904 191010 390960
rect 191066 390904 191071 390960
rect 76649 390902 191071 390904
rect 76649 390899 76715 390902
rect 191005 390899 191071 390902
rect 71129 390826 71195 390829
rect 195973 390826 196039 390829
rect 71129 390824 196039 390826
rect 71129 390768 71134 390824
rect 71190 390768 195978 390824
rect 196034 390768 196039 390824
rect 71129 390766 196039 390768
rect 71129 390763 71195 390766
rect 195973 390763 196039 390766
rect 82077 390692 82143 390693
rect 82077 390690 82124 390692
rect 82032 390688 82124 390690
rect 82032 390632 82082 390688
rect 82032 390630 82124 390632
rect 82077 390628 82124 390630
rect 82188 390628 82194 390692
rect 95325 390690 95391 390693
rect 96705 390692 96771 390693
rect 104249 390692 104315 390693
rect 96470 390690 96476 390692
rect 95325 390688 96476 390690
rect 95325 390632 95330 390688
rect 95386 390632 96476 390688
rect 95325 390630 96476 390632
rect 82077 390627 82143 390628
rect 95325 390627 95391 390630
rect 96470 390628 96476 390630
rect 96540 390628 96546 390692
rect 96654 390628 96660 390692
rect 96724 390690 96771 390692
rect 96724 390688 96816 390690
rect 96766 390632 96816 390688
rect 96724 390630 96816 390632
rect 96724 390628 96771 390630
rect 104198 390628 104204 390692
rect 104268 390690 104315 390692
rect 105077 390692 105143 390693
rect 107745 390692 107811 390693
rect 111977 390692 112043 390693
rect 105077 390690 105124 390692
rect 104268 390688 104360 390690
rect 104310 390632 104360 390688
rect 104268 390630 104360 390632
rect 105032 390688 105124 390690
rect 105032 390632 105082 390688
rect 105032 390630 105124 390632
rect 104268 390628 104315 390630
rect 96705 390627 96771 390628
rect 104249 390627 104315 390628
rect 105077 390628 105124 390630
rect 105188 390628 105194 390692
rect 107694 390628 107700 390692
rect 107764 390690 107811 390692
rect 107764 390688 107856 390690
rect 107806 390632 107856 390688
rect 107764 390630 107856 390632
rect 107764 390628 107811 390630
rect 111926 390628 111932 390692
rect 111996 390690 112043 390692
rect 111996 390688 112088 390690
rect 112038 390632 112088 390688
rect 111996 390630 112088 390632
rect 111996 390628 112043 390630
rect 105077 390627 105143 390628
rect 107745 390627 107811 390628
rect 111977 390627 112043 390628
rect 88742 390492 88748 390556
rect 88812 390554 88818 390556
rect 89253 390554 89319 390557
rect 88812 390552 89319 390554
rect 88812 390496 89258 390552
rect 89314 390496 89319 390552
rect 88812 390494 89319 390496
rect 88812 390492 88818 390494
rect 89253 390491 89319 390494
rect 100702 390492 100708 390556
rect 100772 390554 100778 390556
rect 100937 390554 101003 390557
rect 100772 390552 101506 390554
rect 100772 390496 100942 390552
rect 100998 390496 101506 390552
rect 100772 390494 101506 390496
rect 100772 390492 100778 390494
rect 100937 390491 101003 390494
rect 91318 390356 91324 390420
rect 91388 390418 91394 390420
rect 91921 390418 91987 390421
rect 91388 390416 91987 390418
rect 91388 390360 91926 390416
rect 91982 390360 91987 390416
rect 91388 390358 91987 390360
rect 91388 390356 91394 390358
rect 91921 390355 91987 390358
rect 96838 390356 96844 390420
rect 96908 390418 96914 390420
rect 96981 390418 97047 390421
rect 96908 390416 97047 390418
rect 96908 390360 96986 390416
rect 97042 390360 97047 390416
rect 96908 390358 97047 390360
rect 96908 390356 96914 390358
rect 96981 390355 97047 390358
rect 101446 390282 101506 390494
rect 104934 390492 104940 390556
rect 105004 390554 105010 390556
rect 105261 390554 105327 390557
rect 582557 390554 582623 390557
rect 105004 390552 105327 390554
rect 105004 390496 105266 390552
rect 105322 390496 105327 390552
rect 105004 390494 105327 390496
rect 105004 390492 105010 390494
rect 105261 390491 105327 390494
rect 258030 390552 582623 390554
rect 258030 390496 582562 390552
rect 582618 390496 582623 390552
rect 258030 390494 582623 390496
rect 102041 390282 102107 390285
rect 101446 390280 102107 390282
rect 101446 390224 102046 390280
rect 102102 390224 102107 390280
rect 101446 390222 102107 390224
rect 102041 390219 102107 390222
rect 249701 390282 249767 390285
rect 258030 390282 258090 390494
rect 582557 390491 582623 390494
rect 249701 390280 258090 390282
rect 249701 390224 249706 390280
rect 249762 390224 258090 390280
rect 249701 390222 258090 390224
rect 249701 390219 249767 390222
rect 102409 389466 102475 389469
rect 234061 389466 234127 389469
rect 102409 389464 234127 389466
rect 102409 389408 102414 389464
rect 102470 389408 234066 389464
rect 234122 389408 234127 389464
rect 102409 389406 234127 389408
rect 102409 389403 102475 389406
rect 234061 389403 234127 389406
rect 59169 389330 59235 389333
rect 99465 389330 99531 389333
rect 59169 389328 99531 389330
rect 59169 389272 59174 389328
rect 59230 389272 99470 389328
rect 99526 389272 99531 389328
rect 59169 389270 99531 389272
rect 59169 389267 59235 389270
rect 99465 389267 99531 389270
rect 103881 389330 103947 389333
rect 240133 389330 240199 389333
rect 241053 389330 241119 389333
rect 103881 389328 241119 389330
rect 103881 389272 103886 389328
rect 103942 389272 240138 389328
rect 240194 389272 241058 389328
rect 241114 389272 241119 389328
rect 103881 389270 241119 389272
rect 103881 389267 103947 389270
rect 240133 389267 240199 389270
rect 241053 389267 241119 389270
rect 11697 389194 11763 389197
rect 102041 389194 102107 389197
rect 11697 389192 102107 389194
rect 11697 389136 11702 389192
rect 11758 389136 102046 389192
rect 102102 389136 102107 389192
rect 11697 389134 102107 389136
rect 11697 389131 11763 389134
rect 102041 389131 102107 389134
rect 110413 389194 110479 389197
rect 249977 389194 250043 389197
rect 110413 389192 250043 389194
rect 110413 389136 110418 389192
rect 110474 389136 249982 389192
rect 250038 389136 250043 389192
rect 110413 389134 250043 389136
rect 110413 389131 110479 389134
rect 249977 389131 250043 389134
rect 251909 389194 251975 389197
rect 253974 389194 253980 389196
rect 251909 389192 253980 389194
rect 251909 389136 251914 389192
rect 251970 389136 253980 389192
rect 251909 389134 253980 389136
rect 251909 389131 251975 389134
rect 253974 389132 253980 389134
rect 254044 389132 254050 389196
rect 72417 389058 72483 389061
rect 72734 389058 72740 389060
rect 72417 389056 72740 389058
rect 72417 389000 72422 389056
rect 72478 389000 72740 389056
rect 72417 388998 72740 389000
rect 72417 388995 72483 388998
rect 72734 388996 72740 388998
rect 72804 389058 72810 389060
rect 72969 389058 73035 389061
rect 72804 389056 73035 389058
rect 72804 389000 72974 389056
rect 73030 389000 73035 389056
rect 72804 388998 73035 389000
rect 72804 388996 72810 388998
rect 72969 388995 73035 388998
rect 79133 389058 79199 389061
rect 79726 389058 79732 389060
rect 79133 389056 79732 389058
rect 79133 389000 79138 389056
rect 79194 389000 79732 389056
rect 79133 388998 79732 389000
rect 79133 388995 79199 388998
rect 79726 388996 79732 388998
rect 79796 389058 79802 389060
rect 79961 389058 80027 389061
rect 80145 389060 80211 389061
rect 79796 389056 80027 389058
rect 79796 389000 79966 389056
rect 80022 389000 80027 389056
rect 79796 388998 80027 389000
rect 79796 388996 79802 388998
rect 79961 388995 80027 388998
rect 80094 388996 80100 389060
rect 80164 389058 80211 389060
rect 80973 389058 81039 389061
rect 80164 389056 81039 389058
rect 80206 389000 80978 389056
rect 81034 389000 81039 389056
rect 80164 388998 81039 389000
rect 80164 388996 80211 388998
rect 80145 388995 80211 388996
rect 80973 388995 81039 388998
rect 96889 389058 96955 389061
rect 97625 389058 97691 389061
rect 96889 389056 97691 389058
rect 96889 389000 96894 389056
rect 96950 389000 97630 389056
rect 97686 389000 97691 389056
rect 96889 388998 97691 389000
rect 96889 388995 96955 388998
rect 97625 388995 97691 388998
rect 105169 389058 105235 389061
rect 106089 389058 106155 389061
rect 105169 389056 106155 389058
rect 105169 389000 105174 389056
rect 105230 389000 106094 389056
rect 106150 389000 106155 389056
rect 105169 388998 106155 389000
rect 105169 388995 105235 388998
rect 106089 388995 106155 388998
rect 107929 389058 107995 389061
rect 108849 389058 108915 389061
rect 107929 389056 108915 389058
rect 107929 389000 107934 389056
rect 107990 389000 108854 389056
rect 108910 389000 108915 389056
rect 107929 388998 108915 389000
rect 107929 388995 107995 388998
rect 108849 388995 108915 388998
rect 74441 388922 74507 388925
rect 166349 388922 166415 388925
rect 74441 388920 171150 388922
rect 74441 388864 74446 388920
rect 74502 388864 166354 388920
rect 166410 388864 171150 388920
rect 74441 388862 171150 388864
rect 74441 388859 74507 388862
rect 166349 388859 166415 388862
rect 99557 388514 99623 388517
rect 100150 388514 100156 388516
rect 99557 388512 100156 388514
rect 99557 388456 99562 388512
rect 99618 388456 100156 388512
rect 99557 388454 100156 388456
rect 99557 388451 99623 388454
rect 100150 388452 100156 388454
rect 100220 388452 100226 388516
rect 102542 388452 102548 388516
rect 102612 388514 102618 388516
rect 102777 388514 102843 388517
rect 102612 388512 102843 388514
rect 102612 388456 102782 388512
rect 102838 388456 102843 388512
rect 102612 388454 102843 388456
rect 102612 388452 102618 388454
rect 102777 388451 102843 388454
rect 32397 388378 32463 388381
rect 81249 388378 81315 388381
rect 32397 388376 81315 388378
rect 32397 388320 32402 388376
rect 32458 388320 81254 388376
rect 81310 388320 81315 388376
rect 32397 388318 81315 388320
rect 171090 388378 171150 388862
rect 179505 388514 179571 388517
rect 213453 388514 213519 388517
rect 179505 388512 213519 388514
rect 179505 388456 179510 388512
rect 179566 388456 213458 388512
rect 213514 388456 213519 388512
rect 179505 388454 213519 388456
rect 179505 388451 179571 388454
rect 213453 388451 213519 388454
rect 201125 388378 201191 388381
rect 171090 388376 201191 388378
rect 171090 388320 201130 388376
rect 201186 388320 201191 388376
rect 171090 388318 201191 388320
rect 32397 388315 32463 388318
rect 81249 388315 81315 388318
rect 201125 388315 201191 388318
rect 247033 388378 247099 388381
rect 247677 388378 247743 388381
rect 281574 388378 281580 388380
rect 247033 388376 281580 388378
rect 247033 388320 247038 388376
rect 247094 388320 247682 388376
rect 247738 388320 281580 388376
rect 247033 388318 281580 388320
rect 247033 388315 247099 388318
rect 247677 388315 247743 388318
rect 281574 388316 281580 388318
rect 281644 388378 281650 388380
rect 282177 388378 282243 388381
rect 281644 388376 282243 388378
rect 281644 388320 282182 388376
rect 282238 388320 282243 388376
rect 281644 388318 282243 388320
rect 281644 388316 281650 388318
rect 282177 388315 282243 388318
rect 70342 388180 70348 388244
rect 70412 388242 70418 388244
rect 70669 388242 70735 388245
rect 70412 388240 70735 388242
rect 70412 388184 70674 388240
rect 70730 388184 70735 388240
rect 70412 388182 70735 388184
rect 70412 388180 70418 388182
rect 70669 388179 70735 388182
rect 94313 388242 94379 388245
rect 94998 388242 95004 388244
rect 94313 388240 95004 388242
rect 94313 388184 94318 388240
rect 94374 388184 95004 388240
rect 94313 388182 95004 388184
rect 94313 388179 94379 388182
rect 94998 388180 95004 388182
rect 95068 388180 95074 388244
rect 93894 387908 93900 387972
rect 93964 387970 93970 387972
rect 94773 387970 94839 387973
rect 93964 387968 94839 387970
rect 93964 387912 94778 387968
rect 94834 387912 94839 387968
rect 93964 387910 94839 387912
rect 93964 387908 93970 387910
rect 94773 387907 94839 387910
rect 68870 387772 68876 387836
rect 68940 387834 68946 387836
rect 71221 387834 71287 387837
rect 179505 387834 179571 387837
rect 68940 387832 71287 387834
rect 68940 387776 71226 387832
rect 71282 387776 71287 387832
rect 68940 387774 71287 387776
rect 68940 387772 68946 387774
rect 71221 387771 71287 387774
rect 84150 387832 179571 387834
rect 84150 387776 179510 387832
rect 179566 387776 179571 387832
rect 84150 387774 179571 387776
rect 72509 387562 72575 387565
rect 83181 387562 83247 387565
rect 84150 387562 84210 387774
rect 179505 387771 179571 387774
rect 108665 387698 108731 387701
rect 136541 387698 136607 387701
rect 247033 387698 247099 387701
rect 266302 387698 266308 387700
rect 108665 387696 247099 387698
rect 108665 387640 108670 387696
rect 108726 387640 136546 387696
rect 136602 387640 247038 387696
rect 247094 387640 247099 387696
rect 108665 387638 247099 387640
rect 108665 387635 108731 387638
rect 136541 387635 136607 387638
rect 247033 387635 247099 387638
rect 258030 387638 266308 387698
rect 72509 387560 84210 387562
rect 72509 387504 72514 387560
rect 72570 387504 83186 387560
rect 83242 387504 84210 387560
rect 72509 387502 84210 387504
rect 89161 387562 89227 387565
rect 119981 387562 120047 387565
rect 89161 387560 120047 387562
rect 89161 387504 89166 387560
rect 89222 387504 119986 387560
rect 120042 387504 120047 387560
rect 89161 387502 120047 387504
rect 72509 387499 72575 387502
rect 83181 387499 83247 387502
rect 89161 387499 89227 387502
rect 119981 387499 120047 387502
rect 188286 387500 188292 387564
rect 188356 387562 188362 387564
rect 258030 387562 258090 387638
rect 266302 387636 266308 387638
rect 266372 387698 266378 387700
rect 266445 387698 266511 387701
rect 266372 387696 266511 387698
rect 266372 387640 266450 387696
rect 266506 387640 266511 387696
rect 266372 387638 266511 387640
rect 266372 387636 266378 387638
rect 266445 387635 266511 387638
rect 188356 387502 258090 387562
rect 188356 387500 188362 387502
rect 66069 387426 66135 387429
rect 67541 387426 67607 387429
rect 113817 387426 113883 387429
rect 66069 387424 113883 387426
rect 66069 387368 66074 387424
rect 66130 387368 67546 387424
rect 67602 387368 113822 387424
rect 113878 387368 113883 387424
rect 66069 387366 113883 387368
rect 66069 387363 66135 387366
rect 67541 387363 67607 387366
rect 113817 387363 113883 387366
rect 86718 386956 86724 387020
rect 86788 387018 86794 387020
rect 91093 387018 91159 387021
rect 86788 387016 91159 387018
rect 86788 386960 91098 387016
rect 91154 386960 91159 387016
rect 86788 386958 91159 386960
rect 86788 386956 86794 386958
rect 91093 386955 91159 386958
rect 192937 387018 193003 387021
rect 201534 387018 201540 387020
rect 192937 387016 201540 387018
rect 192937 386960 192942 387016
rect 192998 386960 201540 387016
rect 192937 386958 201540 386960
rect 192937 386955 193003 386958
rect 201534 386956 201540 386958
rect 201604 386956 201610 387020
rect 236269 386474 236335 386477
rect 258073 386474 258139 386477
rect 235950 386472 258139 386474
rect 235950 386416 236274 386472
rect 236330 386416 258078 386472
rect 258134 386416 258139 386472
rect 235950 386414 258139 386416
rect 3509 386338 3575 386341
rect 118693 386338 118759 386341
rect 3509 386336 118759 386338
rect 3509 386280 3514 386336
rect 3570 386280 118698 386336
rect 118754 386280 118759 386336
rect 3509 386278 118759 386280
rect 3509 386275 3575 386278
rect 118693 386275 118759 386278
rect 126881 386338 126947 386341
rect 235950 386338 236010 386414
rect 236269 386411 236335 386414
rect 258073 386411 258139 386414
rect 263542 386338 263548 386340
rect 126881 386336 236010 386338
rect 126881 386280 126886 386336
rect 126942 386280 236010 386336
rect 126881 386278 236010 386280
rect 258030 386278 263548 386338
rect 126881 386275 126947 386278
rect 187049 386202 187115 386205
rect 258030 386202 258090 386278
rect 263542 386276 263548 386278
rect 263612 386338 263618 386340
rect 263777 386338 263843 386341
rect 285673 386340 285739 386341
rect 285622 386338 285628 386340
rect 263612 386336 263843 386338
rect 263612 386280 263782 386336
rect 263838 386280 263843 386336
rect 263612 386278 263843 386280
rect 285582 386278 285628 386338
rect 285692 386336 285739 386340
rect 285734 386280 285739 386336
rect 263612 386276 263618 386278
rect 263777 386275 263843 386278
rect 285622 386276 285628 386278
rect 285692 386276 285739 386280
rect 285673 386275 285739 386276
rect 187049 386200 258090 386202
rect 187049 386144 187054 386200
rect 187110 386144 258090 386200
rect 187049 386142 258090 386144
rect 187049 386139 187115 386142
rect 104801 385658 104867 385661
rect 117313 385658 117379 385661
rect 104801 385656 117379 385658
rect 104801 385600 104806 385656
rect 104862 385600 117318 385656
rect 117374 385600 117379 385656
rect 104801 385598 117379 385600
rect 104801 385595 104867 385598
rect 117313 385595 117379 385598
rect 192845 385658 192911 385661
rect 208342 385658 208348 385660
rect 192845 385656 208348 385658
rect 192845 385600 192850 385656
rect 192906 385600 208348 385656
rect 192845 385598 208348 385600
rect 192845 385595 192911 385598
rect 208342 385596 208348 385598
rect 208412 385596 208418 385660
rect 208485 385658 208551 385661
rect 285622 385658 285628 385660
rect 208485 385656 285628 385658
rect 208485 385600 208490 385656
rect 208546 385600 285628 385656
rect 208485 385598 285628 385600
rect 208485 385595 208551 385598
rect 285622 385596 285628 385598
rect 285692 385596 285698 385660
rect 77201 384978 77267 384981
rect 129089 384978 129155 384981
rect 77201 384976 129155 384978
rect 77201 384920 77206 384976
rect 77262 384920 129094 384976
rect 129150 384920 129155 384976
rect 77201 384918 129155 384920
rect 77201 384915 77267 384918
rect 129089 384915 129155 384918
rect 173249 384978 173315 384981
rect 173801 384978 173867 384981
rect 207749 384978 207815 384981
rect 173249 384976 207815 384978
rect 173249 384920 173254 384976
rect 173310 384920 173806 384976
rect 173862 384920 207754 384976
rect 207810 384920 207815 384976
rect 173249 384918 207815 384920
rect 173249 384915 173315 384918
rect 173801 384915 173867 384918
rect 207749 384915 207815 384918
rect -960 384284 480 384524
rect 238109 384434 238175 384437
rect 244406 384434 244412 384436
rect 238109 384432 244412 384434
rect 238109 384376 238114 384432
rect 238170 384376 244412 384432
rect 238109 384374 244412 384376
rect 238109 384371 238175 384374
rect 244406 384372 244412 384374
rect 244476 384372 244482 384436
rect 66662 384236 66668 384300
rect 66732 384298 66738 384300
rect 88977 384298 89043 384301
rect 66732 384296 89043 384298
rect 66732 384240 88982 384296
rect 89038 384240 89043 384296
rect 66732 384238 89043 384240
rect 66732 384236 66738 384238
rect 88977 384235 89043 384238
rect 101489 384298 101555 384301
rect 113449 384298 113515 384301
rect 101489 384296 113515 384298
rect 101489 384240 101494 384296
rect 101550 384240 113454 384296
rect 113510 384240 113515 384296
rect 101489 384238 113515 384240
rect 101489 384235 101555 384238
rect 113449 384235 113515 384238
rect 233877 384298 233943 384301
rect 242934 384298 242940 384300
rect 233877 384296 242940 384298
rect 233877 384240 233882 384296
rect 233938 384240 242940 384296
rect 233877 384238 242940 384240
rect 233877 384235 233943 384238
rect 242934 384236 242940 384238
rect 243004 384236 243010 384300
rect 216397 384028 216463 384029
rect 216397 384024 216444 384028
rect 216508 384026 216514 384028
rect 216397 383968 216402 384024
rect 216397 383964 216444 383968
rect 216508 383966 216554 384026
rect 216508 383964 216514 383966
rect 216397 383963 216463 383964
rect 197353 383890 197419 383893
rect 582465 383890 582531 383893
rect 197353 383888 582531 383890
rect 197353 383832 197358 383888
rect 197414 383832 582470 383888
rect 582526 383832 582531 383888
rect 197353 383830 582531 383832
rect 197353 383827 197419 383830
rect 582465 383827 582531 383830
rect 69657 383754 69723 383757
rect 74574 383754 74580 383756
rect 69657 383752 74580 383754
rect 69657 383696 69662 383752
rect 69718 383696 74580 383752
rect 69657 383694 74580 383696
rect 69657 383691 69723 383694
rect 74574 383692 74580 383694
rect 74644 383692 74650 383756
rect 91001 383754 91067 383757
rect 96286 383754 96292 383756
rect 91001 383752 96292 383754
rect 91001 383696 91006 383752
rect 91062 383696 96292 383752
rect 91001 383694 96292 383696
rect 91001 383691 91067 383694
rect 96286 383692 96292 383694
rect 96356 383692 96362 383756
rect 105905 383618 105971 383621
rect 242985 383618 243051 383621
rect 243997 383618 244063 383621
rect 105905 383616 244063 383618
rect 105905 383560 105910 383616
rect 105966 383560 242990 383616
rect 243046 383560 244002 383616
rect 244058 383560 244063 383616
rect 105905 383558 244063 383560
rect 105905 383555 105971 383558
rect 242985 383555 243051 383558
rect 243997 383555 244063 383558
rect 81341 382938 81407 382941
rect 87454 382938 87460 382940
rect 81341 382936 87460 382938
rect 81341 382880 81346 382936
rect 81402 382880 87460 382936
rect 81341 382878 87460 382880
rect 81341 382875 81407 382878
rect 87454 382876 87460 382878
rect 87524 382876 87530 382940
rect 105997 382938 106063 382941
rect 114686 382938 114692 382940
rect 105997 382936 114692 382938
rect 105997 382880 106002 382936
rect 106058 382880 114692 382936
rect 105997 382878 114692 382880
rect 105997 382875 106063 382878
rect 114686 382876 114692 382878
rect 114756 382876 114762 382940
rect 190085 382938 190151 382941
rect 282913 382938 282979 382941
rect 190085 382936 282979 382938
rect 190085 382880 190090 382936
rect 190146 382880 282918 382936
rect 282974 382880 282979 382936
rect 190085 382878 282979 382880
rect 190085 382875 190151 382878
rect 282913 382875 282979 382878
rect 188521 382394 188587 382397
rect 190085 382394 190151 382397
rect 188521 382392 190151 382394
rect 188521 382336 188526 382392
rect 188582 382336 190090 382392
rect 190146 382336 190151 382392
rect 188521 382334 190151 382336
rect 188521 382331 188587 382334
rect 190085 382331 190151 382334
rect 119337 382258 119403 382261
rect 258349 382258 258415 382261
rect 119337 382256 258415 382258
rect 119337 382200 119342 382256
rect 119398 382200 258354 382256
rect 258410 382200 258415 382256
rect 119337 382198 258415 382200
rect 119337 382195 119403 382198
rect 258349 382195 258415 382198
rect 168373 381714 168439 381717
rect 197353 381714 197419 381717
rect 168373 381712 197419 381714
rect 168373 381656 168378 381712
rect 168434 381656 197358 381712
rect 197414 381656 197419 381712
rect 168373 381654 197419 381656
rect 168373 381651 168439 381654
rect 197353 381651 197419 381654
rect 89529 381578 89595 381581
rect 189073 381578 189139 381581
rect 89529 381576 189139 381578
rect 89529 381520 89534 381576
rect 89590 381520 189078 381576
rect 189134 381520 189139 381576
rect 89529 381518 189139 381520
rect 89529 381515 89595 381518
rect 189073 381515 189139 381518
rect 69606 380836 69612 380900
rect 69676 380898 69682 380900
rect 127617 380898 127683 380901
rect 69676 380896 127683 380898
rect 69676 380840 127622 380896
rect 127678 380840 127683 380896
rect 69676 380838 127683 380840
rect 69676 380836 69682 380838
rect 127617 380835 127683 380838
rect 144177 380898 144243 380901
rect 276197 380898 276263 380901
rect 144177 380896 276263 380898
rect 144177 380840 144182 380896
rect 144238 380840 276202 380896
rect 276258 380840 276263 380896
rect 144177 380838 276263 380840
rect 144177 380835 144243 380838
rect 276197 380835 276263 380838
rect 106457 380762 106523 380765
rect 124305 380762 124371 380765
rect 124857 380762 124923 380765
rect 106457 380760 124923 380762
rect 106457 380704 106462 380760
rect 106518 380704 124310 380760
rect 124366 380704 124862 380760
rect 124918 380704 124923 380760
rect 106457 380702 124923 380704
rect 106457 380699 106523 380702
rect 124305 380699 124371 380702
rect 124857 380699 124923 380702
rect 192702 380156 192708 380220
rect 192772 380218 192778 380220
rect 244365 380218 244431 380221
rect 192772 380216 244431 380218
rect 192772 380160 244370 380216
rect 244426 380160 244431 380216
rect 192772 380158 244431 380160
rect 192772 380156 192778 380158
rect 244365 380155 244431 380158
rect 276197 379540 276263 379541
rect 276197 379538 276244 379540
rect 276152 379536 276244 379538
rect 276152 379480 276202 379536
rect 276152 379478 276244 379480
rect 276197 379476 276244 379478
rect 276308 379476 276314 379540
rect 276197 379475 276263 379476
rect 109033 379402 109099 379405
rect 109677 379402 109743 379405
rect 124397 379402 124463 379405
rect 248689 379402 248755 379405
rect 249057 379402 249123 379405
rect 109033 379400 249123 379402
rect 109033 379344 109038 379400
rect 109094 379344 109682 379400
rect 109738 379344 124402 379400
rect 124458 379344 248694 379400
rect 248750 379344 249062 379400
rect 249118 379344 249123 379400
rect 109033 379342 249123 379344
rect 109033 379339 109099 379342
rect 109677 379339 109743 379342
rect 124397 379339 124463 379342
rect 248689 379339 248755 379342
rect 249057 379339 249123 379342
rect 582465 378450 582531 378453
rect 583520 378450 584960 378540
rect 582465 378448 584960 378450
rect 582465 378392 582470 378448
rect 582526 378392 584960 378448
rect 582465 378390 584960 378392
rect 582465 378387 582531 378390
rect 583520 378300 584960 378390
rect 242750 377980 242756 378044
rect 242820 378042 242826 378044
rect 249977 378042 250043 378045
rect 242820 378040 250043 378042
rect 242820 377984 249982 378040
rect 250038 377984 250043 378040
rect 242820 377982 250043 377984
rect 242820 377980 242826 377982
rect 249977 377979 250043 377982
rect 166257 377362 166323 377365
rect 256693 377362 256759 377365
rect 166257 377360 256759 377362
rect 166257 377304 166262 377360
rect 166318 377304 256698 377360
rect 256754 377304 256759 377360
rect 166257 377302 256759 377304
rect 166257 377299 166323 377302
rect 256693 377299 256759 377302
rect 67766 376620 67772 376684
rect 67836 376682 67842 376684
rect 158713 376682 158779 376685
rect 159449 376682 159515 376685
rect 67836 376680 159515 376682
rect 67836 376624 158718 376680
rect 158774 376624 159454 376680
rect 159510 376624 159515 376680
rect 67836 376622 159515 376624
rect 67836 376620 67842 376622
rect 158713 376619 158779 376622
rect 159449 376619 159515 376622
rect 204253 376682 204319 376685
rect 205541 376682 205607 376685
rect 582373 376682 582439 376685
rect 204253 376680 582439 376682
rect 204253 376624 204258 376680
rect 204314 376624 205546 376680
rect 205602 376624 582378 376680
rect 582434 376624 582439 376680
rect 204253 376622 582439 376624
rect 204253 376619 204319 376622
rect 205541 376619 205607 376622
rect 582373 376619 582439 376622
rect 155217 376546 155283 376549
rect 260925 376546 260991 376549
rect 261477 376546 261543 376549
rect 155217 376544 261543 376546
rect 155217 376488 155222 376544
rect 155278 376488 260930 376544
rect 260986 376488 261482 376544
rect 261538 376488 261543 376544
rect 155217 376486 261543 376488
rect 155217 376483 155283 376486
rect 260925 376483 260991 376486
rect 261477 376483 261543 376486
rect 197118 375940 197124 376004
rect 197188 376002 197194 376004
rect 203006 376002 203012 376004
rect 197188 375942 203012 376002
rect 197188 375940 197194 375942
rect 203006 375940 203012 375942
rect 203076 375940 203082 376004
rect 169017 375322 169083 375325
rect 258257 375322 258323 375325
rect 258390 375322 258396 375324
rect 169017 375320 258396 375322
rect 169017 375264 169022 375320
rect 169078 375264 258262 375320
rect 258318 375264 258396 375320
rect 169017 375262 258396 375264
rect 169017 375259 169083 375262
rect 258257 375259 258323 375262
rect 258390 375260 258396 375262
rect 258460 375260 258466 375324
rect 65885 373962 65951 373965
rect 188521 373962 188587 373965
rect 65885 373960 188587 373962
rect 65885 373904 65890 373960
rect 65946 373904 188526 373960
rect 188582 373904 188587 373960
rect 65885 373902 188587 373904
rect 65885 373899 65951 373902
rect 188521 373899 188587 373902
rect 67173 372602 67239 372605
rect 160686 372602 160692 372604
rect 67173 372600 160692 372602
rect 67173 372544 67178 372600
rect 67234 372544 160692 372600
rect 67173 372542 160692 372544
rect 67173 372539 67239 372542
rect 160686 372540 160692 372542
rect 160756 372540 160762 372604
rect 117221 371922 117287 371925
rect 212533 371922 212599 371925
rect 117221 371920 212599 371922
rect 117221 371864 117226 371920
rect 117282 371864 212538 371920
rect 212594 371864 212599 371920
rect 117221 371862 212599 371864
rect 117221 371859 117287 371862
rect 212533 371859 212599 371862
rect -960 371378 480 371468
rect 3417 371378 3483 371381
rect -960 371376 3483 371378
rect -960 371320 3422 371376
rect 3478 371320 3483 371376
rect -960 371318 3483 371320
rect -960 371228 480 371318
rect 3417 371315 3483 371318
rect 236494 370636 236500 370700
rect 236564 370698 236570 370700
rect 247718 370698 247724 370700
rect 236564 370638 247724 370698
rect 236564 370636 236570 370638
rect 247718 370636 247724 370638
rect 247788 370636 247794 370700
rect 126329 370562 126395 370565
rect 237373 370562 237439 370565
rect 126329 370560 237439 370562
rect 126329 370504 126334 370560
rect 126390 370504 237378 370560
rect 237434 370504 237439 370560
rect 126329 370502 237439 370504
rect 126329 370499 126395 370502
rect 237373 370499 237439 370502
rect 237373 369882 237439 369885
rect 238017 369882 238083 369885
rect 237373 369880 238083 369882
rect 237373 369824 237378 369880
rect 237434 369824 238022 369880
rect 238078 369824 238083 369880
rect 237373 369822 238083 369824
rect 237373 369819 237439 369822
rect 238017 369819 238083 369822
rect 83457 369746 83523 369749
rect 180149 369746 180215 369749
rect 83457 369744 180215 369746
rect 83457 369688 83462 369744
rect 83518 369688 180154 369744
rect 180210 369688 180215 369744
rect 83457 369686 180215 369688
rect 83457 369683 83523 369686
rect 180149 369683 180215 369686
rect 79961 368386 80027 368389
rect 173249 368386 173315 368389
rect 79961 368384 173315 368386
rect 79961 368328 79966 368384
rect 80022 368328 173254 368384
rect 173310 368328 173315 368384
rect 79961 368326 173315 368328
rect 79961 368323 80027 368326
rect 173249 368323 173315 368326
rect 252553 368386 252619 368389
rect 252686 368386 252692 368388
rect 252553 368384 252692 368386
rect 252553 368328 252558 368384
rect 252614 368328 252692 368384
rect 252553 368326 252692 368328
rect 252553 368323 252619 368326
rect 252686 368324 252692 368326
rect 252756 368324 252762 368388
rect 208485 367706 208551 367709
rect 284569 367706 284635 367709
rect 208485 367704 284635 367706
rect 208485 367648 208490 367704
rect 208546 367648 284574 367704
rect 284630 367648 284635 367704
rect 208485 367646 284635 367648
rect 208485 367643 208551 367646
rect 284569 367643 284635 367646
rect 189073 367162 189139 367165
rect 190177 367162 190243 367165
rect 198089 367162 198155 367165
rect 189073 367160 198155 367162
rect 189073 367104 189078 367160
rect 189134 367104 190182 367160
rect 190238 367104 198094 367160
rect 198150 367104 198155 367160
rect 189073 367102 198155 367104
rect 189073 367099 189139 367102
rect 190177 367099 190243 367102
rect 198089 367099 198155 367102
rect 122097 367026 122163 367029
rect 289813 367026 289879 367029
rect 122097 367024 289879 367026
rect 122097 366968 122102 367024
rect 122158 366968 289818 367024
rect 289874 366968 289879 367024
rect 122097 366966 289879 366968
rect 122097 366963 122163 366966
rect 289813 366963 289879 366966
rect 218646 366284 218652 366348
rect 218716 366346 218722 366348
rect 249742 366346 249748 366348
rect 218716 366286 249748 366346
rect 218716 366284 218722 366286
rect 249742 366284 249748 366286
rect 249812 366284 249818 366348
rect 582373 365122 582439 365125
rect 583520 365122 584960 365212
rect 582373 365120 584960 365122
rect 582373 365064 582378 365120
rect 582434 365064 584960 365120
rect 582373 365062 584960 365064
rect 582373 365059 582439 365062
rect 120717 364986 120783 364989
rect 170489 364986 170555 364989
rect 120717 364984 170555 364986
rect 120717 364928 120722 364984
rect 120778 364928 170494 364984
rect 170550 364928 170555 364984
rect 120717 364926 170555 364928
rect 120717 364923 120783 364926
rect 170489 364923 170555 364926
rect 215150 364924 215156 364988
rect 215220 364986 215226 364988
rect 253933 364986 253999 364989
rect 215220 364984 253999 364986
rect 215220 364928 253938 364984
rect 253994 364928 253999 364984
rect 583520 364972 584960 365062
rect 215220 364926 253999 364928
rect 215220 364924 215226 364926
rect 253933 364923 253999 364926
rect 193121 363626 193187 363629
rect 245745 363626 245811 363629
rect 193121 363624 245811 363626
rect 193121 363568 193126 363624
rect 193182 363568 245750 363624
rect 245806 363568 245811 363624
rect 193121 363566 245811 363568
rect 193121 363563 193187 363566
rect 245745 363563 245811 363566
rect 261477 363082 261543 363085
rect 269246 363082 269252 363084
rect 261477 363080 269252 363082
rect 261477 363024 261482 363080
rect 261538 363024 269252 363080
rect 261477 363022 269252 363024
rect 261477 363019 261543 363022
rect 269246 363020 269252 363022
rect 269316 363020 269322 363084
rect 187693 361586 187759 361589
rect 188981 361586 189047 361589
rect 219433 361586 219499 361589
rect 187693 361584 219499 361586
rect 187693 361528 187698 361584
rect 187754 361528 188986 361584
rect 189042 361528 219438 361584
rect 219494 361528 219499 361584
rect 187693 361526 219499 361528
rect 187693 361523 187759 361526
rect 188981 361523 189047 361526
rect 219433 361523 219499 361526
rect 221222 360844 221228 360908
rect 221292 360906 221298 360908
rect 251265 360906 251331 360909
rect 221292 360904 251331 360906
rect 221292 360848 251270 360904
rect 251326 360848 251331 360904
rect 221292 360846 251331 360848
rect 221292 360844 221298 360846
rect 251265 360843 251331 360846
rect -960 358458 480 358548
rect 3233 358458 3299 358461
rect -960 358456 3299 358458
rect -960 358400 3238 358456
rect 3294 358400 3299 358456
rect -960 358398 3299 358400
rect -960 358308 480 358398
rect 3233 358395 3299 358398
rect 56409 358050 56475 358053
rect 193806 358050 193812 358052
rect 56409 358048 193812 358050
rect 56409 357992 56414 358048
rect 56470 357992 193812 358048
rect 56409 357990 193812 357992
rect 56409 357987 56475 357990
rect 193806 357988 193812 357990
rect 193876 357988 193882 358052
rect 232589 358050 232655 358053
rect 267958 358050 267964 358052
rect 232589 358048 267964 358050
rect 232589 357992 232594 358048
rect 232650 357992 267964 358048
rect 232589 357990 267964 357992
rect 232589 357987 232655 357990
rect 267958 357988 267964 357990
rect 268028 357988 268034 358052
rect 72734 356628 72740 356692
rect 72804 356690 72810 356692
rect 73061 356690 73127 356693
rect 200113 356690 200179 356693
rect 72804 356688 200179 356690
rect 72804 356632 73066 356688
rect 73122 356632 200118 356688
rect 200174 356632 200179 356688
rect 72804 356630 200179 356632
rect 72804 356628 72810 356630
rect 73061 356627 73127 356630
rect 200113 356627 200179 356630
rect 195973 356010 196039 356013
rect 196617 356010 196683 356013
rect 195973 356008 196683 356010
rect 195973 355952 195978 356008
rect 196034 355952 196622 356008
rect 196678 355952 196683 356008
rect 195973 355950 196683 355952
rect 195973 355947 196039 355950
rect 196617 355947 196683 355950
rect 188838 355404 188844 355468
rect 188908 355466 188914 355468
rect 231117 355466 231183 355469
rect 188908 355464 231183 355466
rect 188908 355408 231122 355464
rect 231178 355408 231183 355464
rect 188908 355406 231183 355408
rect 188908 355404 188914 355406
rect 231117 355403 231183 355406
rect 68870 355268 68876 355332
rect 68940 355330 68946 355332
rect 196617 355330 196683 355333
rect 68940 355328 196683 355330
rect 68940 355272 196622 355328
rect 196678 355272 196683 355328
rect 68940 355270 196683 355272
rect 68940 355268 68946 355270
rect 196617 355267 196683 355270
rect 193489 353970 193555 353973
rect 244273 353970 244339 353973
rect 193489 353968 244339 353970
rect 193489 353912 193494 353968
rect 193550 353912 244278 353968
rect 244334 353912 244339 353968
rect 193489 353910 244339 353912
rect 193489 353907 193555 353910
rect 244273 353907 244339 353910
rect 582649 351930 582715 351933
rect 583520 351930 584960 352020
rect 582649 351928 584960 351930
rect 582649 351872 582654 351928
rect 582710 351872 584960 351928
rect 582649 351870 584960 351872
rect 582649 351867 582715 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 3417 345402 3483 345405
rect -960 345400 3483 345402
rect -960 345344 3422 345400
rect 3478 345344 3483 345400
rect -960 345342 3483 345344
rect -960 345252 480 345342
rect 3417 345339 3483 345342
rect 266445 339556 266511 339557
rect 266445 339554 266492 339556
rect 266400 339552 266492 339554
rect 266400 339496 266450 339552
rect 266400 339494 266492 339496
rect 266445 339492 266492 339494
rect 266556 339492 266562 339556
rect 266445 339491 266511 339492
rect 193806 338676 193812 338740
rect 193876 338738 193882 338740
rect 228357 338738 228423 338741
rect 193876 338736 228423 338738
rect 193876 338680 228362 338736
rect 228418 338680 228423 338736
rect 193876 338678 228423 338680
rect 193876 338676 193882 338678
rect 228357 338675 228423 338678
rect 583520 338452 584960 338692
rect 72417 338194 72483 338197
rect 72550 338194 72556 338196
rect 72417 338192 72556 338194
rect 72417 338136 72422 338192
rect 72478 338136 72556 338192
rect 72417 338134 72556 338136
rect 72417 338131 72483 338134
rect 72550 338132 72556 338134
rect 72620 338194 72626 338196
rect 73061 338194 73127 338197
rect 72620 338192 73127 338194
rect 72620 338136 73066 338192
rect 73122 338136 73127 338192
rect 72620 338134 73127 338136
rect 72620 338132 72626 338134
rect 73061 338131 73127 338134
rect 252553 338060 252619 338061
rect 252502 337996 252508 338060
rect 252572 338058 252619 338060
rect 252572 338056 252664 338058
rect 252614 338000 252664 338056
rect 252572 337998 252664 338000
rect 252572 337996 252619 337998
rect 252553 337995 252619 337996
rect 208393 337378 208459 337381
rect 238886 337378 238892 337380
rect 208393 337376 238892 337378
rect 208393 337320 208398 337376
rect 208454 337320 238892 337376
rect 208393 337318 238892 337320
rect 208393 337315 208459 337318
rect 238886 337316 238892 337318
rect 238956 337316 238962 337380
rect 249701 336698 249767 336701
rect 252686 336698 252692 336700
rect 249701 336696 252692 336698
rect 249701 336640 249706 336696
rect 249762 336640 252692 336696
rect 249701 336638 252692 336640
rect 249701 336635 249767 336638
rect 252686 336636 252692 336638
rect 252756 336636 252762 336700
rect 213913 334658 213979 334661
rect 252502 334658 252508 334660
rect 213913 334656 252508 334658
rect 213913 334600 213918 334656
rect 213974 334600 252508 334656
rect 213913 334598 252508 334600
rect 213913 334595 213979 334598
rect 252502 334596 252508 334598
rect 252572 334596 252578 334660
rect 159357 332618 159423 332621
rect 262438 332618 262444 332620
rect 159357 332616 262444 332618
rect 159357 332560 159362 332616
rect 159418 332560 262444 332616
rect 159357 332558 262444 332560
rect 159357 332555 159423 332558
rect 262438 332556 262444 332558
rect 262508 332556 262514 332620
rect -960 332196 480 332436
rect 211797 331802 211863 331805
rect 260966 331802 260972 331804
rect 211797 331800 260972 331802
rect 211797 331744 211802 331800
rect 211858 331744 260972 331800
rect 211797 331742 260972 331744
rect 211797 331739 211863 331742
rect 260966 331740 260972 331742
rect 261036 331740 261042 331804
rect 146937 331258 147003 331261
rect 227805 331258 227871 331261
rect 146937 331256 227871 331258
rect 146937 331200 146942 331256
rect 146998 331200 227810 331256
rect 227866 331200 227871 331256
rect 146937 331198 227871 331200
rect 146937 331195 147003 331198
rect 227805 331195 227871 331198
rect 174721 329898 174787 329901
rect 244365 329898 244431 329901
rect 174721 329896 244431 329898
rect 174721 329840 174726 329896
rect 174782 329840 244370 329896
rect 244426 329840 244431 329896
rect 174721 329838 244431 329840
rect 174721 329835 174787 329838
rect 244365 329835 244431 329838
rect 135897 328538 135963 328541
rect 208393 328538 208459 328541
rect 135897 328536 208459 328538
rect 135897 328480 135902 328536
rect 135958 328480 208398 328536
rect 208454 328480 208459 328536
rect 135897 328478 208459 328480
rect 135897 328475 135963 328478
rect 208393 328475 208459 328478
rect 252318 328340 252324 328404
rect 252388 328402 252394 328404
rect 255497 328402 255563 328405
rect 252388 328400 255563 328402
rect 252388 328344 255502 328400
rect 255558 328344 255563 328400
rect 252388 328342 255563 328344
rect 252388 328340 252394 328342
rect 255497 328339 255563 328342
rect 155401 327178 155467 327181
rect 252318 327178 252324 327180
rect 155401 327176 252324 327178
rect 155401 327120 155406 327176
rect 155462 327120 252324 327176
rect 155401 327118 252324 327120
rect 155401 327115 155467 327118
rect 252318 327116 252324 327118
rect 252388 327116 252394 327180
rect 73061 326362 73127 326365
rect 77334 326362 77340 326364
rect 73061 326360 77340 326362
rect 73061 326304 73066 326360
rect 73122 326304 77340 326360
rect 73061 326302 77340 326304
rect 73061 326299 73127 326302
rect 77334 326300 77340 326302
rect 77404 326300 77410 326364
rect 137461 326362 137527 326365
rect 223481 326362 223547 326365
rect 137461 326360 223547 326362
rect 137461 326304 137466 326360
rect 137522 326304 223486 326360
rect 223542 326304 223547 326360
rect 137461 326302 223547 326304
rect 137461 326299 137527 326302
rect 223481 326299 223547 326302
rect 215937 325818 216003 325821
rect 256785 325818 256851 325821
rect 215937 325816 256851 325818
rect 215937 325760 215942 325816
rect 215998 325760 256790 325816
rect 256846 325760 256851 325816
rect 215937 325758 256851 325760
rect 215937 325755 216003 325758
rect 256785 325755 256851 325758
rect 580257 325274 580323 325277
rect 583520 325274 584960 325364
rect 580257 325272 584960 325274
rect 580257 325216 580262 325272
rect 580318 325216 584960 325272
rect 580257 325214 584960 325216
rect 580257 325211 580323 325214
rect 583520 325124 584960 325214
rect 22001 324458 22067 324461
rect 202321 324458 202387 324461
rect 22001 324456 202387 324458
rect 22001 324400 22006 324456
rect 22062 324400 202326 324456
rect 202382 324400 202387 324456
rect 22001 324398 202387 324400
rect 22001 324395 22067 324398
rect 202321 324395 202387 324398
rect 97901 323642 97967 323645
rect 110638 323642 110644 323644
rect 97901 323640 110644 323642
rect 97901 323584 97906 323640
rect 97962 323584 110644 323640
rect 97901 323582 110644 323584
rect 97901 323579 97967 323582
rect 110638 323580 110644 323582
rect 110708 323580 110714 323644
rect 198733 323098 198799 323101
rect 199326 323098 199332 323100
rect 198733 323096 199332 323098
rect 198733 323040 198738 323096
rect 198794 323040 199332 323096
rect 198733 323038 199332 323040
rect 198733 323035 198799 323038
rect 199326 323036 199332 323038
rect 199396 323036 199402 323100
rect 167637 322962 167703 322965
rect 168281 322962 168347 322965
rect 217174 322962 217180 322964
rect 167637 322960 217180 322962
rect 167637 322904 167642 322960
rect 167698 322904 168286 322960
rect 168342 322904 217180 322960
rect 167637 322902 217180 322904
rect 167637 322899 167703 322902
rect 168281 322899 168347 322902
rect 217174 322900 217180 322902
rect 217244 322900 217250 322964
rect 66478 322084 66484 322148
rect 66548 322146 66554 322148
rect 161933 322146 161999 322149
rect 66548 322144 161999 322146
rect 66548 322088 161938 322144
rect 161994 322088 161999 322144
rect 66548 322086 161999 322088
rect 66548 322084 66554 322086
rect 161933 322083 161999 322086
rect 249609 321738 249675 321741
rect 252553 321738 252619 321741
rect 249609 321736 252619 321738
rect 249609 321680 249614 321736
rect 249670 321680 252558 321736
rect 252614 321680 252619 321736
rect 249609 321678 252619 321680
rect 249609 321675 249675 321678
rect 252553 321675 252619 321678
rect 159541 321602 159607 321605
rect 270585 321602 270651 321605
rect 159541 321600 270651 321602
rect 159541 321544 159546 321600
rect 159602 321544 270590 321600
rect 270646 321544 270651 321600
rect 159541 321542 270651 321544
rect 159541 321539 159607 321542
rect 270585 321539 270651 321542
rect 86861 320786 86927 320789
rect 94446 320786 94452 320788
rect 86861 320784 94452 320786
rect 86861 320728 86866 320784
rect 86922 320728 94452 320784
rect 86861 320726 94452 320728
rect 86861 320723 86927 320726
rect 94446 320724 94452 320726
rect 94516 320724 94522 320788
rect 111057 320786 111123 320789
rect 116025 320786 116091 320789
rect 111057 320784 116091 320786
rect 111057 320728 111062 320784
rect 111118 320728 116030 320784
rect 116086 320728 116091 320784
rect 111057 320726 116091 320728
rect 111057 320723 111123 320726
rect 116025 320723 116091 320726
rect 271873 320650 271939 320653
rect 272149 320650 272215 320653
rect 271873 320648 272215 320650
rect 271873 320592 271878 320648
rect 271934 320592 272154 320648
rect 272210 320592 272215 320648
rect 271873 320590 272215 320592
rect 271873 320587 271939 320590
rect 272149 320587 272215 320590
rect 77385 320242 77451 320245
rect 77385 320240 84210 320242
rect 77385 320184 77390 320240
rect 77446 320184 84210 320240
rect 77385 320182 84210 320184
rect 77385 320179 77451 320182
rect 84150 320106 84210 320182
rect 85798 320180 85804 320244
rect 85868 320180 85874 320244
rect 95141 320242 95207 320245
rect 100753 320242 100819 320245
rect 95141 320240 100819 320242
rect 95141 320184 95146 320240
rect 95202 320184 100758 320240
rect 100814 320184 100819 320240
rect 95141 320182 100819 320184
rect 85806 320106 85866 320180
rect 95141 320179 95207 320182
rect 100753 320179 100819 320182
rect 102685 320244 102751 320245
rect 102685 320240 102732 320244
rect 102796 320242 102802 320244
rect 129089 320242 129155 320245
rect 272149 320242 272215 320245
rect 102685 320184 102690 320240
rect 102685 320180 102732 320184
rect 102796 320182 102842 320242
rect 129089 320240 272215 320242
rect 129089 320184 129094 320240
rect 129150 320184 272154 320240
rect 272210 320184 272215 320240
rect 129089 320182 272215 320184
rect 102796 320180 102802 320182
rect 102685 320179 102751 320180
rect 129089 320179 129155 320182
rect 272149 320179 272215 320182
rect 184933 320106 184999 320109
rect 185669 320106 185735 320109
rect 84150 320104 185735 320106
rect 84150 320048 184938 320104
rect 184994 320048 185674 320104
rect 185730 320048 185735 320104
rect 84150 320046 185735 320048
rect 184933 320043 184999 320046
rect 185669 320043 185735 320046
rect 263593 320106 263659 320109
rect 263777 320106 263843 320109
rect 263593 320104 263843 320106
rect 263593 320048 263598 320104
rect 263654 320048 263782 320104
rect 263838 320048 263843 320104
rect 263593 320046 263843 320048
rect 263593 320043 263659 320046
rect 263777 320043 263843 320046
rect 90909 319426 90975 319429
rect 98126 319426 98132 319428
rect 90909 319424 98132 319426
rect -960 319290 480 319380
rect 90909 319368 90914 319424
rect 90970 319368 98132 319424
rect 90909 319366 98132 319368
rect 90909 319363 90975 319366
rect 98126 319364 98132 319366
rect 98196 319364 98202 319428
rect 99281 319426 99347 319429
rect 111742 319426 111748 319428
rect 99281 319424 111748 319426
rect 99281 319368 99286 319424
rect 99342 319368 111748 319424
rect 99281 319366 111748 319368
rect 99281 319363 99347 319366
rect 111742 319364 111748 319366
rect 111812 319364 111818 319428
rect 4061 319290 4127 319293
rect -960 319288 4127 319290
rect -960 319232 4066 319288
rect 4122 319232 4127 319288
rect -960 319230 4127 319232
rect -960 319140 480 319230
rect 4061 319227 4127 319230
rect 188613 319018 188679 319021
rect 263777 319018 263843 319021
rect 188613 319016 263843 319018
rect 188613 318960 188618 319016
rect 188674 318960 263782 319016
rect 263838 318960 263843 319016
rect 188613 318958 263843 318960
rect 188613 318955 188679 318958
rect 263777 318955 263843 318958
rect 163497 318882 163563 318885
rect 263685 318882 263751 318885
rect 163497 318880 263751 318882
rect 163497 318824 163502 318880
rect 163558 318824 263690 318880
rect 263746 318824 263751 318880
rect 163497 318822 263751 318824
rect 163497 318819 163563 318822
rect 263685 318819 263751 318822
rect 84694 318684 84700 318748
rect 84764 318746 84770 318748
rect 84837 318746 84903 318749
rect 183461 318746 183527 318749
rect 84764 318744 183527 318746
rect 84764 318688 84842 318744
rect 84898 318688 183466 318744
rect 183522 318688 183527 318744
rect 84764 318686 183527 318688
rect 84764 318684 84770 318686
rect 84837 318683 84903 318686
rect 183461 318683 183527 318686
rect 95049 318066 95115 318069
rect 106406 318066 106412 318068
rect 95049 318064 106412 318066
rect 95049 318008 95054 318064
rect 95110 318008 106412 318064
rect 95049 318006 106412 318008
rect 95049 318003 95115 318006
rect 106406 318004 106412 318006
rect 106476 318004 106482 318068
rect 183461 318066 183527 318069
rect 216213 318066 216279 318069
rect 183461 318064 216279 318066
rect 183461 318008 183466 318064
rect 183522 318008 216218 318064
rect 216274 318008 216279 318064
rect 183461 318006 216279 318008
rect 183461 318003 183527 318006
rect 216213 318003 216279 318006
rect 254577 318066 254643 318069
rect 270718 318066 270724 318068
rect 254577 318064 270724 318066
rect 254577 318008 254582 318064
rect 254638 318008 270724 318064
rect 254577 318006 270724 318008
rect 254577 318003 254643 318006
rect 270718 318004 270724 318006
rect 270788 318004 270794 318068
rect 81934 317460 81940 317524
rect 82004 317522 82010 317524
rect 82721 317522 82787 317525
rect 82004 317520 82787 317522
rect 82004 317464 82726 317520
rect 82782 317464 82787 317520
rect 82004 317462 82787 317464
rect 82004 317460 82010 317462
rect 82721 317459 82787 317462
rect 145557 317522 145623 317525
rect 207013 317522 207079 317525
rect 145557 317520 207079 317522
rect 145557 317464 145562 317520
rect 145618 317464 207018 317520
rect 207074 317464 207079 317520
rect 145557 317462 207079 317464
rect 145557 317459 145623 317462
rect 207013 317459 207079 317462
rect 182081 317386 182147 317389
rect 184197 317386 184263 317389
rect 182081 317384 184263 317386
rect 182081 317328 182086 317384
rect 182142 317328 184202 317384
rect 184258 317328 184263 317384
rect 182081 317326 184263 317328
rect 182081 317323 182147 317326
rect 184197 317323 184263 317326
rect 82721 316842 82787 316845
rect 90214 316842 90220 316844
rect 82721 316840 90220 316842
rect 82721 316784 82726 316840
rect 82782 316784 90220 316840
rect 82721 316782 90220 316784
rect 82721 316779 82787 316782
rect 90214 316780 90220 316782
rect 90284 316780 90290 316844
rect 86217 316706 86283 316709
rect 118734 316706 118740 316708
rect 86217 316704 118740 316706
rect 86217 316648 86222 316704
rect 86278 316648 118740 316704
rect 86217 316646 118740 316648
rect 86217 316643 86283 316646
rect 118734 316644 118740 316646
rect 118804 316706 118810 316708
rect 182081 316706 182147 316709
rect 118804 316704 182147 316706
rect 118804 316648 182086 316704
rect 182142 316648 182147 316704
rect 118804 316646 182147 316648
rect 118804 316644 118810 316646
rect 182081 316643 182147 316646
rect 191598 316644 191604 316708
rect 191668 316706 191674 316708
rect 232497 316706 232563 316709
rect 191668 316704 232563 316706
rect 191668 316648 232502 316704
rect 232558 316648 232563 316704
rect 191668 316646 232563 316648
rect 191668 316644 191674 316646
rect 232497 316643 232563 316646
rect 249057 316706 249123 316709
rect 263726 316706 263732 316708
rect 249057 316704 263732 316706
rect 249057 316648 249062 316704
rect 249118 316648 263732 316704
rect 249057 316646 263732 316648
rect 249057 316643 249123 316646
rect 263726 316644 263732 316646
rect 263796 316644 263802 316708
rect 259453 316570 259519 316573
rect 260046 316570 260052 316572
rect 259453 316568 260052 316570
rect 259453 316512 259458 316568
rect 259514 316512 260052 316568
rect 259453 316510 260052 316512
rect 259453 316507 259519 316510
rect 260046 316508 260052 316510
rect 260116 316508 260122 316572
rect 144177 316162 144243 316165
rect 200297 316162 200363 316165
rect 144177 316160 200363 316162
rect 144177 316104 144182 316160
rect 144238 316104 200302 316160
rect 200358 316104 200363 316160
rect 144177 316102 200363 316104
rect 144177 316099 144243 316102
rect 200297 316099 200363 316102
rect 170673 314938 170739 314941
rect 170949 314938 171015 314941
rect 244457 314938 244523 314941
rect 170673 314936 244523 314938
rect 170673 314880 170678 314936
rect 170734 314880 170954 314936
rect 171010 314880 244462 314936
rect 244518 314880 244523 314936
rect 170673 314878 244523 314880
rect 170673 314875 170739 314878
rect 170949 314875 171015 314878
rect 244457 314875 244523 314878
rect 33777 314802 33843 314805
rect 223113 314802 223179 314805
rect 33777 314800 223179 314802
rect 33777 314744 33782 314800
rect 33838 314744 223118 314800
rect 223174 314744 223179 314800
rect 33777 314742 223179 314744
rect 33777 314739 33843 314742
rect 223113 314739 223179 314742
rect 235257 314122 235323 314125
rect 254577 314122 254643 314125
rect 235257 314120 254643 314122
rect 235257 314064 235262 314120
rect 235318 314064 254582 314120
rect 254638 314064 254643 314120
rect 235257 314062 254643 314064
rect 235257 314059 235323 314062
rect 254577 314059 254643 314062
rect 205541 313986 205607 313989
rect 253933 313986 253999 313989
rect 205541 313984 253999 313986
rect 205541 313928 205546 313984
rect 205602 313928 253938 313984
rect 253994 313928 253999 313984
rect 205541 313926 253999 313928
rect 205541 313923 205607 313926
rect 253933 313923 253999 313926
rect 254761 313986 254827 313989
rect 259494 313986 259500 313988
rect 254761 313984 259500 313986
rect 254761 313928 254766 313984
rect 254822 313928 259500 313984
rect 254761 313926 259500 313928
rect 254761 313923 254827 313926
rect 259494 313924 259500 313926
rect 259564 313924 259570 313988
rect 262857 313986 262923 313989
rect 277158 313986 277164 313988
rect 262857 313984 277164 313986
rect 262857 313928 262862 313984
rect 262918 313928 277164 313984
rect 262857 313926 277164 313928
rect 262857 313923 262923 313926
rect 277158 313924 277164 313926
rect 277228 313924 277234 313988
rect 162117 313442 162183 313445
rect 162761 313442 162827 313445
rect 250713 313442 250779 313445
rect 162117 313440 250779 313442
rect 162117 313384 162122 313440
rect 162178 313384 162766 313440
rect 162822 313384 250718 313440
rect 250774 313384 250779 313440
rect 162117 313382 250779 313384
rect 162117 313379 162183 313382
rect 162761 313379 162827 313382
rect 250713 313379 250779 313382
rect 22737 313306 22803 313309
rect 220813 313306 220879 313309
rect 22737 313304 220879 313306
rect 22737 313248 22742 313304
rect 22798 313248 220818 313304
rect 220874 313248 220879 313304
rect 22737 313246 220879 313248
rect 22737 313243 22803 313246
rect 220813 313243 220879 313246
rect 82905 312490 82971 312493
rect 188613 312490 188679 312493
rect 82905 312488 188679 312490
rect 82905 312432 82910 312488
rect 82966 312432 188618 312488
rect 188674 312432 188679 312488
rect 82905 312430 188679 312432
rect 82905 312427 82971 312430
rect 188613 312427 188679 312430
rect 211797 312490 211863 312493
rect 261109 312490 261175 312493
rect 211797 312488 261175 312490
rect 211797 312432 211802 312488
rect 211858 312432 261114 312488
rect 261170 312432 261175 312488
rect 211797 312430 261175 312432
rect 211797 312427 211863 312430
rect 261109 312427 261175 312430
rect 188429 312082 188495 312085
rect 197445 312082 197511 312085
rect 188429 312080 197511 312082
rect 188429 312024 188434 312080
rect 188490 312024 197450 312080
rect 197506 312024 197511 312080
rect 188429 312022 197511 312024
rect 188429 312019 188495 312022
rect 197445 312019 197511 312022
rect 582557 312082 582623 312085
rect 583520 312082 584960 312172
rect 582557 312080 584960 312082
rect 582557 312024 582562 312080
rect 582618 312024 584960 312080
rect 582557 312022 584960 312024
rect 582557 312019 582623 312022
rect 30281 311946 30347 311949
rect 203425 311946 203491 311949
rect 30281 311944 203491 311946
rect 30281 311888 30286 311944
rect 30342 311888 203430 311944
rect 203486 311888 203491 311944
rect 583520 311932 584960 312022
rect 30281 311886 203491 311888
rect 30281 311883 30347 311886
rect 203425 311883 203491 311886
rect 216213 311266 216279 311269
rect 280245 311266 280311 311269
rect 281441 311266 281507 311269
rect 216213 311264 281507 311266
rect 216213 311208 216218 311264
rect 216274 311208 280250 311264
rect 280306 311208 281446 311264
rect 281502 311208 281507 311264
rect 216213 311206 281507 311208
rect 216213 311203 216279 311206
rect 280245 311203 280311 311206
rect 281441 311203 281507 311206
rect 61653 311130 61719 311133
rect 61837 311130 61903 311133
rect 280337 311130 280403 311133
rect 280797 311130 280863 311133
rect 61653 311128 280863 311130
rect 61653 311072 61658 311128
rect 61714 311072 61842 311128
rect 61898 311072 280342 311128
rect 280398 311072 280802 311128
rect 280858 311072 280863 311128
rect 61653 311070 280863 311072
rect 61653 311067 61719 311070
rect 61837 311067 61903 311070
rect 280337 311067 280403 311070
rect 280797 311067 280863 311070
rect 122741 310722 122807 310725
rect 219985 310722 220051 310725
rect 122741 310720 220051 310722
rect 122741 310664 122746 310720
rect 122802 310664 219990 310720
rect 220046 310664 220051 310720
rect 122741 310662 220051 310664
rect 122741 310659 122807 310662
rect 219985 310659 220051 310662
rect 41137 310586 41203 310589
rect 205633 310586 205699 310589
rect 41137 310584 205699 310586
rect 41137 310528 41142 310584
rect 41198 310528 205638 310584
rect 205694 310528 205699 310584
rect 41137 310526 205699 310528
rect 41137 310523 41203 310526
rect 205633 310523 205699 310526
rect 185669 309498 185735 309501
rect 256734 309498 256740 309500
rect 185669 309496 256740 309498
rect 185669 309440 185674 309496
rect 185730 309440 256740 309496
rect 185669 309438 256740 309440
rect 185669 309435 185735 309438
rect 256734 309436 256740 309438
rect 256804 309436 256810 309500
rect 177297 309362 177363 309365
rect 267733 309362 267799 309365
rect 177297 309360 267799 309362
rect 177297 309304 177302 309360
rect 177358 309304 267738 309360
rect 267794 309304 267799 309360
rect 177297 309302 267799 309304
rect 177297 309299 177363 309302
rect 267733 309299 267799 309302
rect 1301 309226 1367 309229
rect 200205 309226 200271 309229
rect 1301 309224 200271 309226
rect 1301 309168 1306 309224
rect 1362 309168 200210 309224
rect 200266 309168 200271 309224
rect 1301 309166 200271 309168
rect 1301 309163 1367 309166
rect 200205 309163 200271 309166
rect 269113 309090 269179 309093
rect 269389 309090 269455 309093
rect 269113 309088 269455 309090
rect 269113 309032 269118 309088
rect 269174 309032 269394 309088
rect 269450 309032 269455 309088
rect 269113 309030 269455 309032
rect 269113 309027 269179 309030
rect 269389 309027 269455 309030
rect 246297 308546 246363 308549
rect 254209 308546 254275 308549
rect 246297 308544 254275 308546
rect 246297 308488 246302 308544
rect 246358 308488 254214 308544
rect 254270 308488 254275 308544
rect 246297 308486 254275 308488
rect 246297 308483 246363 308486
rect 254209 308483 254275 308486
rect 218053 308410 218119 308413
rect 244549 308410 244615 308413
rect 218053 308408 244615 308410
rect 218053 308352 218058 308408
rect 218114 308352 244554 308408
rect 244610 308352 244615 308408
rect 218053 308350 244615 308352
rect 218053 308347 218119 308350
rect 244549 308347 244615 308350
rect 251909 308410 251975 308413
rect 267917 308410 267983 308413
rect 251909 308408 267983 308410
rect 251909 308352 251914 308408
rect 251970 308352 267922 308408
rect 267978 308352 267983 308408
rect 251909 308350 267983 308352
rect 251909 308347 251975 308350
rect 267917 308347 267983 308350
rect 184197 308138 184263 308141
rect 212717 308138 212783 308141
rect 184197 308136 212783 308138
rect 184197 308080 184202 308136
rect 184258 308080 212722 308136
rect 212778 308080 212783 308136
rect 184197 308078 212783 308080
rect 184197 308075 184263 308078
rect 212717 308075 212783 308078
rect 88977 308002 89043 308005
rect 88977 308000 258090 308002
rect 88977 307944 88982 308000
rect 89038 307944 258090 308000
rect 88977 307942 258090 307944
rect 88977 307939 89043 307942
rect 17861 307866 17927 307869
rect 202045 307866 202111 307869
rect 17861 307864 202111 307866
rect 17861 307808 17866 307864
rect 17922 307808 202050 307864
rect 202106 307808 202111 307864
rect 17861 307806 202111 307808
rect 258030 307866 258090 307942
rect 269389 307866 269455 307869
rect 258030 307864 269455 307866
rect 258030 307808 269394 307864
rect 269450 307808 269455 307864
rect 258030 307806 269455 307808
rect 17861 307803 17927 307806
rect 202045 307803 202111 307806
rect 269389 307803 269455 307806
rect 206134 307668 206140 307732
rect 206204 307730 206210 307732
rect 207105 307730 207171 307733
rect 206204 307728 207171 307730
rect 206204 307672 207110 307728
rect 207166 307672 207171 307728
rect 206204 307670 207171 307672
rect 206204 307668 206210 307670
rect 207105 307667 207171 307670
rect 222193 307730 222259 307733
rect 224166 307730 224172 307732
rect 222193 307728 224172 307730
rect 222193 307672 222198 307728
rect 222254 307672 224172 307728
rect 222193 307670 224172 307672
rect 222193 307667 222259 307670
rect 224166 307668 224172 307670
rect 224236 307668 224242 307732
rect 249333 307730 249399 307733
rect 249701 307730 249767 307733
rect 249333 307728 249767 307730
rect 249333 307672 249338 307728
rect 249394 307672 249706 307728
rect 249762 307672 249767 307728
rect 249333 307670 249767 307672
rect 249333 307667 249399 307670
rect 249701 307667 249767 307670
rect 238109 307186 238175 307189
rect 251265 307186 251331 307189
rect 238109 307184 251331 307186
rect 238109 307128 238114 307184
rect 238170 307128 251270 307184
rect 251326 307128 251331 307184
rect 238109 307126 251331 307128
rect 238109 307123 238175 307126
rect 251265 307123 251331 307126
rect 207105 307050 207171 307053
rect 255262 307050 255268 307052
rect 207105 307048 255268 307050
rect 207105 306992 207110 307048
rect 207166 306992 255268 307048
rect 207105 306990 255268 306992
rect 207105 306987 207171 306990
rect 255262 306988 255268 306990
rect 255332 306988 255338 307052
rect 32397 306778 32463 306781
rect 221549 306778 221615 306781
rect 32397 306776 221615 306778
rect 32397 306720 32402 306776
rect 32458 306720 221554 306776
rect 221610 306720 221615 306776
rect 32397 306718 221615 306720
rect 32397 306715 32463 306718
rect 221549 306715 221615 306718
rect 192569 306642 192635 306645
rect 210233 306642 210299 306645
rect 192569 306640 210299 306642
rect 192569 306584 192574 306640
rect 192630 306584 210238 306640
rect 210294 306584 210299 306640
rect 192569 306582 210299 306584
rect 192569 306579 192635 306582
rect 210233 306579 210299 306582
rect 189993 306506 190059 306509
rect 199469 306506 199535 306509
rect 189993 306504 199535 306506
rect 189993 306448 189998 306504
rect 190054 306448 199474 306504
rect 199530 306448 199535 306504
rect 189993 306446 199535 306448
rect 189993 306443 190059 306446
rect 199469 306443 199535 306446
rect 230238 306444 230244 306508
rect 230308 306506 230314 306508
rect 245837 306506 245903 306509
rect 230308 306504 245903 306506
rect 230308 306448 245842 306504
rect 245898 306448 245903 306504
rect 230308 306446 245903 306448
rect 230308 306444 230314 306446
rect 245837 306443 245903 306446
rect 249333 306506 249399 306509
rect 277669 306506 277735 306509
rect 249333 306504 277735 306506
rect 249333 306448 249338 306504
rect 249394 306448 277674 306504
rect 277730 306448 277735 306504
rect 249333 306446 277735 306448
rect 249333 306443 249399 306446
rect 277669 306443 277735 306446
rect -960 306234 480 306324
rect 3233 306234 3299 306237
rect -960 306232 3299 306234
rect -960 306176 3238 306232
rect 3294 306176 3299 306232
rect -960 306174 3299 306176
rect -960 306084 480 306174
rect 3233 306171 3299 306174
rect 260097 305826 260163 305829
rect 273294 305826 273300 305828
rect 260097 305824 273300 305826
rect 260097 305768 260102 305824
rect 260158 305768 273300 305824
rect 260097 305766 273300 305768
rect 260097 305763 260163 305766
rect 273294 305764 273300 305766
rect 273364 305764 273370 305828
rect 96521 305690 96587 305693
rect 108982 305690 108988 305692
rect 96521 305688 108988 305690
rect 96521 305632 96526 305688
rect 96582 305632 108988 305688
rect 96521 305630 108988 305632
rect 96521 305627 96587 305630
rect 108982 305628 108988 305630
rect 109052 305628 109058 305692
rect 233877 305690 233943 305693
rect 265065 305690 265131 305693
rect 233877 305688 265131 305690
rect 233877 305632 233882 305688
rect 233938 305632 265070 305688
rect 265126 305632 265131 305688
rect 233877 305630 265131 305632
rect 233877 305627 233943 305630
rect 265065 305627 265131 305630
rect 184054 305220 184060 305284
rect 184124 305282 184130 305284
rect 209589 305282 209655 305285
rect 184124 305280 209655 305282
rect 184124 305224 209594 305280
rect 209650 305224 209655 305280
rect 184124 305222 209655 305224
rect 184124 305220 184130 305222
rect 209589 305219 209655 305222
rect 220486 305220 220492 305284
rect 220556 305282 220562 305284
rect 220556 305222 229110 305282
rect 220556 305220 220562 305222
rect 91134 305146 91140 305148
rect 84150 305086 91140 305146
rect 75177 305010 75243 305013
rect 81934 305010 81940 305012
rect 75177 305008 81940 305010
rect 75177 304952 75182 305008
rect 75238 304952 81940 305008
rect 75177 304950 81940 304952
rect 75177 304947 75243 304950
rect 81934 304948 81940 304950
rect 82004 304948 82010 305012
rect 83457 305010 83523 305013
rect 84150 305010 84210 305086
rect 91134 305084 91140 305086
rect 91204 305084 91210 305148
rect 187693 305146 187759 305149
rect 214005 305146 214071 305149
rect 187693 305144 214071 305146
rect 187693 305088 187698 305144
rect 187754 305088 214010 305144
rect 214066 305088 214071 305144
rect 187693 305086 214071 305088
rect 187693 305083 187759 305086
rect 214005 305083 214071 305086
rect 226190 305084 226196 305148
rect 226260 305146 226266 305148
rect 227713 305146 227779 305149
rect 226260 305144 227779 305146
rect 226260 305088 227718 305144
rect 227774 305088 227779 305144
rect 226260 305086 227779 305088
rect 229050 305146 229110 305222
rect 241462 305146 241468 305148
rect 229050 305086 241468 305146
rect 226260 305084 226266 305086
rect 227713 305083 227779 305086
rect 241462 305084 241468 305086
rect 241532 305084 241538 305148
rect 83457 305008 84210 305010
rect 83457 304952 83462 305008
rect 83518 304952 84210 305008
rect 83457 304950 84210 304952
rect 83457 304947 83523 304950
rect 90950 304948 90956 305012
rect 91020 305010 91026 305012
rect 95233 305010 95299 305013
rect 91020 305008 95299 305010
rect 91020 304952 95238 305008
rect 95294 304952 95299 305008
rect 91020 304950 95299 304952
rect 91020 304948 91026 304950
rect 95233 304947 95299 304950
rect 176009 305010 176075 305013
rect 176561 305010 176627 305013
rect 269113 305010 269179 305013
rect 176009 305008 269179 305010
rect 176009 304952 176014 305008
rect 176070 304952 176566 305008
rect 176622 304952 269118 305008
rect 269174 304952 269179 305008
rect 176009 304950 269179 304952
rect 176009 304947 176075 304950
rect 176561 304947 176627 304950
rect 269113 304947 269179 304950
rect 101673 304194 101739 304197
rect 122925 304194 122991 304197
rect 101673 304192 122991 304194
rect 101673 304136 101678 304192
rect 101734 304136 122930 304192
rect 122986 304136 122991 304192
rect 101673 304134 122991 304136
rect 101673 304131 101739 304134
rect 122925 304131 122991 304134
rect 241646 304132 241652 304196
rect 241716 304194 241722 304196
rect 242801 304194 242867 304197
rect 241716 304192 242867 304194
rect 241716 304136 242806 304192
rect 242862 304136 242867 304192
rect 241716 304134 242867 304136
rect 241716 304132 241722 304134
rect 242801 304131 242867 304134
rect 152457 303922 152523 303925
rect 213361 303922 213427 303925
rect 152457 303920 213427 303922
rect 152457 303864 152462 303920
rect 152518 303864 213366 303920
rect 213422 303864 213427 303920
rect 152457 303862 213427 303864
rect 152457 303859 152523 303862
rect 213361 303859 213427 303862
rect 217542 303860 217548 303924
rect 217612 303922 217618 303924
rect 251909 303922 251975 303925
rect 217612 303920 251975 303922
rect 217612 303864 251914 303920
rect 251970 303864 251975 303920
rect 217612 303862 251975 303864
rect 217612 303860 217618 303862
rect 251909 303859 251975 303862
rect 186814 303724 186820 303788
rect 186884 303786 186890 303788
rect 195697 303786 195763 303789
rect 186884 303784 195763 303786
rect 186884 303728 195702 303784
rect 195758 303728 195763 303784
rect 186884 303726 195763 303728
rect 186884 303724 186890 303726
rect 195697 303723 195763 303726
rect 213678 303724 213684 303788
rect 213748 303786 213754 303788
rect 229185 303786 229251 303789
rect 274582 303786 274588 303788
rect 213748 303784 229251 303786
rect 213748 303728 229190 303784
rect 229246 303728 229251 303784
rect 213748 303726 229251 303728
rect 213748 303724 213754 303726
rect 229185 303723 229251 303726
rect 248370 303726 274588 303786
rect 211654 303588 211660 303652
rect 211724 303650 211730 303652
rect 218053 303650 218119 303653
rect 211724 303648 218119 303650
rect 211724 303592 218058 303648
rect 218114 303592 218119 303648
rect 211724 303590 218119 303592
rect 211724 303588 211730 303590
rect 218053 303587 218119 303590
rect 240869 303650 240935 303653
rect 245561 303650 245627 303653
rect 248370 303650 248430 303726
rect 274582 303724 274588 303726
rect 274652 303724 274658 303788
rect 240869 303648 248430 303650
rect 240869 303592 240874 303648
rect 240930 303592 245566 303648
rect 245622 303592 248430 303648
rect 240869 303590 248430 303592
rect 251265 303650 251331 303653
rect 282913 303650 282979 303653
rect 251265 303648 282979 303650
rect 251265 303592 251270 303648
rect 251326 303592 282918 303648
rect 282974 303592 282979 303648
rect 251265 303590 282979 303592
rect 240869 303587 240935 303590
rect 245561 303587 245627 303590
rect 251265 303587 251331 303590
rect 282913 303587 282979 303590
rect 198089 303514 198155 303517
rect 200614 303514 200620 303516
rect 198089 303512 200620 303514
rect 198089 303456 198094 303512
rect 198150 303456 200620 303512
rect 198089 303454 200620 303456
rect 198089 303451 198155 303454
rect 200614 303452 200620 303454
rect 200684 303514 200690 303516
rect 201401 303514 201467 303517
rect 200684 303512 201467 303514
rect 200684 303456 201406 303512
rect 201462 303456 201467 303512
rect 200684 303454 201467 303456
rect 200684 303452 200690 303454
rect 201401 303451 201467 303454
rect 89529 302834 89595 302837
rect 99966 302834 99972 302836
rect 89529 302832 99972 302834
rect 89529 302776 89534 302832
rect 89590 302776 99972 302832
rect 89529 302774 99972 302776
rect 89529 302771 89595 302774
rect 99966 302772 99972 302774
rect 100036 302772 100042 302836
rect 250713 302834 250779 302837
rect 259729 302834 259795 302837
rect 250713 302832 259795 302834
rect 250713 302776 250718 302832
rect 250774 302776 259734 302832
rect 259790 302776 259795 302832
rect 250713 302774 259795 302776
rect 250713 302771 250779 302774
rect 259729 302771 259795 302774
rect 26141 302562 26207 302565
rect 200113 302562 200179 302565
rect 26141 302560 200179 302562
rect 26141 302504 26146 302560
rect 26202 302504 200118 302560
rect 200174 302504 200179 302560
rect 26141 302502 200179 302504
rect 26141 302499 26207 302502
rect 200113 302499 200179 302502
rect 131757 302426 131823 302429
rect 207657 302426 207723 302429
rect 131757 302424 207723 302426
rect 131757 302368 131762 302424
rect 131818 302368 207662 302424
rect 207718 302368 207723 302424
rect 131757 302366 207723 302368
rect 131757 302363 131823 302366
rect 207657 302363 207723 302366
rect 248781 302426 248847 302429
rect 249609 302426 249675 302429
rect 278773 302426 278839 302429
rect 248781 302424 278839 302426
rect 248781 302368 248786 302424
rect 248842 302368 249614 302424
rect 249670 302368 278778 302424
rect 278834 302368 278839 302424
rect 248781 302366 278839 302368
rect 248781 302363 248847 302366
rect 249609 302363 249675 302366
rect 278773 302363 278839 302366
rect 192753 302292 192819 302293
rect 192702 302290 192708 302292
rect 192662 302230 192708 302290
rect 192772 302288 192819 302292
rect 192814 302232 192819 302288
rect 192702 302228 192708 302230
rect 192772 302228 192819 302232
rect 192753 302227 192819 302228
rect 192937 302290 193003 302293
rect 194542 302290 194548 302292
rect 192937 302288 194548 302290
rect 192937 302232 192942 302288
rect 192998 302232 194548 302288
rect 192937 302230 194548 302232
rect 192937 302227 193003 302230
rect 194542 302228 194548 302230
rect 194612 302228 194618 302292
rect 214414 302228 214420 302292
rect 214484 302290 214490 302292
rect 229829 302290 229895 302293
rect 214484 302288 229895 302290
rect 214484 302232 229834 302288
rect 229890 302232 229895 302288
rect 214484 302230 229895 302232
rect 214484 302228 214490 302230
rect 229829 302227 229895 302230
rect 236085 302290 236151 302293
rect 240726 302290 240732 302292
rect 236085 302288 240732 302290
rect 236085 302232 236090 302288
rect 236146 302232 240732 302288
rect 236085 302230 240732 302232
rect 236085 302227 236151 302230
rect 240726 302228 240732 302230
rect 240796 302228 240802 302292
rect 241145 302290 241211 302293
rect 582465 302290 582531 302293
rect 241145 302288 582531 302290
rect 241145 302232 241150 302288
rect 241206 302232 582470 302288
rect 582526 302232 582531 302288
rect 241145 302230 582531 302232
rect 241145 302227 241211 302230
rect 582465 302227 582531 302230
rect 220854 301820 220860 301884
rect 220924 301882 220930 301884
rect 225045 301882 225111 301885
rect 220924 301880 225111 301882
rect 220924 301824 225050 301880
rect 225106 301824 225111 301880
rect 220924 301822 225111 301824
rect 220924 301820 220930 301822
rect 225045 301819 225111 301822
rect 240225 301746 240291 301749
rect 241053 301746 241119 301749
rect 245745 301746 245811 301749
rect 219390 301744 241119 301746
rect 219390 301688 240230 301744
rect 240286 301688 241058 301744
rect 241114 301688 241119 301744
rect 219390 301686 241119 301688
rect 191097 301610 191163 301613
rect 191598 301610 191604 301612
rect 191097 301608 191604 301610
rect 191097 301552 191102 301608
rect 191158 301552 191604 301608
rect 191097 301550 191604 301552
rect 191097 301547 191163 301550
rect 191598 301548 191604 301550
rect 191668 301548 191674 301612
rect 193254 301548 193260 301612
rect 193324 301610 193330 301612
rect 194133 301610 194199 301613
rect 193324 301608 194199 301610
rect 193324 301552 194138 301608
rect 194194 301552 194199 301608
rect 193324 301550 194199 301552
rect 193324 301548 193330 301550
rect 194133 301547 194199 301550
rect 91134 301412 91140 301476
rect 91204 301474 91210 301476
rect 122833 301474 122899 301477
rect 91204 301472 122899 301474
rect 91204 301416 122838 301472
rect 122894 301416 122899 301472
rect 91204 301414 122899 301416
rect 91204 301412 91210 301414
rect 122833 301411 122899 301414
rect 148409 301474 148475 301477
rect 203057 301474 203123 301477
rect 204345 301476 204411 301477
rect 204294 301474 204300 301476
rect 148409 301472 203123 301474
rect 148409 301416 148414 301472
rect 148470 301416 203062 301472
rect 203118 301416 203123 301472
rect 148409 301414 203123 301416
rect 204254 301414 204300 301474
rect 204364 301472 204411 301476
rect 204406 301416 204411 301472
rect 148409 301411 148475 301414
rect 203057 301411 203123 301414
rect 204294 301412 204300 301414
rect 204364 301412 204411 301416
rect 204345 301411 204411 301412
rect 207013 301476 207079 301477
rect 210601 301476 210667 301477
rect 207013 301472 207060 301476
rect 207124 301474 207130 301476
rect 210550 301474 210556 301476
rect 207013 301416 207018 301472
rect 207013 301412 207060 301416
rect 207124 301414 207170 301474
rect 210510 301414 210556 301474
rect 210620 301472 210667 301476
rect 210662 301416 210667 301472
rect 207124 301412 207130 301414
rect 210550 301412 210556 301414
rect 210620 301412 210667 301416
rect 215886 301412 215892 301476
rect 215956 301474 215962 301476
rect 216765 301474 216831 301477
rect 215956 301472 216831 301474
rect 215956 301416 216770 301472
rect 216826 301416 216831 301472
rect 215956 301414 216831 301416
rect 215956 301412 215962 301414
rect 207013 301411 207079 301412
rect 210601 301411 210667 301412
rect 216765 301411 216831 301414
rect 219198 301412 219204 301476
rect 219268 301474 219274 301476
rect 219390 301474 219450 301686
rect 240225 301683 240291 301686
rect 241053 301683 241119 301686
rect 245702 301744 245811 301746
rect 245702 301688 245750 301744
rect 245806 301688 245811 301744
rect 245702 301683 245811 301688
rect 222326 301548 222332 301612
rect 222396 301610 222402 301612
rect 222561 301610 222627 301613
rect 222396 301608 222627 301610
rect 222396 301552 222566 301608
rect 222622 301552 222627 301608
rect 222396 301550 222627 301552
rect 222396 301548 222402 301550
rect 222561 301547 222627 301550
rect 226558 301548 226564 301612
rect 226628 301610 226634 301612
rect 226977 301610 227043 301613
rect 226628 301608 227043 301610
rect 226628 301552 226982 301608
rect 227038 301552 227043 301608
rect 226628 301550 227043 301552
rect 226628 301548 226634 301550
rect 226977 301547 227043 301550
rect 230422 301548 230428 301612
rect 230492 301610 230498 301612
rect 231301 301610 231367 301613
rect 230492 301608 231367 301610
rect 230492 301552 231306 301608
rect 231362 301552 231367 301608
rect 230492 301550 231367 301552
rect 230492 301548 230498 301550
rect 231301 301547 231367 301550
rect 234654 301548 234660 301612
rect 234724 301610 234730 301612
rect 235257 301610 235323 301613
rect 234724 301608 235323 301610
rect 234724 301552 235262 301608
rect 235318 301552 235323 301608
rect 234724 301550 235323 301552
rect 234724 301548 234730 301550
rect 235257 301547 235323 301550
rect 237598 301548 237604 301612
rect 237668 301610 237674 301612
rect 237741 301610 237807 301613
rect 237668 301608 237807 301610
rect 237668 301552 237746 301608
rect 237802 301552 237807 301608
rect 237668 301550 237807 301552
rect 237668 301548 237674 301550
rect 237741 301547 237807 301550
rect 219268 301414 219450 301474
rect 222561 301474 222627 301477
rect 222694 301474 222700 301476
rect 222561 301472 222700 301474
rect 222561 301416 222566 301472
rect 222622 301416 222700 301472
rect 222561 301414 222700 301416
rect 219268 301412 219274 301414
rect 222561 301411 222627 301414
rect 222694 301412 222700 301414
rect 222764 301412 222770 301476
rect 223614 301412 223620 301476
rect 223684 301474 223690 301476
rect 223849 301474 223915 301477
rect 223684 301472 223915 301474
rect 223684 301416 223854 301472
rect 223910 301416 223915 301472
rect 223684 301414 223915 301416
rect 223684 301412 223690 301414
rect 223849 301411 223915 301414
rect 224902 301412 224908 301476
rect 224972 301474 224978 301476
rect 225781 301474 225847 301477
rect 224972 301472 225847 301474
rect 224972 301416 225786 301472
rect 225842 301416 225847 301472
rect 224972 301414 225847 301416
rect 224972 301412 224978 301414
rect 225781 301411 225847 301414
rect 226701 301476 226767 301477
rect 226701 301472 226748 301476
rect 226812 301474 226818 301476
rect 226701 301416 226706 301472
rect 226701 301412 226748 301416
rect 226812 301414 226858 301474
rect 226812 301412 226818 301414
rect 227662 301412 227668 301476
rect 227732 301474 227738 301476
rect 228265 301474 228331 301477
rect 227732 301472 228331 301474
rect 227732 301416 228270 301472
rect 228326 301416 228331 301472
rect 227732 301414 228331 301416
rect 227732 301412 227738 301414
rect 226701 301411 226767 301412
rect 228265 301411 228331 301414
rect 229686 301412 229692 301476
rect 229756 301474 229762 301476
rect 230105 301474 230171 301477
rect 229756 301472 230171 301474
rect 229756 301416 230110 301472
rect 230166 301416 230171 301472
rect 229756 301414 230171 301416
rect 229756 301412 229762 301414
rect 230105 301411 230171 301414
rect 230565 301476 230631 301477
rect 232129 301476 232195 301477
rect 230565 301472 230612 301476
rect 230676 301474 230682 301476
rect 232078 301474 232084 301476
rect 230565 301416 230570 301472
rect 230565 301412 230612 301416
rect 230676 301414 230722 301474
rect 232038 301414 232084 301474
rect 232148 301472 232195 301476
rect 232190 301416 232195 301472
rect 230676 301412 230682 301414
rect 232078 301412 232084 301414
rect 232148 301412 232195 301416
rect 232262 301412 232268 301476
rect 232332 301474 232338 301476
rect 232681 301474 232747 301477
rect 232332 301472 232747 301474
rect 232332 301416 232686 301472
rect 232742 301416 232747 301472
rect 232332 301414 232747 301416
rect 232332 301412 232338 301414
rect 230565 301411 230631 301412
rect 232129 301411 232195 301412
rect 232681 301411 232747 301414
rect 233182 301412 233188 301476
rect 233252 301474 233258 301476
rect 233325 301474 233391 301477
rect 233252 301472 233391 301474
rect 233252 301416 233330 301472
rect 233386 301416 233391 301472
rect 233252 301414 233391 301416
rect 233252 301412 233258 301414
rect 233325 301411 233391 301414
rect 233550 301412 233556 301476
rect 233620 301474 233626 301476
rect 233969 301474 234035 301477
rect 233620 301472 234035 301474
rect 233620 301416 233974 301472
rect 234030 301416 234035 301472
rect 233620 301414 234035 301416
rect 233620 301412 233626 301414
rect 233969 301411 234035 301414
rect 234797 301476 234863 301477
rect 236637 301476 236703 301477
rect 234797 301472 234844 301476
rect 234908 301474 234914 301476
rect 234797 301416 234802 301472
rect 234797 301412 234844 301416
rect 234908 301414 234954 301474
rect 236637 301472 236684 301476
rect 236748 301474 236754 301476
rect 237649 301474 237715 301477
rect 237782 301474 237788 301476
rect 236637 301416 236642 301472
rect 234908 301412 234914 301414
rect 236637 301412 236684 301416
rect 236748 301414 236794 301474
rect 237649 301472 237788 301474
rect 237649 301416 237654 301472
rect 237710 301416 237788 301472
rect 237649 301414 237788 301416
rect 236748 301412 236754 301414
rect 234797 301411 234863 301412
rect 236637 301411 236703 301412
rect 237649 301411 237715 301414
rect 237782 301412 237788 301414
rect 237852 301412 237858 301476
rect 238518 301412 238524 301476
rect 238588 301474 238594 301476
rect 239673 301474 239739 301477
rect 238588 301472 239739 301474
rect 238588 301416 239678 301472
rect 239734 301416 239739 301472
rect 238588 301414 239739 301416
rect 238588 301412 238594 301414
rect 239673 301411 239739 301414
rect 242934 301412 242940 301476
rect 243004 301474 243010 301476
rect 243445 301474 243511 301477
rect 243004 301472 243511 301474
rect 243004 301416 243450 301472
rect 243506 301416 243511 301472
rect 243004 301414 243511 301416
rect 243004 301412 243010 301414
rect 243445 301411 243511 301414
rect 245510 301412 245516 301476
rect 245580 301474 245586 301476
rect 245702 301474 245762 301683
rect 245878 301548 245884 301612
rect 245948 301610 245954 301612
rect 246481 301610 246547 301613
rect 245948 301608 246547 301610
rect 245948 301552 246486 301608
rect 246542 301552 246547 301608
rect 245948 301550 246547 301552
rect 245948 301548 245954 301550
rect 246481 301547 246547 301550
rect 246573 301474 246639 301477
rect 245580 301472 246639 301474
rect 245580 301416 246578 301472
rect 246634 301416 246639 301472
rect 245580 301414 246639 301416
rect 245580 301412 245586 301414
rect 246573 301411 246639 301414
rect 247718 301412 247724 301476
rect 247788 301474 247794 301476
rect 247861 301474 247927 301477
rect 247788 301472 247927 301474
rect 247788 301416 247866 301472
rect 247922 301416 247927 301472
rect 247788 301414 247927 301416
rect 247788 301412 247794 301414
rect 247861 301411 247927 301414
rect 250253 301474 250319 301477
rect 258390 301474 258396 301476
rect 250253 301472 258396 301474
rect 250253 301416 250258 301472
rect 250314 301416 258396 301472
rect 250253 301414 258396 301416
rect 250253 301411 250319 301414
rect 258390 301412 258396 301414
rect 258460 301412 258466 301476
rect 253657 301338 253723 301341
rect 253430 301336 253723 301338
rect 253430 301280 253662 301336
rect 253718 301280 253723 301336
rect 253430 301278 253723 301280
rect 253430 301172 253490 301278
rect 253657 301275 253723 301278
rect 191097 301066 191163 301069
rect 191097 301064 193690 301066
rect 191097 301008 191102 301064
rect 191158 301008 193690 301064
rect 191097 301006 193690 301008
rect 191097 301003 191163 301006
rect 133137 300930 133203 300933
rect 191741 300930 191807 300933
rect 133137 300928 191807 300930
rect 133137 300872 133142 300928
rect 133198 300872 191746 300928
rect 191802 300872 191807 300928
rect 193630 300900 193690 301006
rect 133137 300870 191807 300872
rect 133137 300867 133203 300870
rect 191741 300867 191807 300870
rect 84694 300732 84700 300796
rect 84764 300794 84770 300796
rect 87045 300794 87111 300797
rect 84764 300792 87111 300794
rect 84764 300736 87050 300792
rect 87106 300736 87111 300792
rect 84764 300734 87111 300736
rect 84764 300732 84770 300734
rect 87045 300731 87111 300734
rect 87454 300732 87460 300796
rect 87524 300794 87530 300796
rect 89713 300794 89779 300797
rect 256601 300794 256667 300797
rect 87524 300792 89779 300794
rect 87524 300736 89718 300792
rect 89774 300736 89779 300792
rect 252908 300792 256667 300794
rect 252908 300764 256606 300792
rect 87524 300734 89779 300736
rect 87524 300732 87530 300734
rect 89713 300731 89779 300734
rect 252878 300736 256606 300764
rect 256662 300736 256667 300792
rect 252878 300734 256667 300736
rect 252878 300660 252938 300734
rect 256601 300731 256667 300734
rect 252870 300596 252876 300660
rect 252940 300596 252946 300660
rect 256509 300386 256575 300389
rect 253460 300384 256575 300386
rect 253460 300328 256514 300384
rect 256570 300328 256575 300384
rect 253460 300326 256575 300328
rect 256509 300323 256575 300326
rect 252829 300250 252895 300253
rect 252829 300248 252938 300250
rect 252829 300192 252834 300248
rect 252890 300192 252938 300248
rect 252829 300187 252938 300192
rect 181529 300114 181595 300117
rect 193254 300114 193260 300116
rect 181529 300112 193260 300114
rect 181529 300056 181534 300112
rect 181590 300056 193260 300112
rect 181529 300054 193260 300056
rect 181529 300051 181595 300054
rect 193254 300052 193260 300054
rect 193324 300052 193330 300116
rect 191741 299978 191807 299981
rect 191741 299976 193660 299978
rect 191741 299920 191746 299976
rect 191802 299920 193660 299976
rect 252878 299948 252938 300187
rect 191741 299918 193660 299920
rect 191741 299915 191807 299918
rect 191966 299508 191972 299572
rect 192036 299570 192042 299572
rect 192201 299570 192267 299573
rect 273253 299570 273319 299573
rect 192036 299568 192267 299570
rect 192036 299512 192206 299568
rect 192262 299512 192267 299568
rect 192036 299510 192267 299512
rect 253460 299568 273319 299570
rect 253460 299512 273258 299568
rect 273314 299512 273319 299568
rect 253460 299510 273319 299512
rect 192036 299508 192042 299510
rect 192201 299507 192267 299510
rect 273253 299507 273319 299510
rect 272517 299436 272583 299437
rect 272517 299432 272564 299436
rect 272628 299434 272634 299436
rect 272517 299376 272522 299432
rect 272517 299372 272564 299376
rect 272628 299374 272674 299434
rect 272628 299372 272634 299374
rect 272517 299371 272583 299372
rect 253460 299102 253950 299162
rect 190637 299026 190703 299029
rect 253105 299026 253171 299029
rect 190637 299024 193660 299026
rect 190637 298968 190642 299024
rect 190698 298968 193660 299024
rect 190637 298966 193660 298968
rect 253062 299024 253171 299026
rect 253062 298968 253110 299024
rect 253166 298968 253171 299024
rect 190637 298963 190703 298966
rect 253062 298963 253171 298968
rect 173014 298828 173020 298892
rect 173084 298890 173090 298892
rect 187693 298890 187759 298893
rect 173084 298888 187759 298890
rect 173084 298832 187698 298888
rect 187754 298832 187759 298888
rect 173084 298830 187759 298832
rect 173084 298828 173090 298830
rect 187693 298827 187759 298830
rect 91502 298692 91508 298756
rect 91572 298754 91578 298756
rect 96613 298754 96679 298757
rect 91572 298752 96679 298754
rect 91572 298696 96618 298752
rect 96674 298696 96679 298752
rect 91572 298694 96679 298696
rect 91572 298692 91578 298694
rect 96613 298691 96679 298694
rect 126237 298754 126303 298757
rect 193581 298754 193647 298757
rect 126237 298752 193647 298754
rect 126237 298696 126242 298752
rect 126298 298696 193586 298752
rect 193642 298696 193647 298752
rect 253062 298724 253122 298963
rect 253890 298754 253950 299102
rect 256969 298754 257035 298757
rect 265750 298754 265756 298756
rect 253890 298752 265756 298754
rect 126237 298694 193647 298696
rect 253890 298696 256974 298752
rect 257030 298696 265756 298752
rect 253890 298694 265756 298696
rect 126237 298691 126303 298694
rect 193581 298691 193647 298694
rect 256969 298691 257035 298694
rect 265750 298692 265756 298694
rect 265820 298692 265826 298756
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect 256601 298346 256667 298349
rect 253460 298344 256667 298346
rect 253460 298288 256606 298344
rect 256662 298288 256667 298344
rect 253460 298286 256667 298288
rect 256601 298283 256667 298286
rect 39941 298210 40007 298213
rect 113817 298210 113883 298213
rect 39941 298208 113883 298210
rect 39941 298152 39946 298208
rect 40002 298152 113822 298208
rect 113878 298152 113883 298208
rect 39941 298150 113883 298152
rect 39941 298147 40007 298150
rect 113817 298147 113883 298150
rect 188286 298148 188292 298212
rect 188356 298210 188362 298212
rect 192569 298210 192635 298213
rect 188356 298208 192635 298210
rect 188356 298152 192574 298208
rect 192630 298152 192635 298208
rect 188356 298150 192635 298152
rect 188356 298148 188362 298150
rect 192569 298147 192635 298150
rect 191465 298076 191531 298077
rect 191414 298074 191420 298076
rect 191338 298014 191420 298074
rect 191484 298074 191531 298076
rect 266353 298074 266419 298077
rect 267774 298074 267780 298076
rect 191484 298072 193660 298074
rect 191526 298016 193660 298072
rect 191414 298012 191420 298014
rect 191484 298014 193660 298016
rect 266353 298072 267780 298074
rect 266353 298016 266358 298072
rect 266414 298016 267780 298072
rect 266353 298014 267780 298016
rect 191484 298012 191531 298014
rect 191465 298011 191531 298012
rect 266353 298011 266419 298014
rect 267774 298012 267780 298014
rect 267844 298074 267850 298076
rect 272057 298074 272123 298077
rect 267844 298072 272123 298074
rect 267844 298016 272062 298072
rect 272118 298016 272123 298072
rect 267844 298014 272123 298016
rect 267844 298012 267850 298014
rect 272057 298011 272123 298014
rect 256601 297938 256667 297941
rect 253460 297936 256667 297938
rect 253460 297880 256606 297936
rect 256662 297880 256667 297936
rect 253460 297878 256667 297880
rect 256601 297875 256667 297878
rect 256509 297530 256575 297533
rect 253460 297528 256575 297530
rect 253460 297472 256514 297528
rect 256570 297472 256575 297528
rect 253460 297470 256575 297472
rect 256509 297467 256575 297470
rect 16481 297394 16547 297397
rect 192702 297394 192708 297396
rect 16481 297392 192708 297394
rect 16481 297336 16486 297392
rect 16542 297336 192708 297392
rect 16481 297334 192708 297336
rect 16481 297331 16547 297334
rect 192702 297332 192708 297334
rect 192772 297332 192778 297396
rect 191741 297122 191807 297125
rect 255865 297122 255931 297125
rect 191741 297120 193660 297122
rect 191741 297064 191746 297120
rect 191802 297064 193660 297120
rect 191741 297062 193660 297064
rect 253460 297120 255931 297122
rect 253460 297064 255870 297120
rect 255926 297064 255931 297120
rect 253460 297062 255931 297064
rect 191741 297059 191807 297062
rect 255865 297059 255931 297062
rect 252829 296986 252895 296989
rect 253197 296986 253263 296989
rect 252829 296984 253263 296986
rect 252829 296928 252834 296984
rect 252890 296928 253202 296984
rect 253258 296928 253263 296984
rect 252829 296926 253263 296928
rect 252829 296923 252895 296926
rect 253197 296923 253263 296926
rect 256601 296986 256667 296989
rect 264881 296986 264947 296989
rect 256601 296984 264947 296986
rect 256601 296928 256606 296984
rect 256662 296928 264886 296984
rect 264942 296928 264947 296984
rect 256601 296926 264947 296928
rect 256601 296923 256667 296926
rect 264881 296923 264947 296926
rect 280429 296714 280495 296717
rect 253460 296712 280495 296714
rect 253460 296656 280434 296712
rect 280490 296656 280495 296712
rect 253460 296654 280495 296656
rect 280429 296651 280495 296654
rect 252829 296578 252895 296581
rect 253013 296578 253079 296581
rect 252829 296576 253079 296578
rect 252829 296520 252834 296576
rect 252890 296520 253018 296576
rect 253074 296520 253079 296576
rect 252829 296518 253079 296520
rect 252829 296515 252938 296518
rect 253013 296515 253079 296518
rect 252878 296276 252938 296515
rect 193029 296170 193095 296173
rect 193029 296168 193660 296170
rect 193029 296112 193034 296168
rect 193090 296112 193660 296168
rect 193029 296110 193660 296112
rect 193029 296107 193095 296110
rect 255262 295898 255268 295900
rect 253460 295838 255268 295898
rect 255262 295836 255268 295838
rect 255332 295836 255338 295900
rect 256601 295490 256667 295493
rect 253460 295488 256667 295490
rect 253460 295432 256606 295488
rect 256662 295432 256667 295488
rect 253460 295430 256667 295432
rect 256601 295427 256667 295430
rect 268326 295292 268332 295356
rect 268396 295354 268402 295356
rect 269113 295354 269179 295357
rect 268396 295352 269179 295354
rect 268396 295296 269118 295352
rect 269174 295296 269179 295352
rect 268396 295294 269179 295296
rect 268396 295292 268402 295294
rect 269113 295291 269179 295294
rect 280429 295354 280495 295357
rect 284477 295354 284543 295357
rect 280429 295352 284543 295354
rect 280429 295296 280434 295352
rect 280490 295296 284482 295352
rect 284538 295296 284543 295352
rect 280429 295294 284543 295296
rect 280429 295291 280495 295294
rect 284477 295291 284543 295294
rect 192477 295218 192543 295221
rect 193305 295218 193371 295221
rect 278865 295218 278931 295221
rect 192477 295216 193660 295218
rect 192477 295160 192482 295216
rect 192538 295160 193310 295216
rect 193366 295160 193660 295216
rect 192477 295158 193660 295160
rect 263550 295216 278931 295218
rect 263550 295160 278870 295216
rect 278926 295160 278931 295216
rect 263550 295158 278931 295160
rect 192477 295155 192543 295158
rect 193305 295155 193371 295158
rect 255589 295082 255655 295085
rect 256601 295082 256667 295085
rect 253460 295080 256667 295082
rect 253460 295024 255594 295080
rect 255650 295024 256606 295080
rect 256662 295024 256667 295080
rect 253460 295022 256667 295024
rect 255589 295019 255655 295022
rect 256601 295019 256667 295022
rect 263550 294946 263610 295158
rect 278865 295155 278931 295158
rect 253430 294886 263610 294946
rect 253430 294644 253490 294886
rect 79961 294538 80027 294541
rect 87086 294538 87092 294540
rect 79961 294536 87092 294538
rect 79961 294480 79966 294536
rect 80022 294480 87092 294536
rect 79961 294478 87092 294480
rect 79961 294475 80027 294478
rect 87086 294476 87092 294478
rect 87156 294476 87162 294540
rect 93761 294538 93827 294541
rect 98310 294538 98316 294540
rect 93761 294536 98316 294538
rect 93761 294480 93766 294536
rect 93822 294480 98316 294536
rect 93761 294478 98316 294480
rect 93761 294475 93827 294478
rect 98310 294476 98316 294478
rect 98380 294476 98386 294540
rect 120717 294538 120783 294541
rect 189993 294538 190059 294541
rect 120717 294536 190059 294538
rect 120717 294480 120722 294536
rect 120778 294480 189998 294536
rect 190054 294480 190059 294536
rect 120717 294478 190059 294480
rect 120717 294475 120783 294478
rect 189993 294475 190059 294478
rect 191741 294266 191807 294269
rect 256601 294266 256667 294269
rect 191741 294264 193660 294266
rect 191741 294208 191746 294264
rect 191802 294208 193660 294264
rect 191741 294206 193660 294208
rect 253460 294264 256667 294266
rect 253460 294208 256606 294264
rect 256662 294208 256667 294264
rect 253460 294206 256667 294208
rect 191741 294203 191807 294206
rect 256601 294203 256667 294206
rect 75678 293932 75684 293996
rect 75748 293994 75754 293996
rect 176653 293994 176719 293997
rect 177205 293994 177271 293997
rect 75748 293992 177271 293994
rect 75748 293936 176658 293992
rect 176714 293936 177210 293992
rect 177266 293936 177271 293992
rect 75748 293934 177271 293936
rect 75748 293932 75754 293934
rect 176653 293931 176719 293934
rect 177205 293931 177271 293934
rect 278865 293994 278931 293997
rect 285673 293994 285739 293997
rect 278865 293992 285739 293994
rect 278865 293936 278870 293992
rect 278926 293936 285678 293992
rect 285734 293936 285739 293992
rect 278865 293934 285739 293936
rect 278865 293931 278931 293934
rect 285673 293931 285739 293934
rect 255497 293858 255563 293861
rect 253460 293856 255563 293858
rect 253460 293800 255502 293856
rect 255558 293800 255563 293856
rect 253460 293798 255563 293800
rect 255497 293795 255563 293798
rect 255681 293450 255747 293453
rect 253460 293448 255747 293450
rect 253460 293392 255686 293448
rect 255742 293392 255747 293448
rect 253460 293390 255747 293392
rect 255681 293387 255747 293390
rect -960 293178 480 293268
rect 3417 293178 3483 293181
rect -960 293176 3483 293178
rect -960 293120 3422 293176
rect 3478 293120 3483 293176
rect -960 293118 3483 293120
rect -960 293028 480 293118
rect 3417 293115 3483 293118
rect 155309 293178 155375 293181
rect 191966 293178 191972 293180
rect 155309 293176 191972 293178
rect 155309 293120 155314 293176
rect 155370 293120 191972 293176
rect 155309 293118 191972 293120
rect 155309 293115 155375 293118
rect 191966 293116 191972 293118
rect 192036 293116 192042 293180
rect 192702 293116 192708 293180
rect 192772 293178 192778 293180
rect 192772 293118 193660 293178
rect 192772 293116 192778 293118
rect 256601 293042 256667 293045
rect 253460 293040 256667 293042
rect 253460 292984 256606 293040
rect 256662 292984 256667 293040
rect 253460 292982 256667 292984
rect 256601 292979 256667 292982
rect 86534 292572 86540 292636
rect 86604 292634 86610 292636
rect 91093 292634 91159 292637
rect 86604 292632 91159 292634
rect 86604 292576 91098 292632
rect 91154 292576 91159 292632
rect 86604 292574 91159 292576
rect 86604 292572 86610 292574
rect 91093 292571 91159 292574
rect 191741 292634 191807 292637
rect 192702 292634 192708 292636
rect 191741 292632 192708 292634
rect 191741 292576 191746 292632
rect 191802 292576 192708 292632
rect 191741 292574 192708 292576
rect 191741 292571 191807 292574
rect 192702 292572 192708 292574
rect 192772 292572 192778 292636
rect 255405 292634 255471 292637
rect 253460 292632 255471 292634
rect 253460 292576 255410 292632
rect 255466 292576 255471 292632
rect 253460 292574 255471 292576
rect 255405 292571 255471 292574
rect 191741 292226 191807 292229
rect 255405 292226 255471 292229
rect 191741 292224 193660 292226
rect 191741 292168 191746 292224
rect 191802 292168 193660 292224
rect 191741 292166 193660 292168
rect 253460 292224 255471 292226
rect 253460 292168 255410 292224
rect 255466 292168 255471 292224
rect 253460 292166 255471 292168
rect 191741 292163 191807 292166
rect 255405 292163 255471 292166
rect 83089 291954 83155 291957
rect 92974 291954 92980 291956
rect 83089 291952 92980 291954
rect 83089 291896 83094 291952
rect 83150 291896 92980 291952
rect 83089 291894 92980 291896
rect 83089 291891 83155 291894
rect 92974 291892 92980 291894
rect 93044 291954 93050 291956
rect 100017 291954 100083 291957
rect 93044 291952 100083 291954
rect 93044 291896 100022 291952
rect 100078 291896 100083 291952
rect 93044 291894 100083 291896
rect 93044 291892 93050 291894
rect 100017 291891 100083 291894
rect 178677 291954 178743 291957
rect 183461 291954 183527 291957
rect 178677 291952 183527 291954
rect 178677 291896 178682 291952
rect 178738 291896 183466 291952
rect 183522 291896 183527 291952
rect 178677 291894 183527 291896
rect 178677 291891 178743 291894
rect 183461 291891 183527 291894
rect 64597 291818 64663 291821
rect 80145 291818 80211 291821
rect 64597 291816 80211 291818
rect 64597 291760 64602 291816
rect 64658 291760 80150 291816
rect 80206 291760 80211 291816
rect 64597 291758 80211 291760
rect 64597 291755 64663 291758
rect 80145 291755 80211 291758
rect 83958 291756 83964 291820
rect 84028 291818 84034 291820
rect 106457 291818 106523 291821
rect 84028 291816 106523 291818
rect 84028 291760 106462 291816
rect 106518 291760 106523 291816
rect 84028 291758 106523 291760
rect 84028 291756 84034 291758
rect 106457 291755 106523 291758
rect 134609 291818 134675 291821
rect 181529 291818 181595 291821
rect 257061 291818 257127 291821
rect 267917 291818 267983 291821
rect 134609 291816 181595 291818
rect 134609 291760 134614 291816
rect 134670 291760 181534 291816
rect 181590 291760 181595 291816
rect 134609 291758 181595 291760
rect 253460 291816 257127 291818
rect 253460 291760 257066 291816
rect 257122 291760 257127 291816
rect 253460 291758 257127 291760
rect 134609 291755 134675 291758
rect 181529 291755 181595 291758
rect 257061 291755 257127 291758
rect 258030 291816 267983 291818
rect 258030 291760 267922 291816
rect 267978 291760 267983 291816
rect 258030 291758 267983 291760
rect 258030 291682 258090 291758
rect 267917 291755 267983 291758
rect 253430 291622 258090 291682
rect 80881 291274 80947 291277
rect 83958 291274 83964 291276
rect 80881 291272 83964 291274
rect 80881 291216 80886 291272
rect 80942 291216 83964 291272
rect 80881 291214 83964 291216
rect 80881 291211 80947 291214
rect 83958 291212 83964 291214
rect 84028 291212 84034 291276
rect 85849 291274 85915 291277
rect 86769 291274 86835 291277
rect 104157 291274 104223 291277
rect 191557 291276 191623 291277
rect 191557 291274 191604 291276
rect 85849 291272 104223 291274
rect 85849 291216 85854 291272
rect 85910 291216 86774 291272
rect 86830 291216 104162 291272
rect 104218 291216 104223 291272
rect 85849 291214 104223 291216
rect 191476 291272 191604 291274
rect 191668 291274 191674 291276
rect 191476 291216 191562 291272
rect 191476 291214 191604 291216
rect 85849 291211 85915 291214
rect 86769 291211 86835 291214
rect 104157 291211 104223 291214
rect 191557 291212 191604 291214
rect 191668 291214 193660 291274
rect 253430 291244 253490 291622
rect 191668 291212 191674 291214
rect 191557 291211 191623 291212
rect 255405 290866 255471 290869
rect 253460 290864 255471 290866
rect 253460 290808 255410 290864
rect 255466 290808 255471 290864
rect 253460 290806 255471 290808
rect 255405 290803 255471 290806
rect 262438 290730 262444 290732
rect 253430 290670 262444 290730
rect 83181 290458 83247 290461
rect 92606 290458 92612 290460
rect 83181 290456 92612 290458
rect 83181 290400 83186 290456
rect 83242 290400 92612 290456
rect 83181 290398 92612 290400
rect 83181 290395 83247 290398
rect 92606 290396 92612 290398
rect 92676 290396 92682 290460
rect 166441 290458 166507 290461
rect 184841 290458 184907 290461
rect 166441 290456 184907 290458
rect 166441 290400 166446 290456
rect 166502 290400 184846 290456
rect 184902 290400 184907 290456
rect 253430 290428 253490 290670
rect 262438 290668 262444 290670
rect 262508 290730 262514 290732
rect 263593 290730 263659 290733
rect 262508 290728 263659 290730
rect 262508 290672 263598 290728
rect 263654 290672 263659 290728
rect 262508 290670 263659 290672
rect 262508 290668 262514 290670
rect 263593 290667 263659 290670
rect 166441 290398 184907 290400
rect 166441 290395 166507 290398
rect 184841 290395 184907 290398
rect 191741 290322 191807 290325
rect 191741 290320 193660 290322
rect 191741 290264 191746 290320
rect 191802 290264 193660 290320
rect 191741 290262 193660 290264
rect 191741 290259 191807 290262
rect 73286 289988 73292 290052
rect 73356 290050 73362 290052
rect 74533 290050 74599 290053
rect 73356 290048 74599 290050
rect 73356 289992 74538 290048
rect 74594 289992 74599 290048
rect 73356 289990 74599 289992
rect 73356 289988 73362 289990
rect 74533 289987 74599 289990
rect 82629 290050 82695 290053
rect 104893 290050 104959 290053
rect 256785 290050 256851 290053
rect 82629 290048 104959 290050
rect 82629 289992 82634 290048
rect 82690 289992 104898 290048
rect 104954 289992 104959 290048
rect 82629 289990 104959 289992
rect 253460 290048 256851 290050
rect 253460 289992 256790 290048
rect 256846 289992 256851 290048
rect 253460 289990 256851 289992
rect 82629 289987 82695 289990
rect 104893 289987 104959 289990
rect 256785 289987 256851 289990
rect 73153 289914 73219 289917
rect 73470 289914 73476 289916
rect 73153 289912 73476 289914
rect 73153 289856 73158 289912
rect 73214 289856 73476 289912
rect 73153 289854 73476 289856
rect 73153 289851 73219 289854
rect 73470 289852 73476 289854
rect 73540 289852 73546 289916
rect 90909 289914 90975 289917
rect 166441 289914 166507 289917
rect 253197 289914 253263 289917
rect 90909 289912 166507 289914
rect 90909 289856 90914 289912
rect 90970 289856 166446 289912
rect 166502 289856 166507 289912
rect 90909 289854 166507 289856
rect 90909 289851 90975 289854
rect 166441 289851 166507 289854
rect 252878 289912 253263 289914
rect 252878 289856 253202 289912
rect 253258 289856 253263 289912
rect 252878 289854 253263 289856
rect 252878 289778 252938 289854
rect 253197 289851 253263 289854
rect 252878 289718 253490 289778
rect 253430 289642 253490 289718
rect 253841 289642 253907 289645
rect 253430 289640 253907 289642
rect 253430 289612 253846 289640
rect 253460 289584 253846 289612
rect 253902 289584 253907 289640
rect 253460 289582 253907 289584
rect 253841 289579 253907 289582
rect 252870 289444 252876 289508
rect 252940 289444 252946 289508
rect 191557 289370 191623 289373
rect 191557 289368 193660 289370
rect 191557 289312 191562 289368
rect 191618 289312 193660 289368
rect 191557 289310 193660 289312
rect 191557 289307 191623 289310
rect 55121 289234 55187 289237
rect 79317 289234 79383 289237
rect 55121 289232 79383 289234
rect 55121 289176 55126 289232
rect 55182 289176 79322 289232
rect 79378 289176 79383 289232
rect 55121 289174 79383 289176
rect 55121 289171 55187 289174
rect 79317 289171 79383 289174
rect 79685 289098 79751 289101
rect 120165 289098 120231 289101
rect 156597 289098 156663 289101
rect 169753 289098 169819 289101
rect 79685 289096 169819 289098
rect 79685 289040 79690 289096
rect 79746 289040 120170 289096
rect 120226 289040 156602 289096
rect 156658 289040 169758 289096
rect 169814 289040 169819 289096
rect 79685 289038 169819 289040
rect 252878 289098 252938 289444
rect 270769 289098 270835 289101
rect 252878 289096 270835 289098
rect 252878 289040 270774 289096
rect 270830 289040 270835 289096
rect 252878 289038 270835 289040
rect 79685 289035 79751 289038
rect 120165 289035 120231 289038
rect 156597 289035 156663 289038
rect 169753 289035 169819 289038
rect 270769 289035 270835 289038
rect 255497 288826 255563 288829
rect 253460 288824 255563 288826
rect 253460 288768 255502 288824
rect 255558 288768 255563 288824
rect 253460 288766 255563 288768
rect 255497 288763 255563 288766
rect 65793 288418 65859 288421
rect 66069 288418 66135 288421
rect 65793 288416 66135 288418
rect 65793 288360 65798 288416
rect 65854 288360 66074 288416
rect 66130 288360 66135 288416
rect 65793 288358 66135 288360
rect 65793 288355 65859 288358
rect 66069 288355 66135 288358
rect 191741 288418 191807 288421
rect 191741 288416 193660 288418
rect 191741 288360 191746 288416
rect 191802 288360 193660 288416
rect 191741 288358 193660 288360
rect 191741 288355 191807 288358
rect 253430 288282 253490 288388
rect 263869 288282 263935 288285
rect 253430 288280 263935 288282
rect 253430 288224 263874 288280
rect 263930 288224 263935 288280
rect 253430 288222 263935 288224
rect 263869 288219 263935 288222
rect 253430 287874 253490 287980
rect 253430 287814 258090 287874
rect 129089 287738 129155 287741
rect 141509 287738 141575 287741
rect 129089 287736 141575 287738
rect 129089 287680 129094 287736
rect 129150 287680 141514 287736
rect 141570 287680 141575 287736
rect 129089 287678 141575 287680
rect 129089 287675 129155 287678
rect 141509 287675 141575 287678
rect 255313 287602 255379 287605
rect 253460 287600 255379 287602
rect 253460 287544 255318 287600
rect 255374 287544 255379 287600
rect 253460 287542 255379 287544
rect 255313 287539 255379 287542
rect 86401 287466 86467 287469
rect 86861 287466 86927 287469
rect 100109 287466 100175 287469
rect 86401 287464 100175 287466
rect 86401 287408 86406 287464
rect 86462 287408 86866 287464
rect 86922 287408 100114 287464
rect 100170 287408 100175 287464
rect 86401 287406 100175 287408
rect 86401 287403 86467 287406
rect 86861 287403 86927 287406
rect 100109 287403 100175 287406
rect 190637 287466 190703 287469
rect 258030 287466 258090 287814
rect 270585 287466 270651 287469
rect 278865 287466 278931 287469
rect 190637 287464 193660 287466
rect 190637 287408 190642 287464
rect 190698 287408 193660 287464
rect 190637 287406 193660 287408
rect 258030 287464 278931 287466
rect 258030 287408 270590 287464
rect 270646 287408 278870 287464
rect 278926 287408 278931 287464
rect 258030 287406 278931 287408
rect 190637 287403 190703 287406
rect 270585 287403 270651 287406
rect 278865 287403 278931 287406
rect 66069 287330 66135 287333
rect 98494 287330 98500 287332
rect 66069 287328 98500 287330
rect 66069 287272 66074 287328
rect 66130 287272 98500 287328
rect 66069 287270 98500 287272
rect 66069 287267 66135 287270
rect 98494 287268 98500 287270
rect 98564 287268 98570 287332
rect 95785 287194 95851 287197
rect 129089 287194 129155 287197
rect 255497 287194 255563 287197
rect 95785 287192 129155 287194
rect 95785 287136 95790 287192
rect 95846 287136 129094 287192
rect 129150 287136 129155 287192
rect 95785 287134 129155 287136
rect 253460 287192 255563 287194
rect 253460 287136 255502 287192
rect 255558 287136 255563 287192
rect 253460 287134 255563 287136
rect 95785 287131 95851 287134
rect 129089 287131 129155 287134
rect 255497 287131 255563 287134
rect 72049 287058 72115 287061
rect 73061 287058 73127 287061
rect 157241 287058 157307 287061
rect 270493 287058 270559 287061
rect 72049 287056 157307 287058
rect 72049 287000 72054 287056
rect 72110 287000 73066 287056
rect 73122 287000 157246 287056
rect 157302 287000 157307 287056
rect 72049 286998 157307 287000
rect 72049 286995 72115 286998
rect 73061 286995 73127 286998
rect 157241 286995 157307 286998
rect 253430 287056 270559 287058
rect 253430 287000 270498 287056
rect 270554 287000 270559 287056
rect 253430 286998 270559 287000
rect 253430 286756 253490 286998
rect 270493 286995 270559 286998
rect 191005 286514 191071 286517
rect 191005 286512 193660 286514
rect 191005 286456 191010 286512
rect 191066 286456 193660 286512
rect 191005 286454 193660 286456
rect 191005 286451 191071 286454
rect 255497 286378 255563 286381
rect 253460 286376 255563 286378
rect 253460 286320 255502 286376
rect 255558 286320 255563 286376
rect 253460 286318 255563 286320
rect 255497 286315 255563 286318
rect 255405 285970 255471 285973
rect 253460 285968 255471 285970
rect 253460 285912 255410 285968
rect 255466 285912 255471 285968
rect 253460 285910 255471 285912
rect 255405 285907 255471 285910
rect 75913 285834 75979 285837
rect 64830 285832 75979 285834
rect 64830 285776 75918 285832
rect 75974 285776 75979 285832
rect 64830 285774 75979 285776
rect 61837 285698 61903 285701
rect 64830 285698 64890 285774
rect 75913 285771 75979 285774
rect 91921 285834 91987 285837
rect 157241 285834 157307 285837
rect 160921 285834 160987 285837
rect 91921 285832 99390 285834
rect 91921 285776 91926 285832
rect 91982 285776 99390 285832
rect 91921 285774 99390 285776
rect 91921 285771 91987 285774
rect 61837 285696 64890 285698
rect 61837 285640 61842 285696
rect 61898 285640 64890 285696
rect 61837 285638 64890 285640
rect 87505 285698 87571 285701
rect 90909 285698 90975 285701
rect 87505 285696 90975 285698
rect 87505 285640 87510 285696
rect 87566 285640 90914 285696
rect 90970 285640 90975 285696
rect 87505 285638 90975 285640
rect 61837 285635 61903 285638
rect 87505 285635 87571 285638
rect 90909 285635 90975 285638
rect 93853 285698 93919 285701
rect 98678 285698 98684 285700
rect 93853 285696 98684 285698
rect 93853 285640 93858 285696
rect 93914 285640 98684 285696
rect 93853 285638 98684 285640
rect 93853 285635 93919 285638
rect 98678 285636 98684 285638
rect 98748 285636 98754 285700
rect 99330 285698 99390 285774
rect 157241 285832 160987 285834
rect 157241 285776 157246 285832
rect 157302 285776 160926 285832
rect 160982 285776 160987 285832
rect 157241 285774 160987 285776
rect 157241 285771 157307 285774
rect 160921 285771 160987 285774
rect 102133 285698 102199 285701
rect 102961 285698 103027 285701
rect 99330 285696 103027 285698
rect 99330 285640 102138 285696
rect 102194 285640 102966 285696
rect 103022 285640 103027 285696
rect 99330 285638 103027 285640
rect 102133 285635 102199 285638
rect 102961 285635 103027 285638
rect 113817 285562 113883 285565
rect 181437 285562 181503 285565
rect 113817 285560 181503 285562
rect 113817 285504 113822 285560
rect 113878 285504 181442 285560
rect 181498 285504 181503 285560
rect 113817 285502 181503 285504
rect 113817 285499 113883 285502
rect 181437 285499 181503 285502
rect 191649 285562 191715 285565
rect 255405 285562 255471 285565
rect 263685 285562 263751 285565
rect 191649 285560 193660 285562
rect 191649 285504 191654 285560
rect 191710 285504 193660 285560
rect 255405 285560 263751 285562
rect 191649 285502 193660 285504
rect 191649 285499 191715 285502
rect 252829 285426 252895 285429
rect 253430 285426 253490 285532
rect 255405 285504 255410 285560
rect 255466 285504 263690 285560
rect 263746 285504 263751 285560
rect 255405 285502 263751 285504
rect 255405 285499 255471 285502
rect 263685 285499 263751 285502
rect 265341 285426 265407 285429
rect 252829 285424 252938 285426
rect 252829 285368 252834 285424
rect 252890 285368 252938 285424
rect 252829 285363 252938 285368
rect 253430 285424 265407 285426
rect 253430 285368 265346 285424
rect 265402 285368 265407 285424
rect 253430 285366 265407 285368
rect 265341 285363 265407 285366
rect 252878 285124 252938 285363
rect 583520 285276 584960 285516
rect 76005 284882 76071 284885
rect 76414 284882 76420 284884
rect 76005 284880 76420 284882
rect 76005 284824 76010 284880
rect 76066 284824 76420 284880
rect 76005 284822 76420 284824
rect 76005 284819 76071 284822
rect 76414 284820 76420 284822
rect 76484 284882 76490 284884
rect 100293 284882 100359 284885
rect 76484 284880 100359 284882
rect 76484 284824 100298 284880
rect 100354 284824 100359 284880
rect 76484 284822 100359 284824
rect 76484 284820 76490 284822
rect 100293 284819 100359 284822
rect 256877 284746 256943 284749
rect 253460 284744 256943 284746
rect 253460 284688 256882 284744
rect 256938 284688 256943 284744
rect 253460 284686 256943 284688
rect 256877 284683 256943 284686
rect 89161 284474 89227 284477
rect 89621 284474 89687 284477
rect 111149 284474 111215 284477
rect 89161 284472 111215 284474
rect 89161 284416 89166 284472
rect 89222 284416 89626 284472
rect 89682 284416 111154 284472
rect 111210 284416 111215 284472
rect 89161 284414 111215 284416
rect 89161 284411 89227 284414
rect 89621 284411 89687 284414
rect 111149 284411 111215 284414
rect 191741 284474 191807 284477
rect 191741 284472 193660 284474
rect 191741 284416 191746 284472
rect 191802 284416 193660 284472
rect 191741 284414 193660 284416
rect 191741 284411 191807 284414
rect 70158 284276 70164 284340
rect 70228 284338 70234 284340
rect 72417 284338 72483 284341
rect 70228 284336 72483 284338
rect 70228 284280 72422 284336
rect 72478 284280 72483 284336
rect 70228 284278 72483 284280
rect 70228 284276 70234 284278
rect 72417 284275 72483 284278
rect 72918 284276 72924 284340
rect 72988 284338 72994 284340
rect 74901 284338 74967 284341
rect 72988 284336 74967 284338
rect 72988 284280 74906 284336
rect 74962 284280 74967 284336
rect 72988 284278 74967 284280
rect 72988 284276 72994 284278
rect 74901 284275 74967 284278
rect 97441 284338 97507 284341
rect 178861 284338 178927 284341
rect 97441 284336 178927 284338
rect 97441 284280 97446 284336
rect 97502 284280 178866 284336
rect 178922 284280 178927 284336
rect 97441 284278 178927 284280
rect 97441 284275 97507 284278
rect 178861 284275 178927 284278
rect 191097 284338 191163 284341
rect 191649 284338 191715 284341
rect 255405 284338 255471 284341
rect 191097 284336 191715 284338
rect 191097 284280 191102 284336
rect 191158 284280 191654 284336
rect 191710 284280 191715 284336
rect 191097 284278 191715 284280
rect 253460 284336 255471 284338
rect 253460 284280 255410 284336
rect 255466 284280 255471 284336
rect 253460 284278 255471 284280
rect 191097 284275 191163 284278
rect 191649 284275 191715 284278
rect 255405 284275 255471 284278
rect 265341 284338 265407 284341
rect 266353 284338 266419 284341
rect 265341 284336 266419 284338
rect 265341 284280 265346 284336
rect 265402 284280 266358 284336
rect 266414 284280 266419 284336
rect 265341 284278 266419 284280
rect 265341 284275 265407 284278
rect 266353 284275 266419 284278
rect 73153 284204 73219 284205
rect 73102 284202 73108 284204
rect 73062 284142 73108 284202
rect 73172 284200 73219 284204
rect 73214 284144 73219 284200
rect 73102 284140 73108 284142
rect 73172 284140 73219 284144
rect 87086 284140 87092 284204
rect 87156 284202 87162 284204
rect 87597 284202 87663 284205
rect 87156 284200 87663 284202
rect 87156 284144 87602 284200
rect 87658 284144 87663 284200
rect 87156 284142 87663 284144
rect 87156 284140 87162 284142
rect 73153 284139 73219 284140
rect 87597 284139 87663 284142
rect 253657 283930 253723 283933
rect 253460 283928 253723 283930
rect 253460 283872 253662 283928
rect 253718 283872 253723 283928
rect 253460 283870 253723 283872
rect 253657 283867 253723 283870
rect 67081 283794 67147 283797
rect 67541 283794 67607 283797
rect 67081 283792 67607 283794
rect 67081 283736 67086 283792
rect 67142 283736 67546 283792
rect 67602 283736 67607 283792
rect 67081 283734 67607 283736
rect 67081 283731 67147 283734
rect 67541 283731 67607 283734
rect 68553 283522 68619 283525
rect 69381 283522 69447 283525
rect 69974 283522 69980 283524
rect 68553 283520 69980 283522
rect 68553 283464 68558 283520
rect 68614 283464 69386 283520
rect 69442 283464 69980 283520
rect 68553 283462 69980 283464
rect 68553 283459 68619 283462
rect 69381 283459 69447 283462
rect 69974 283460 69980 283462
rect 70044 283460 70050 283524
rect 71313 283522 71379 283525
rect 71630 283522 71636 283524
rect 71313 283520 71636 283522
rect 71313 283464 71318 283520
rect 71374 283464 71636 283520
rect 71313 283462 71636 283464
rect 71313 283459 71379 283462
rect 71630 283460 71636 283462
rect 71700 283460 71706 283524
rect 88609 283522 88675 283525
rect 89478 283522 89484 283524
rect 88609 283520 89484 283522
rect 88609 283464 88614 283520
rect 88670 283464 89484 283520
rect 88609 283462 89484 283464
rect 88609 283459 88675 283462
rect 89478 283460 89484 283462
rect 89548 283460 89554 283524
rect 193029 283522 193095 283525
rect 258165 283522 258231 283525
rect 266445 283522 266511 283525
rect 193029 283520 193660 283522
rect 193029 283464 193034 283520
rect 193090 283464 193660 283520
rect 193029 283462 193660 283464
rect 253460 283520 266511 283522
rect 253460 283464 258170 283520
rect 258226 283464 266450 283520
rect 266506 283464 266511 283520
rect 253460 283462 266511 283464
rect 193029 283459 193095 283462
rect 258165 283459 258231 283462
rect 266445 283459 266511 283462
rect 68686 283324 68692 283388
rect 68756 283386 68762 283388
rect 69749 283386 69815 283389
rect 83457 283388 83523 283389
rect 83406 283386 83412 283388
rect 68756 283384 69815 283386
rect 68756 283328 69754 283384
rect 69810 283328 69815 283384
rect 68756 283326 69815 283328
rect 83366 283326 83412 283386
rect 83476 283384 83523 283388
rect 83518 283328 83523 283384
rect 68756 283324 68762 283326
rect 69749 283323 69815 283326
rect 83406 283324 83412 283326
rect 83476 283324 83523 283328
rect 83457 283323 83523 283324
rect 3509 283250 3575 283253
rect 87086 283250 87092 283252
rect 3509 283248 87092 283250
rect 3509 283192 3514 283248
rect 3570 283192 87092 283248
rect 3509 283190 87092 283192
rect 3509 283187 3575 283190
rect 87086 283188 87092 283190
rect 87156 283188 87162 283252
rect 69974 283052 69980 283116
rect 70044 283114 70050 283116
rect 71037 283114 71103 283117
rect 70044 283112 71103 283114
rect 70044 283056 71042 283112
rect 71098 283056 71103 283112
rect 70044 283054 71103 283056
rect 70044 283052 70050 283054
rect 71037 283051 71103 283054
rect 75361 283114 75427 283117
rect 75678 283114 75684 283116
rect 75361 283112 75684 283114
rect 75361 283056 75366 283112
rect 75422 283056 75684 283112
rect 75361 283054 75684 283056
rect 75361 283051 75427 283054
rect 75678 283052 75684 283054
rect 75748 283052 75754 283116
rect 97901 283114 97967 283117
rect 117957 283114 118023 283117
rect 255497 283114 255563 283117
rect 97901 283112 118023 283114
rect 97901 283056 97906 283112
rect 97962 283056 117962 283112
rect 118018 283056 118023 283112
rect 97901 283054 118023 283056
rect 253460 283112 255563 283114
rect 253460 283056 255502 283112
rect 255558 283056 255563 283112
rect 253460 283054 255563 283056
rect 97901 283051 97967 283054
rect 117957 283051 118023 283054
rect 255497 283051 255563 283054
rect 66805 282978 66871 282981
rect 85297 282978 85363 282981
rect 188337 282978 188403 282981
rect 66805 282976 68908 282978
rect 66805 282920 66810 282976
rect 66866 282920 68908 282976
rect 66805 282918 68908 282920
rect 85297 282976 188403 282978
rect 85297 282920 85302 282976
rect 85358 282920 188342 282976
rect 188398 282920 188403 282976
rect 85297 282918 188403 282920
rect 66805 282915 66871 282918
rect 85297 282915 85363 282918
rect 188337 282915 188403 282918
rect 98913 282842 98979 282845
rect 161381 282842 161447 282845
rect 162301 282842 162367 282845
rect 98913 282840 162367 282842
rect 98913 282784 98918 282840
rect 98974 282784 161386 282840
rect 161442 282784 162306 282840
rect 162362 282784 162367 282840
rect 98913 282782 162367 282784
rect 98913 282779 98979 282782
rect 161381 282779 161447 282782
rect 162301 282779 162367 282782
rect 100753 282706 100819 282709
rect 255497 282706 255563 282709
rect 98716 282704 100819 282706
rect 98716 282648 100758 282704
rect 100814 282648 100819 282704
rect 98716 282646 100819 282648
rect 253460 282704 255563 282706
rect 253460 282648 255502 282704
rect 255558 282648 255563 282704
rect 253460 282646 255563 282648
rect 100753 282643 100819 282646
rect 255497 282643 255563 282646
rect 191557 282570 191623 282573
rect 191557 282568 193660 282570
rect 191557 282512 191562 282568
rect 191618 282512 193660 282568
rect 191557 282510 193660 282512
rect 191557 282507 191623 282510
rect 67081 282162 67147 282165
rect 253430 282162 253490 282268
rect 277577 282162 277643 282165
rect 67081 282160 68908 282162
rect 67081 282104 67086 282160
rect 67142 282104 68908 282160
rect 67081 282102 68908 282104
rect 253430 282160 277643 282162
rect 253430 282104 277582 282160
rect 277638 282104 277643 282160
rect 253430 282102 277643 282104
rect 67081 282099 67147 282102
rect 277577 282099 277643 282102
rect 255405 281890 255471 281893
rect 253460 281888 255471 281890
rect 67265 281618 67331 281621
rect 67398 281618 67404 281620
rect 67265 281616 67404 281618
rect 67265 281560 67270 281616
rect 67326 281560 67404 281616
rect 67265 281558 67404 281560
rect 67265 281555 67331 281558
rect 67398 281556 67404 281558
rect 67468 281556 67474 281620
rect 98686 281618 98746 281860
rect 253460 281832 255410 281888
rect 255466 281832 255471 281888
rect 253460 281830 255471 281832
rect 255405 281827 255471 281830
rect 113817 281618 113883 281621
rect 98686 281616 113883 281618
rect 98686 281560 113822 281616
rect 113878 281560 113883 281616
rect 98686 281558 113883 281560
rect 113817 281555 113883 281558
rect 162301 281618 162367 281621
rect 168465 281618 168531 281621
rect 162301 281616 168531 281618
rect 162301 281560 162306 281616
rect 162362 281560 168470 281616
rect 168526 281560 168531 281616
rect 162301 281558 168531 281560
rect 162301 281555 162367 281558
rect 168465 281555 168531 281558
rect 191741 281618 191807 281621
rect 191741 281616 193660 281618
rect 191741 281560 191746 281616
rect 191802 281560 193660 281616
rect 191741 281558 193660 281560
rect 191741 281555 191807 281558
rect 66529 281482 66595 281485
rect 68277 281482 68343 281485
rect 66529 281480 68938 281482
rect 66529 281424 66534 281480
rect 66590 281424 68282 281480
rect 68338 281424 68938 281480
rect 66529 281422 68938 281424
rect 66529 281419 66595 281422
rect 68277 281419 68343 281422
rect 68878 281316 68938 281422
rect 255405 281346 255471 281349
rect 253460 281344 255471 281346
rect 253460 281288 255410 281344
rect 255466 281288 255471 281344
rect 253460 281286 255471 281288
rect 255405 281283 255471 281286
rect 100845 281074 100911 281077
rect 98716 281072 100911 281074
rect 98716 281016 100850 281072
rect 100906 281016 100911 281072
rect 98716 281014 100911 281016
rect 100845 281011 100911 281014
rect 258809 280938 258875 280941
rect 268326 280938 268332 280940
rect 258809 280936 268332 280938
rect 151169 280802 151235 280805
rect 184197 280802 184263 280805
rect 151169 280800 184263 280802
rect 151169 280744 151174 280800
rect 151230 280744 184202 280800
rect 184258 280744 184263 280800
rect 151169 280742 184263 280744
rect 253430 280802 253490 280908
rect 258809 280880 258814 280936
rect 258870 280880 268332 280936
rect 258809 280878 268332 280880
rect 258809 280875 258875 280878
rect 268326 280876 268332 280878
rect 268396 280876 268402 280940
rect 258257 280802 258323 280805
rect 274909 280802 274975 280805
rect 253430 280800 274975 280802
rect 253430 280744 258262 280800
rect 258318 280744 274914 280800
rect 274970 280744 274975 280800
rect 253430 280742 274975 280744
rect 151169 280739 151235 280742
rect 184197 280739 184263 280742
rect 258257 280739 258323 280742
rect 274909 280739 274975 280742
rect 191281 280666 191347 280669
rect 192937 280666 193003 280669
rect 191281 280664 193660 280666
rect 191281 280608 191286 280664
rect 191342 280608 192942 280664
rect 192998 280608 193660 280664
rect 191281 280606 193660 280608
rect 191281 280603 191347 280606
rect 192937 280603 193003 280606
rect 66897 280530 66963 280533
rect 255405 280530 255471 280533
rect 66897 280528 68908 280530
rect 66897 280472 66902 280528
rect 66958 280472 68908 280528
rect 66897 280470 68908 280472
rect 253460 280528 255471 280530
rect 253460 280472 255410 280528
rect 255466 280472 255471 280528
rect 253460 280470 255471 280472
rect 66897 280467 66963 280470
rect 255405 280467 255471 280470
rect 100753 280258 100819 280261
rect 98716 280256 100819 280258
rect -960 279972 480 280212
rect 98716 280200 100758 280256
rect 100814 280200 100819 280256
rect 98716 280198 100819 280200
rect 100753 280195 100819 280198
rect 255405 280122 255471 280125
rect 253460 280120 255471 280122
rect 253460 280064 255410 280120
rect 255466 280064 255471 280120
rect 253460 280062 255471 280064
rect 255405 280059 255471 280062
rect 67541 279714 67607 279717
rect 191557 279714 191623 279717
rect 258717 279714 258783 279717
rect 67541 279712 68908 279714
rect 67541 279656 67546 279712
rect 67602 279656 68908 279712
rect 67541 279654 68908 279656
rect 191557 279712 193660 279714
rect 191557 279656 191562 279712
rect 191618 279656 193660 279712
rect 191557 279654 193660 279656
rect 253460 279712 258783 279714
rect 253460 279656 258722 279712
rect 258778 279656 258783 279712
rect 253460 279654 258783 279656
rect 67541 279651 67607 279654
rect 191557 279651 191623 279654
rect 258717 279651 258783 279654
rect 100753 279442 100819 279445
rect 98716 279440 100819 279442
rect 98716 279384 100758 279440
rect 100814 279384 100819 279440
rect 98716 279382 100819 279384
rect 100753 279379 100819 279382
rect 256693 279306 256759 279309
rect 253460 279304 256759 279306
rect 253460 279248 256698 279304
rect 256754 279248 256759 279304
rect 253460 279246 256759 279248
rect 256693 279243 256759 279246
rect 66621 278898 66687 278901
rect 255497 278898 255563 278901
rect 66621 278896 68908 278898
rect 66621 278840 66626 278896
rect 66682 278840 68908 278896
rect 66621 278838 68908 278840
rect 253460 278896 255563 278898
rect 253460 278840 255502 278896
rect 255558 278840 255563 278896
rect 253460 278838 255563 278840
rect 66621 278835 66687 278838
rect 255497 278835 255563 278838
rect 193121 278762 193187 278765
rect 193397 278762 193463 278765
rect 193121 278760 193660 278762
rect 193121 278704 193126 278760
rect 193182 278704 193402 278760
rect 193458 278704 193660 278760
rect 193121 278702 193660 278704
rect 193121 278699 193187 278702
rect 193397 278699 193463 278702
rect 101673 278626 101739 278629
rect 98716 278624 101739 278626
rect 98716 278568 101678 278624
rect 101734 278568 101739 278624
rect 98716 278566 101739 278568
rect 101673 278563 101739 278566
rect 253430 278354 253490 278460
rect 266629 278354 266695 278357
rect 253430 278352 267750 278354
rect 253430 278296 266634 278352
rect 266690 278296 267750 278352
rect 253430 278294 267750 278296
rect 266629 278291 266695 278294
rect 66805 278082 66871 278085
rect 66805 278080 68908 278082
rect 66805 278024 66810 278080
rect 66866 278024 68908 278080
rect 66805 278022 68908 278024
rect 66805 278019 66871 278022
rect 253430 277946 253490 278052
rect 263685 277946 263751 277949
rect 253430 277944 263751 277946
rect 253430 277888 263690 277944
rect 263746 277888 263751 277944
rect 253430 277886 263751 277888
rect 267690 277946 267750 278294
rect 276197 277946 276263 277949
rect 267690 277944 276263 277946
rect 267690 277888 276202 277944
rect 276258 277888 276263 277944
rect 267690 277886 276263 277888
rect 263685 277883 263751 277886
rect 276197 277883 276263 277886
rect 100753 277810 100819 277813
rect 98716 277808 100819 277810
rect 98716 277752 100758 277808
rect 100814 277752 100819 277808
rect 98716 277750 100819 277752
rect 100753 277747 100819 277750
rect 192845 277810 192911 277813
rect 192845 277808 193660 277810
rect 192845 277752 192850 277808
rect 192906 277752 193660 277808
rect 192845 277750 193660 277752
rect 192845 277747 192911 277750
rect 255405 277674 255471 277677
rect 253460 277672 255471 277674
rect 253460 277616 255410 277672
rect 255466 277616 255471 277672
rect 253460 277614 255471 277616
rect 255405 277611 255471 277614
rect 67357 277266 67423 277269
rect 259545 277266 259611 277269
rect 262305 277266 262371 277269
rect 67357 277264 68908 277266
rect 67357 277208 67362 277264
rect 67418 277208 68908 277264
rect 67357 277206 68908 277208
rect 253460 277264 262371 277266
rect 253460 277208 259550 277264
rect 259606 277208 262310 277264
rect 262366 277208 262371 277264
rect 253460 277206 262371 277208
rect 67357 277203 67423 277206
rect 259545 277203 259611 277206
rect 262305 277203 262371 277206
rect 101489 276994 101555 276997
rect 98716 276992 101555 276994
rect 98716 276936 101494 276992
rect 101550 276936 101555 276992
rect 98716 276934 101555 276936
rect 101489 276931 101555 276934
rect 193213 276858 193279 276861
rect 258073 276858 258139 276861
rect 260966 276858 260972 276860
rect 193213 276856 193660 276858
rect 193213 276800 193218 276856
rect 193274 276800 193660 276856
rect 193213 276798 193660 276800
rect 253460 276856 260972 276858
rect 253460 276800 258078 276856
rect 258134 276800 260972 276856
rect 253460 276798 260972 276800
rect 193213 276795 193279 276798
rect 258073 276795 258139 276798
rect 260966 276796 260972 276798
rect 261036 276796 261042 276860
rect 100845 276722 100911 276725
rect 128997 276722 129063 276725
rect 100845 276720 129063 276722
rect 100845 276664 100850 276720
rect 100906 276664 129002 276720
rect 129058 276664 129063 276720
rect 100845 276662 129063 276664
rect 100845 276659 100911 276662
rect 128997 276659 129063 276662
rect 66897 276450 66963 276453
rect 255405 276450 255471 276453
rect 66897 276448 68908 276450
rect 66897 276392 66902 276448
rect 66958 276392 68908 276448
rect 66897 276390 68908 276392
rect 253460 276448 255471 276450
rect 253460 276392 255410 276448
rect 255466 276392 255471 276448
rect 253460 276390 255471 276392
rect 66897 276387 66963 276390
rect 255405 276387 255471 276390
rect 100753 276178 100819 276181
rect 98716 276176 100819 276178
rect 98716 276120 100758 276176
rect 100814 276120 100819 276176
rect 98716 276118 100819 276120
rect 100753 276115 100819 276118
rect 255497 276042 255563 276045
rect 253460 276040 255563 276042
rect 253460 275984 255502 276040
rect 255558 275984 255563 276040
rect 253460 275982 255563 275984
rect 255497 275979 255563 275982
rect 66161 275634 66227 275637
rect 66161 275632 68908 275634
rect 66161 275576 66166 275632
rect 66222 275576 68908 275632
rect 66161 275574 68908 275576
rect 66161 275571 66227 275574
rect 66069 274818 66135 274821
rect 98686 274818 98746 275332
rect 193630 275090 193690 275740
rect 256734 275634 256740 275636
rect 253460 275574 256740 275634
rect 256734 275572 256740 275574
rect 256804 275572 256810 275636
rect 255405 275226 255471 275229
rect 253460 275224 255471 275226
rect 253460 275168 255410 275224
rect 255466 275168 255471 275224
rect 253460 275166 255471 275168
rect 255405 275163 255471 275166
rect 190870 275030 193690 275090
rect 149881 274818 149947 274821
rect 66069 274816 68908 274818
rect 66069 274760 66074 274816
rect 66130 274760 68908 274816
rect 66069 274758 68908 274760
rect 98686 274816 149947 274818
rect 98686 274760 149886 274816
rect 149942 274760 149947 274816
rect 98686 274758 149947 274760
rect 66069 274755 66135 274758
rect 149881 274755 149947 274758
rect 190310 274620 190316 274684
rect 190380 274682 190386 274684
rect 190870 274682 190930 275030
rect 191189 274818 191255 274821
rect 191557 274818 191623 274821
rect 255405 274818 255471 274821
rect 191189 274816 193660 274818
rect 191189 274760 191194 274816
rect 191250 274760 191562 274816
rect 191618 274760 193660 274816
rect 191189 274758 193660 274760
rect 253460 274816 255471 274818
rect 253460 274760 255410 274816
rect 255466 274760 255471 274816
rect 253460 274758 255471 274760
rect 191189 274755 191255 274758
rect 191557 274755 191623 274758
rect 255405 274755 255471 274758
rect 190380 274622 190930 274682
rect 190380 274620 190386 274622
rect 101489 274546 101555 274549
rect 98716 274544 101555 274546
rect 98716 274488 101494 274544
rect 101550 274488 101555 274544
rect 98716 274486 101555 274488
rect 101489 274483 101555 274486
rect 255405 274410 255471 274413
rect 253460 274408 255471 274410
rect 253460 274352 255410 274408
rect 255466 274352 255471 274408
rect 253460 274350 255471 274352
rect 255405 274347 255471 274350
rect 66529 274002 66595 274005
rect 255497 274002 255563 274005
rect 66529 274000 68908 274002
rect 66529 273944 66534 274000
rect 66590 273944 68908 274000
rect 66529 273942 68908 273944
rect 253460 274000 255563 274002
rect 253460 273944 255502 274000
rect 255558 273944 255563 274000
rect 253460 273942 255563 273944
rect 66529 273939 66595 273942
rect 255497 273939 255563 273942
rect 141509 273866 141575 273869
rect 180241 273866 180307 273869
rect 260925 273866 260991 273869
rect 270585 273866 270651 273869
rect 141509 273864 180307 273866
rect 141509 273808 141514 273864
rect 141570 273808 180246 273864
rect 180302 273808 180307 273864
rect 258030 273864 270651 273866
rect 141509 273806 180307 273808
rect 141509 273803 141575 273806
rect 180241 273803 180307 273806
rect 100753 273730 100819 273733
rect 98716 273728 100819 273730
rect 98716 273672 100758 273728
rect 100814 273672 100819 273728
rect 98716 273670 100819 273672
rect 100753 273667 100819 273670
rect 188838 273260 188844 273324
rect 188908 273322 188914 273324
rect 193630 273322 193690 273836
rect 258030 273808 260930 273864
rect 260986 273808 270590 273864
rect 270646 273808 270651 273864
rect 258030 273806 270651 273808
rect 253430 273458 253490 273564
rect 258030 273458 258090 273806
rect 260925 273803 260991 273806
rect 270585 273803 270651 273806
rect 253430 273398 258090 273458
rect 188908 273262 193690 273322
rect 188908 273260 188914 273262
rect 67398 273124 67404 273188
rect 67468 273186 67474 273188
rect 255405 273186 255471 273189
rect 67468 273126 68908 273186
rect 253460 273184 255471 273186
rect 253460 273128 255410 273184
rect 255466 273128 255471 273184
rect 253460 273126 255471 273128
rect 67468 273124 67474 273126
rect 255405 273123 255471 273126
rect 259453 273186 259519 273189
rect 260046 273186 260052 273188
rect 259453 273184 260052 273186
rect 259453 273128 259458 273184
rect 259514 273128 260052 273184
rect 259453 273126 260052 273128
rect 259453 273123 259519 273126
rect 260046 273124 260052 273126
rect 260116 273124 260122 273188
rect 100753 272914 100819 272917
rect 98716 272912 100819 272914
rect 98716 272856 100758 272912
rect 100814 272856 100819 272912
rect 98716 272854 100819 272856
rect 100753 272851 100819 272854
rect 191649 272914 191715 272917
rect 191649 272912 193660 272914
rect 191649 272856 191654 272912
rect 191710 272856 193660 272912
rect 191649 272854 193660 272856
rect 191649 272851 191715 272854
rect 255497 272778 255563 272781
rect 253460 272776 255563 272778
rect 253460 272720 255502 272776
rect 255558 272720 255563 272776
rect 253460 272718 255563 272720
rect 255497 272715 255563 272718
rect 161105 272506 161171 272509
rect 189717 272506 189783 272509
rect 161105 272504 189783 272506
rect 161105 272448 161110 272504
rect 161166 272448 189722 272504
rect 189778 272448 189783 272504
rect 161105 272446 189783 272448
rect 161105 272443 161171 272446
rect 189717 272443 189783 272446
rect 66621 272370 66687 272373
rect 66621 272368 68908 272370
rect 66621 272312 66626 272368
rect 66682 272312 68908 272368
rect 66621 272310 68908 272312
rect 66621 272307 66687 272310
rect 253430 272234 253490 272340
rect 267733 272234 267799 272237
rect 270493 272234 270559 272237
rect 253430 272232 270559 272234
rect 253430 272176 267738 272232
rect 267794 272176 270498 272232
rect 270554 272176 270559 272232
rect 253430 272174 270559 272176
rect 267733 272171 267799 272174
rect 270493 272171 270559 272174
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 100845 272098 100911 272101
rect 98716 272096 100911 272098
rect 98716 272040 100850 272096
rect 100906 272040 100911 272096
rect 583520 272084 584960 272174
rect 98716 272038 100911 272040
rect 100845 272035 100911 272038
rect 191741 271962 191807 271965
rect 256877 271962 256943 271965
rect 191741 271960 193660 271962
rect 191741 271904 191746 271960
rect 191802 271904 193660 271960
rect 191741 271902 193660 271904
rect 253460 271960 256943 271962
rect 253460 271904 256882 271960
rect 256938 271904 256943 271960
rect 253460 271902 256943 271904
rect 191741 271899 191807 271902
rect 256877 271899 256943 271902
rect 66253 271554 66319 271557
rect 66253 271552 68908 271554
rect 66253 271496 66258 271552
rect 66314 271496 68908 271552
rect 66253 271494 68908 271496
rect 66253 271491 66319 271494
rect 255405 271418 255471 271421
rect 253460 271416 255471 271418
rect 253460 271360 255410 271416
rect 255466 271360 255471 271416
rect 253460 271358 255471 271360
rect 255405 271355 255471 271358
rect 100753 271282 100819 271285
rect 98716 271280 100819 271282
rect 98716 271224 100758 271280
rect 100814 271224 100819 271280
rect 98716 271222 100819 271224
rect 100753 271219 100819 271222
rect 98678 271084 98684 271148
rect 98748 271146 98754 271148
rect 152549 271146 152615 271149
rect 281717 271146 281783 271149
rect 98748 271144 152615 271146
rect 98748 271088 152554 271144
rect 152610 271088 152615 271144
rect 98748 271086 152615 271088
rect 98748 271084 98754 271086
rect 152549 271083 152615 271086
rect 267690 271144 281783 271146
rect 267690 271088 281722 271144
rect 281778 271088 281783 271144
rect 267690 271086 281783 271088
rect 191741 271010 191807 271013
rect 191741 271008 193660 271010
rect 191741 270952 191746 271008
rect 191802 270952 193660 271008
rect 191741 270950 193660 270952
rect 191741 270947 191807 270950
rect 253430 270874 253490 270980
rect 263777 270874 263843 270877
rect 267690 270874 267750 271086
rect 281717 271083 281783 271086
rect 253430 270872 267750 270874
rect 253430 270816 263782 270872
rect 263838 270816 267750 270872
rect 253430 270814 267750 270816
rect 263777 270811 263843 270814
rect 60457 270738 60523 270741
rect 60457 270736 68908 270738
rect 60457 270680 60462 270736
rect 60518 270680 68908 270736
rect 60457 270678 68908 270680
rect 60457 270675 60523 270678
rect 106089 270602 106155 270605
rect 129181 270602 129247 270605
rect 255405 270602 255471 270605
rect 106089 270600 129247 270602
rect 106089 270544 106094 270600
rect 106150 270544 129186 270600
rect 129242 270544 129247 270600
rect 106089 270542 129247 270544
rect 253460 270600 255471 270602
rect 253460 270544 255410 270600
rect 255466 270544 255471 270600
rect 253460 270542 255471 270544
rect 106089 270539 106155 270542
rect 129181 270539 129247 270542
rect 255405 270539 255471 270542
rect 258257 270602 258323 270605
rect 258390 270602 258396 270604
rect 258257 270600 258396 270602
rect 258257 270544 258262 270600
rect 258318 270544 258396 270600
rect 258257 270542 258396 270544
rect 258257 270539 258323 270542
rect 258390 270540 258396 270542
rect 258460 270540 258466 270604
rect 100753 270466 100819 270469
rect 98716 270464 100819 270466
rect 98716 270408 100758 270464
rect 100814 270408 100819 270464
rect 98716 270406 100819 270408
rect 100753 270403 100819 270406
rect 255497 270194 255563 270197
rect 253460 270192 255563 270194
rect 253460 270136 255502 270192
rect 255558 270136 255563 270192
rect 253460 270134 255563 270136
rect 255497 270131 255563 270134
rect 190821 270058 190887 270061
rect 190821 270056 193660 270058
rect 190821 270000 190826 270056
rect 190882 270000 193660 270056
rect 190821 269998 193660 270000
rect 190821 269995 190887 269998
rect 68878 269378 68938 269892
rect 100017 269786 100083 269789
rect 142981 269786 143047 269789
rect 100017 269784 143047 269786
rect 100017 269728 100022 269784
rect 100078 269728 142986 269784
rect 143042 269728 143047 269784
rect 100017 269726 143047 269728
rect 100017 269723 100083 269726
rect 142981 269723 143047 269726
rect 158621 269786 158687 269789
rect 172605 269786 172671 269789
rect 255405 269786 255471 269789
rect 158621 269784 172671 269786
rect 158621 269728 158626 269784
rect 158682 269728 172610 269784
rect 172666 269728 172671 269784
rect 158621 269726 172671 269728
rect 253460 269784 255471 269786
rect 253460 269728 255410 269784
rect 255466 269728 255471 269784
rect 253460 269726 255471 269728
rect 158621 269723 158687 269726
rect 172605 269723 172671 269726
rect 255405 269723 255471 269726
rect 257337 269786 257403 269789
rect 291653 269786 291719 269789
rect 257337 269784 291719 269786
rect 257337 269728 257342 269784
rect 257398 269728 291658 269784
rect 291714 269728 291719 269784
rect 257337 269726 291719 269728
rect 257337 269723 257403 269726
rect 291653 269723 291719 269726
rect 101581 269650 101647 269653
rect 98716 269648 101647 269650
rect 98716 269592 101586 269648
rect 101642 269592 101647 269648
rect 98716 269590 101647 269592
rect 101581 269587 101647 269590
rect 256693 269378 256759 269381
rect 259494 269378 259500 269380
rect 64830 269318 68938 269378
rect 253460 269376 259500 269378
rect 253460 269320 256698 269376
rect 256754 269320 259500 269376
rect 253460 269318 259500 269320
rect 60641 269242 60707 269245
rect 64830 269242 64890 269318
rect 256693 269315 256759 269318
rect 259494 269316 259500 269318
rect 259564 269316 259570 269380
rect 60641 269240 64890 269242
rect 60641 269184 60646 269240
rect 60702 269184 64890 269240
rect 60641 269182 64890 269184
rect 60641 269179 60707 269182
rect 66897 269106 66963 269109
rect 191465 269106 191531 269109
rect 66897 269104 68908 269106
rect 66897 269048 66902 269104
rect 66958 269048 68908 269104
rect 66897 269046 68908 269048
rect 191465 269104 193660 269106
rect 191465 269048 191470 269104
rect 191526 269048 193660 269104
rect 191465 269046 193660 269048
rect 66897 269043 66963 269046
rect 191465 269043 191531 269046
rect 255405 268970 255471 268973
rect 253460 268968 255471 268970
rect 253460 268912 255410 268968
rect 255466 268912 255471 268968
rect 253460 268910 255471 268912
rect 255405 268907 255471 268910
rect 100753 268834 100819 268837
rect 98716 268832 100819 268834
rect 98716 268776 100758 268832
rect 100814 268776 100819 268832
rect 98716 268774 100819 268776
rect 100753 268771 100819 268774
rect 140037 268562 140103 268565
rect 188286 268562 188292 268564
rect 140037 268560 188292 268562
rect 140037 268504 140042 268560
rect 140098 268504 188292 268560
rect 140037 268502 188292 268504
rect 140037 268499 140103 268502
rect 188286 268500 188292 268502
rect 188356 268500 188362 268564
rect 100293 268426 100359 268429
rect 159541 268426 159607 268429
rect 100293 268424 159607 268426
rect 100293 268368 100298 268424
rect 100354 268368 159546 268424
rect 159602 268368 159607 268424
rect 100293 268366 159607 268368
rect 253430 268426 253490 268532
rect 277393 268426 277459 268429
rect 253430 268424 277459 268426
rect 253430 268368 277398 268424
rect 277454 268368 277459 268424
rect 253430 268366 277459 268368
rect 100293 268363 100359 268366
rect 159541 268363 159607 268366
rect 66805 268290 66871 268293
rect 66805 268288 68908 268290
rect 66805 268232 66810 268288
rect 66866 268232 68908 268288
rect 66805 268230 68908 268232
rect 66805 268227 66871 268230
rect 191741 268154 191807 268157
rect 255497 268154 255563 268157
rect 191741 268152 193660 268154
rect 191741 268096 191746 268152
rect 191802 268096 193660 268152
rect 191741 268094 193660 268096
rect 253460 268152 255563 268154
rect 253460 268096 255502 268152
rect 255558 268096 255563 268152
rect 253460 268094 255563 268096
rect 191741 268091 191807 268094
rect 255497 268091 255563 268094
rect 100753 268018 100819 268021
rect 98716 268016 100819 268018
rect 98716 267960 100758 268016
rect 100814 267960 100819 268016
rect 98716 267958 100819 267960
rect 267690 268018 267750 268366
rect 277393 268363 277459 268366
rect 268009 268018 268075 268021
rect 267690 268016 268075 268018
rect 267690 267960 268014 268016
rect 268070 267960 268075 268016
rect 267690 267958 268075 267960
rect 100753 267955 100819 267958
rect 268009 267955 268075 267958
rect 100109 267882 100175 267885
rect 104985 267882 105051 267885
rect 100109 267880 105051 267882
rect 100109 267824 100114 267880
rect 100170 267824 104990 267880
rect 105046 267824 105051 267880
rect 100109 267822 105051 267824
rect 100109 267819 100175 267822
rect 104985 267819 105051 267822
rect 255497 267746 255563 267749
rect 253460 267744 255563 267746
rect 253460 267688 255502 267744
rect 255558 267688 255563 267744
rect 253460 267686 255563 267688
rect 255497 267683 255563 267686
rect 66621 267474 66687 267477
rect 66621 267472 68908 267474
rect 66621 267416 66626 267472
rect 66682 267416 68908 267472
rect 66621 267414 68908 267416
rect 66621 267411 66687 267414
rect -960 267202 480 267292
rect 3509 267202 3575 267205
rect 100753 267202 100819 267205
rect -960 267200 3575 267202
rect -960 267144 3514 267200
rect 3570 267144 3575 267200
rect -960 267142 3575 267144
rect 98716 267200 100819 267202
rect 98716 267144 100758 267200
rect 100814 267144 100819 267200
rect 98716 267142 100819 267144
rect -960 267052 480 267142
rect 3509 267139 3575 267142
rect 100753 267139 100819 267142
rect 137369 267202 137435 267205
rect 184054 267202 184060 267204
rect 137369 267200 184060 267202
rect 137369 267144 137374 267200
rect 137430 267144 184060 267200
rect 137369 267142 184060 267144
rect 137369 267139 137435 267142
rect 184054 267140 184060 267142
rect 184124 267140 184130 267204
rect 253430 267202 253490 267308
rect 253430 267142 258090 267202
rect 98862 267004 98868 267068
rect 98932 267066 98938 267068
rect 155953 267066 156019 267069
rect 156413 267066 156479 267069
rect 98932 267064 156479 267066
rect 98932 267008 155958 267064
rect 156014 267008 156418 267064
rect 156474 267008 156479 267064
rect 98932 267006 156479 267008
rect 98932 267004 98938 267006
rect 155953 267003 156019 267006
rect 156413 267003 156479 267006
rect 191741 267066 191807 267069
rect 191741 267064 193660 267066
rect 191741 267008 191746 267064
rect 191802 267008 193660 267064
rect 191741 267006 193660 267008
rect 191741 267003 191807 267006
rect 255405 266930 255471 266933
rect 253460 266928 255471 266930
rect 253460 266872 255410 266928
rect 255466 266872 255471 266928
rect 253460 266870 255471 266872
rect 255405 266867 255471 266870
rect 258030 266794 258090 267142
rect 266813 267068 266879 267069
rect 266813 267064 266860 267068
rect 266924 267066 266930 267068
rect 266813 267008 266818 267064
rect 266813 267004 266860 267008
rect 266924 267006 266970 267066
rect 266924 267004 266930 267006
rect 266813 267003 266879 267004
rect 276238 266794 276244 266796
rect 258030 266734 276244 266794
rect 276238 266732 276244 266734
rect 276308 266794 276314 266796
rect 277393 266794 277459 266797
rect 276308 266792 277459 266794
rect 276308 266736 277398 266792
rect 277454 266736 277459 266792
rect 276308 266734 277459 266736
rect 276308 266732 276314 266734
rect 277393 266731 277459 266734
rect 66437 266658 66503 266661
rect 66437 266656 68908 266658
rect 66437 266600 66442 266656
rect 66498 266600 68908 266656
rect 66437 266598 68908 266600
rect 66437 266595 66503 266598
rect 252878 266389 252938 266492
rect 100937 266386 101003 266389
rect 98716 266384 101003 266386
rect 98716 266328 100942 266384
rect 100998 266328 101003 266384
rect 98716 266326 101003 266328
rect 252878 266384 252987 266389
rect 252878 266328 252926 266384
rect 252982 266328 252987 266384
rect 252878 266326 252987 266328
rect 100937 266323 101003 266326
rect 252921 266323 252987 266326
rect 190821 266114 190887 266117
rect 255497 266114 255563 266117
rect 190821 266112 193660 266114
rect 190821 266056 190826 266112
rect 190882 266056 193660 266112
rect 190821 266054 193660 266056
rect 253460 266112 255563 266114
rect 253460 266056 255502 266112
rect 255558 266056 255563 266112
rect 253460 266054 255563 266056
rect 190821 266051 190887 266054
rect 255497 266051 255563 266054
rect 66805 265842 66871 265845
rect 66805 265840 68908 265842
rect 66805 265784 66810 265840
rect 66866 265784 68908 265840
rect 66805 265782 68908 265784
rect 66805 265779 66871 265782
rect 259729 265706 259795 265709
rect 253460 265704 259795 265706
rect 253460 265648 259734 265704
rect 259790 265648 259795 265704
rect 253460 265646 259795 265648
rect 259729 265643 259795 265646
rect 100753 265570 100819 265573
rect 98716 265568 100819 265570
rect 98716 265512 100758 265568
rect 100814 265512 100819 265568
rect 98716 265510 100819 265512
rect 100753 265507 100819 265510
rect 187601 265570 187667 265573
rect 193438 265570 193444 265572
rect 187601 265568 193444 265570
rect 187601 265512 187606 265568
rect 187662 265512 193444 265568
rect 187601 265510 193444 265512
rect 187601 265507 187667 265510
rect 193438 265508 193444 265510
rect 193508 265508 193514 265572
rect 259269 265570 259335 265573
rect 272149 265570 272215 265573
rect 259269 265568 272215 265570
rect 259269 265512 259274 265568
rect 259330 265512 272154 265568
rect 272210 265512 272215 265568
rect 259269 265510 272215 265512
rect 259269 265507 259335 265510
rect 272149 265507 272215 265510
rect 255405 265298 255471 265301
rect 253460 265296 255471 265298
rect 253460 265240 255410 265296
rect 255466 265240 255471 265296
rect 253460 265238 255471 265240
rect 255405 265235 255471 265238
rect 61929 265162 61995 265165
rect 63125 265162 63191 265165
rect 162117 265162 162183 265165
rect 61929 265160 68938 265162
rect 61929 265104 61934 265160
rect 61990 265104 63130 265160
rect 63186 265104 68938 265160
rect 61929 265102 68938 265104
rect 61929 265099 61995 265102
rect 63125 265099 63191 265102
rect 68878 264996 68938 265102
rect 162117 265160 193660 265162
rect 162117 265104 162122 265160
rect 162178 265104 193660 265160
rect 162117 265102 193660 265104
rect 162117 265099 162183 265102
rect 181437 265026 181503 265029
rect 187049 265026 187115 265029
rect 181437 265024 187115 265026
rect 181437 264968 181442 265024
rect 181498 264968 187054 265024
rect 187110 264968 187115 265024
rect 181437 264966 187115 264968
rect 181437 264963 181503 264966
rect 187049 264963 187115 264966
rect 255589 264890 255655 264893
rect 253460 264888 255655 264890
rect 253460 264832 255594 264888
rect 255650 264832 255655 264888
rect 253460 264830 255655 264832
rect 255589 264827 255655 264830
rect 267181 264890 267247 264893
rect 269062 264890 269068 264892
rect 267181 264888 269068 264890
rect 267181 264832 267186 264888
rect 267242 264832 269068 264888
rect 267181 264830 269068 264832
rect 267181 264827 267247 264830
rect 269062 264828 269068 264830
rect 269132 264828 269138 264892
rect 100845 264754 100911 264757
rect 98716 264752 100911 264754
rect 98716 264696 100850 264752
rect 100906 264696 100911 264752
rect 98716 264694 100911 264696
rect 100845 264691 100911 264694
rect 255405 264482 255471 264485
rect 253460 264480 255471 264482
rect 253460 264424 255410 264480
rect 255466 264424 255471 264480
rect 253460 264422 255471 264424
rect 255405 264419 255471 264422
rect 66805 264210 66871 264213
rect 191741 264210 191807 264213
rect 281574 264210 281580 264212
rect 66805 264208 68908 264210
rect 66805 264152 66810 264208
rect 66866 264152 68908 264208
rect 66805 264150 68908 264152
rect 191741 264208 193660 264210
rect 191741 264152 191746 264208
rect 191802 264152 193660 264208
rect 191741 264150 193660 264152
rect 267690 264150 281580 264210
rect 66805 264147 66871 264150
rect 191741 264147 191807 264150
rect 255405 264074 255471 264077
rect 253460 264072 255471 264074
rect 253460 264016 255410 264072
rect 255466 264016 255471 264072
rect 253460 264014 255471 264016
rect 255405 264011 255471 264014
rect 100753 263938 100819 263941
rect 98716 263936 100819 263938
rect 98716 263880 100758 263936
rect 100814 263880 100819 263936
rect 98716 263878 100819 263880
rect 100753 263875 100819 263878
rect 255497 263802 255563 263805
rect 263869 263802 263935 263805
rect 267690 263802 267750 264150
rect 281574 264148 281580 264150
rect 281644 264148 281650 264212
rect 255497 263800 267750 263802
rect 255497 263744 255502 263800
rect 255558 263744 263874 263800
rect 263930 263744 267750 263800
rect 255497 263742 267750 263744
rect 255497 263739 255563 263742
rect 263869 263739 263935 263742
rect 262438 263666 262444 263668
rect 253460 263606 262444 263666
rect 262438 263604 262444 263606
rect 262508 263604 262514 263668
rect 269849 263666 269915 263669
rect 270718 263666 270724 263668
rect 269849 263664 270724 263666
rect 269849 263608 269854 263664
rect 269910 263608 270724 263664
rect 269849 263606 270724 263608
rect 269849 263603 269915 263606
rect 270718 263604 270724 263606
rect 270788 263666 270794 263668
rect 276238 263666 276244 263668
rect 270788 263606 276244 263666
rect 270788 263604 270794 263606
rect 276238 263604 276244 263606
rect 276308 263604 276314 263668
rect 67081 263394 67147 263397
rect 67449 263394 67515 263397
rect 67081 263392 68908 263394
rect 67081 263336 67086 263392
rect 67142 263336 67454 263392
rect 67510 263336 68908 263392
rect 67081 263334 68908 263336
rect 67081 263331 67147 263334
rect 67449 263331 67515 263334
rect 191005 263258 191071 263261
rect 254117 263258 254183 263261
rect 255037 263258 255103 263261
rect 191005 263256 193660 263258
rect 191005 263200 191010 263256
rect 191066 263200 193660 263256
rect 191005 263198 193660 263200
rect 253460 263256 255103 263258
rect 253460 263200 254122 263256
rect 254178 263200 255042 263256
rect 255098 263200 255103 263256
rect 253460 263198 255103 263200
rect 191005 263195 191071 263198
rect 254117 263195 254183 263198
rect 255037 263195 255103 263198
rect 100753 263122 100819 263125
rect 98716 263120 100819 263122
rect 98716 263064 100758 263120
rect 100814 263064 100819 263120
rect 98716 263062 100819 263064
rect 100753 263059 100819 263062
rect 100937 262850 101003 262853
rect 163681 262850 163747 262853
rect 100937 262848 163747 262850
rect 100937 262792 100942 262848
rect 100998 262792 163686 262848
rect 163742 262792 163747 262848
rect 100937 262790 163747 262792
rect 100937 262787 101003 262790
rect 163681 262787 163747 262790
rect 253430 262714 253490 262820
rect 266486 262714 266492 262716
rect 253430 262654 266492 262714
rect 266486 262652 266492 262654
rect 266556 262652 266562 262716
rect 66897 262578 66963 262581
rect 66897 262576 68908 262578
rect 66897 262520 66902 262576
rect 66958 262520 68908 262576
rect 66897 262518 68908 262520
rect 66897 262515 66963 262518
rect 255497 262442 255563 262445
rect 253460 262440 255563 262442
rect 253460 262384 255502 262440
rect 255558 262384 255563 262440
rect 253460 262382 255563 262384
rect 255497 262379 255563 262382
rect 100753 262306 100819 262309
rect 98716 262304 100819 262306
rect 98716 262248 100758 262304
rect 100814 262248 100819 262304
rect 98716 262246 100819 262248
rect 100753 262243 100819 262246
rect 191741 262306 191807 262309
rect 191741 262304 193660 262306
rect 191741 262248 191746 262304
rect 191802 262248 193660 262304
rect 191741 262246 193660 262248
rect 191741 262243 191807 262246
rect 66253 261762 66319 261765
rect 253430 261762 253490 262004
rect 263542 261762 263548 261764
rect 66253 261760 68908 261762
rect 66253 261704 66258 261760
rect 66314 261704 68908 261760
rect 66253 261702 68908 261704
rect 253430 261702 263548 261762
rect 66253 261699 66319 261702
rect 263542 261700 263548 261702
rect 263612 261700 263618 261764
rect 50797 261490 50863 261493
rect 64781 261490 64847 261493
rect 100845 261492 100911 261493
rect 100845 261490 100892 261492
rect 50797 261488 68938 261490
rect 50797 261432 50802 261488
rect 50858 261432 64786 261488
rect 64842 261432 68938 261488
rect 50797 261430 68938 261432
rect 98716 261488 100892 261490
rect 100956 261490 100962 261492
rect 137277 261490 137343 261493
rect 173014 261490 173020 261492
rect 98716 261432 100850 261488
rect 98716 261430 100892 261432
rect 50797 261427 50863 261430
rect 64781 261427 64847 261430
rect 68878 260916 68938 261430
rect 100845 261428 100892 261430
rect 100956 261430 101038 261490
rect 137277 261488 173020 261490
rect 137277 261432 137282 261488
rect 137338 261432 173020 261488
rect 137277 261430 173020 261432
rect 100956 261428 100962 261430
rect 100845 261427 100911 261428
rect 137277 261427 137343 261430
rect 173014 261428 173020 261430
rect 173084 261428 173090 261492
rect 191557 261354 191623 261357
rect 253430 261354 253490 261460
rect 263726 261354 263732 261356
rect 191557 261352 193660 261354
rect 191557 261296 191562 261352
rect 191618 261296 193660 261352
rect 191557 261294 193660 261296
rect 253430 261294 263732 261354
rect 191557 261291 191623 261294
rect 263726 261292 263732 261294
rect 263796 261292 263802 261356
rect 254526 261082 254532 261084
rect 253460 261022 254532 261082
rect 254526 261020 254532 261022
rect 254596 261020 254602 261084
rect 100845 260674 100911 260677
rect 255262 260674 255268 260676
rect 98716 260672 100911 260674
rect 98716 260616 100850 260672
rect 100906 260616 100911 260672
rect 98716 260614 100911 260616
rect 253460 260614 255268 260674
rect 100845 260611 100911 260614
rect 255262 260612 255268 260614
rect 255332 260674 255338 260676
rect 255405 260674 255471 260677
rect 255332 260672 255471 260674
rect 255332 260616 255410 260672
rect 255466 260616 255471 260672
rect 255332 260614 255471 260616
rect 255332 260612 255338 260614
rect 255405 260611 255471 260614
rect 191741 260402 191807 260405
rect 191741 260400 193660 260402
rect 191741 260344 191746 260400
rect 191802 260344 193660 260400
rect 191741 260342 193660 260344
rect 191741 260339 191807 260342
rect 255589 260266 255655 260269
rect 253460 260264 255655 260266
rect 253460 260208 255594 260264
rect 255650 260208 255655 260264
rect 253460 260206 255655 260208
rect 255589 260203 255655 260206
rect 41229 260130 41295 260133
rect 66805 260130 66871 260133
rect 41229 260128 66871 260130
rect 41229 260072 41234 260128
rect 41290 260072 66810 260128
rect 66866 260072 66871 260128
rect 111149 260130 111215 260133
rect 170765 260130 170831 260133
rect 111149 260128 170831 260130
rect 41229 260070 66871 260072
rect 41229 260067 41295 260070
rect 66805 260067 66871 260070
rect 65885 259586 65951 259589
rect 68878 259586 68938 260100
rect 111149 260072 111154 260128
rect 111210 260072 170770 260128
rect 170826 260072 170831 260128
rect 111149 260070 170831 260072
rect 111149 260067 111215 260070
rect 170765 260067 170831 260070
rect 100753 259858 100819 259861
rect 259494 259858 259500 259860
rect 98716 259856 100819 259858
rect 98716 259800 100758 259856
rect 100814 259800 100819 259856
rect 98716 259798 100819 259800
rect 253460 259798 259500 259858
rect 100753 259795 100819 259798
rect 259494 259796 259500 259798
rect 259564 259796 259570 259860
rect 65885 259584 68938 259586
rect 65885 259528 65890 259584
rect 65946 259528 68938 259584
rect 65885 259526 68938 259528
rect 254577 259586 254643 259589
rect 270677 259588 270743 259589
rect 263726 259586 263732 259588
rect 254577 259584 263732 259586
rect 254577 259528 254582 259584
rect 254638 259528 263732 259584
rect 254577 259526 263732 259528
rect 65885 259523 65951 259526
rect 254577 259523 254643 259526
rect 263726 259524 263732 259526
rect 263796 259524 263802 259588
rect 270677 259584 270724 259588
rect 270788 259586 270794 259588
rect 270677 259528 270682 259584
rect 270677 259524 270724 259528
rect 270788 259526 270834 259586
rect 270788 259524 270794 259526
rect 270677 259523 270743 259524
rect 255405 259450 255471 259453
rect 253460 259448 255471 259450
rect 68185 258770 68251 258773
rect 68878 258770 68938 259284
rect 68185 258768 68938 258770
rect 68185 258712 68190 258768
rect 68246 258712 68938 258768
rect 68185 258710 68938 258712
rect 68185 258707 68251 258710
rect 98134 258501 98194 259012
rect 193397 258906 193463 258909
rect 193630 258906 193690 259420
rect 253460 259392 255410 259448
rect 255466 259392 255471 259448
rect 253460 259390 255471 259392
rect 255405 259387 255471 259390
rect 260741 259450 260807 259453
rect 262254 259450 262260 259452
rect 260741 259448 262260 259450
rect 260741 259392 260746 259448
rect 260802 259392 262260 259448
rect 260741 259390 262260 259392
rect 260741 259387 260807 259390
rect 262254 259388 262260 259390
rect 262324 259388 262330 259452
rect 193397 258904 193690 258906
rect 193397 258848 193402 258904
rect 193458 258848 193690 258904
rect 193397 258846 193690 258848
rect 253430 258906 253490 259012
rect 265065 258906 265131 258909
rect 270534 258906 270540 258908
rect 253430 258846 262874 258906
rect 193397 258843 193463 258846
rect 255589 258770 255655 258773
rect 262814 258770 262874 258846
rect 265065 258904 270540 258906
rect 265065 258848 265070 258904
rect 265126 258848 270540 258904
rect 265065 258846 270540 258848
rect 265065 258843 265131 258846
rect 270534 258844 270540 258846
rect 270604 258844 270610 258908
rect 580165 258906 580231 258909
rect 583520 258906 584960 258996
rect 580165 258904 584960 258906
rect 580165 258848 580170 258904
rect 580226 258848 584960 258904
rect 580165 258846 584960 258848
rect 580165 258843 580231 258846
rect 278129 258770 278195 258773
rect 255589 258768 258090 258770
rect 255589 258712 255594 258768
rect 255650 258712 258090 258768
rect 255589 258710 258090 258712
rect 262814 258768 278195 258770
rect 262814 258712 278134 258768
rect 278190 258712 278195 258768
rect 583520 258756 584960 258846
rect 262814 258710 278195 258712
rect 255589 258707 255655 258710
rect 255497 258634 255563 258637
rect 253460 258632 255563 258634
rect 253460 258576 255502 258632
rect 255558 258576 255563 258632
rect 253460 258574 255563 258576
rect 258030 258634 258090 258710
rect 278129 258707 278195 258710
rect 265065 258634 265131 258637
rect 258030 258632 265131 258634
rect 258030 258576 265070 258632
rect 265126 258576 265131 258632
rect 258030 258574 265131 258576
rect 255497 258571 255563 258574
rect 265065 258571 265131 258574
rect 66805 258498 66871 258501
rect 66805 258496 68908 258498
rect 66805 258440 66810 258496
rect 66866 258440 68908 258496
rect 66805 258438 68908 258440
rect 98085 258496 98194 258501
rect 254577 258498 254643 258501
rect 98085 258440 98090 258496
rect 98146 258440 98194 258496
rect 98085 258438 98194 258440
rect 253430 258496 254643 258498
rect 253430 258440 254582 258496
rect 254638 258440 254643 258496
rect 253430 258438 254643 258440
rect 66805 258435 66871 258438
rect 98085 258435 98151 258438
rect 191741 258362 191807 258365
rect 191741 258360 193660 258362
rect 191741 258304 191746 258360
rect 191802 258304 193660 258360
rect 191741 258302 193660 258304
rect 191741 258299 191807 258302
rect 59118 258164 59124 258228
rect 59188 258226 59194 258228
rect 59261 258226 59327 258229
rect 99281 258226 99347 258229
rect 101397 258226 101463 258229
rect 59188 258224 59327 258226
rect 59188 258168 59266 258224
rect 59322 258168 59327 258224
rect 59188 258166 59327 258168
rect 98716 258224 101463 258226
rect 98716 258168 99286 258224
rect 99342 258168 101402 258224
rect 101458 258168 101463 258224
rect 253430 258196 253490 258438
rect 254577 258435 254643 258438
rect 98716 258166 101463 258168
rect 59188 258164 59194 258166
rect 59261 258163 59327 258166
rect 99281 258163 99347 258166
rect 101397 258163 101463 258166
rect 66110 257892 66116 257956
rect 66180 257954 66186 257956
rect 66253 257954 66319 257957
rect 66180 257952 68938 257954
rect 66180 257896 66258 257952
rect 66314 257896 68938 257952
rect 66180 257894 68938 257896
rect 66180 257892 66186 257894
rect 66253 257891 66319 257894
rect 68878 257652 68938 257894
rect 253430 257682 253490 257788
rect 253430 257622 258090 257682
rect 100109 257410 100175 257413
rect 98716 257408 100175 257410
rect 98716 257352 100114 257408
rect 100170 257352 100175 257408
rect 98716 257350 100175 257352
rect 100109 257347 100175 257350
rect 191649 257410 191715 257413
rect 255405 257410 255471 257413
rect 191649 257408 193660 257410
rect 191649 257352 191654 257408
rect 191710 257352 193660 257408
rect 191649 257350 193660 257352
rect 253460 257408 255471 257410
rect 253460 257352 255410 257408
rect 255466 257352 255471 257408
rect 253460 257350 255471 257352
rect 191649 257347 191715 257350
rect 255405 257347 255471 257350
rect 255405 257002 255471 257005
rect 253460 257000 255471 257002
rect 253460 256944 255410 257000
rect 255466 256944 255471 257000
rect 253460 256942 255471 256944
rect 255405 256939 255471 256942
rect 66621 256868 66687 256869
rect 66621 256866 66668 256868
rect 66540 256864 66668 256866
rect 66732 256866 66738 256868
rect 258030 256866 258090 257622
rect 267958 256866 267964 256868
rect 66540 256808 66626 256864
rect 66540 256806 66668 256808
rect 66621 256804 66668 256806
rect 66732 256806 68908 256866
rect 258030 256806 267964 256866
rect 66732 256804 66738 256806
rect 267958 256804 267964 256806
rect 268028 256804 268034 256868
rect 66621 256803 66687 256804
rect 100845 256594 100911 256597
rect 255405 256594 255471 256597
rect 98716 256592 100911 256594
rect 98716 256536 100850 256592
rect 100906 256536 100911 256592
rect 98716 256534 100911 256536
rect 253460 256592 255471 256594
rect 253460 256536 255410 256592
rect 255466 256536 255471 256592
rect 253460 256534 255471 256536
rect 100845 256531 100911 256534
rect 255405 256531 255471 256534
rect 190821 256458 190887 256461
rect 190821 256456 193660 256458
rect 190821 256400 190826 256456
rect 190882 256400 193660 256456
rect 190821 256398 193660 256400
rect 190821 256395 190887 256398
rect 255589 256186 255655 256189
rect 253460 256184 255655 256186
rect 253460 256128 255594 256184
rect 255650 256128 255655 256184
rect 253460 256126 255655 256128
rect 255589 256123 255655 256126
rect 44081 255914 44147 255917
rect 61878 255914 61884 255916
rect 44081 255912 61884 255914
rect 44081 255856 44086 255912
rect 44142 255856 61884 255912
rect 44081 255854 61884 255856
rect 44081 255851 44147 255854
rect 61878 255852 61884 255854
rect 61948 255914 61954 255916
rect 68878 255914 68938 256020
rect 61948 255854 68938 255914
rect 61948 255852 61954 255854
rect 101397 255778 101463 255781
rect 98716 255776 101463 255778
rect 98716 255720 101402 255776
rect 101458 255720 101463 255776
rect 98716 255718 101463 255720
rect 101397 255715 101463 255718
rect 253430 255642 253490 255748
rect 273529 255642 273595 255645
rect 283097 255642 283163 255645
rect 253430 255640 283163 255642
rect 253430 255584 273534 255640
rect 273590 255584 283102 255640
rect 283158 255584 283163 255640
rect 253430 255582 283163 255584
rect 273529 255579 273595 255582
rect 283097 255579 283163 255582
rect 191005 255506 191071 255509
rect 191005 255504 193660 255506
rect 191005 255448 191010 255504
rect 191066 255448 193660 255504
rect 191005 255446 193660 255448
rect 191005 255443 191071 255446
rect 255497 255370 255563 255373
rect 253460 255368 255563 255370
rect 253460 255312 255502 255368
rect 255558 255312 255563 255368
rect 253460 255310 255563 255312
rect 255497 255307 255563 255310
rect 52361 255234 52427 255237
rect 266905 255234 266971 255237
rect 269246 255234 269252 255236
rect 52361 255232 68908 255234
rect 52361 255176 52366 255232
rect 52422 255176 68908 255232
rect 52361 255174 68908 255176
rect 266905 255232 269252 255234
rect 266905 255176 266910 255232
rect 266966 255176 269252 255232
rect 266905 255174 269252 255176
rect 52361 255171 52427 255174
rect 266905 255171 266971 255174
rect 269246 255172 269252 255174
rect 269316 255172 269322 255236
rect 100845 254962 100911 254965
rect 98164 254960 100911 254962
rect 98164 254932 100850 254960
rect 98134 254904 100850 254932
rect 100906 254904 100911 254960
rect 98134 254902 100911 254904
rect 66805 254418 66871 254421
rect 98134 254420 98194 254902
rect 100845 254899 100911 254902
rect 253430 254826 253490 254932
rect 255221 254826 255287 254829
rect 253430 254824 255287 254826
rect 253430 254768 255226 254824
rect 255282 254768 255287 254824
rect 253430 254766 255287 254768
rect 255221 254763 255287 254766
rect 191649 254554 191715 254557
rect 255405 254554 255471 254557
rect 191649 254552 193660 254554
rect 191649 254496 191654 254552
rect 191710 254496 193660 254552
rect 191649 254494 193660 254496
rect 253460 254552 255471 254554
rect 253460 254496 255410 254552
rect 255466 254496 255471 254552
rect 253460 254494 255471 254496
rect 191649 254491 191715 254494
rect 255405 254491 255471 254494
rect 255589 254554 255655 254557
rect 278957 254554 279023 254557
rect 285622 254554 285628 254556
rect 255589 254552 285628 254554
rect 255589 254496 255594 254552
rect 255650 254496 278962 254552
rect 279018 254496 285628 254552
rect 255589 254494 285628 254496
rect 255589 254491 255655 254494
rect 278957 254491 279023 254494
rect 285622 254492 285628 254494
rect 285692 254492 285698 254556
rect 66805 254416 68908 254418
rect 66805 254360 66810 254416
rect 66866 254360 68908 254416
rect 66805 254358 68908 254360
rect 66805 254355 66871 254358
rect 98126 254356 98132 254420
rect 98196 254356 98202 254420
rect 255221 254418 255287 254421
rect 270677 254418 270743 254421
rect 255221 254416 270743 254418
rect 255221 254360 255226 254416
rect 255282 254360 270682 254416
rect 270738 254360 270743 254416
rect 255221 254358 270743 254360
rect 255221 254355 255287 254358
rect 270677 254355 270743 254358
rect -960 254146 480 254236
rect 3141 254146 3207 254149
rect 100845 254146 100911 254149
rect 255497 254146 255563 254149
rect -960 254144 3207 254146
rect -960 254088 3146 254144
rect 3202 254088 3207 254144
rect -960 254086 3207 254088
rect 98716 254144 100911 254146
rect 98716 254088 100850 254144
rect 100906 254088 100911 254144
rect 98716 254086 100911 254088
rect 253460 254144 255563 254146
rect 253460 254088 255502 254144
rect 255558 254088 255563 254144
rect 253460 254086 255563 254088
rect -960 253996 480 254086
rect 3141 254083 3207 254086
rect 100845 254083 100911 254086
rect 255497 254083 255563 254086
rect 46841 254010 46907 254013
rect 52361 254010 52427 254013
rect 46841 254008 52427 254010
rect 46841 253952 46846 254008
rect 46902 253952 52366 254008
rect 52422 253952 52427 254008
rect 46841 253950 52427 253952
rect 46841 253947 46907 253950
rect 52361 253947 52427 253950
rect 253933 253738 253999 253741
rect 258390 253738 258396 253740
rect 253460 253736 258396 253738
rect 253460 253680 253938 253736
rect 253994 253680 258396 253736
rect 253460 253678 258396 253680
rect 253933 253675 253999 253678
rect 258390 253676 258396 253678
rect 258460 253676 258466 253740
rect 66989 253602 67055 253605
rect 191557 253602 191623 253605
rect 66989 253600 68908 253602
rect 66989 253544 66994 253600
rect 67050 253544 68908 253600
rect 66989 253542 68908 253544
rect 191557 253600 193660 253602
rect 191557 253544 191562 253600
rect 191618 253544 193660 253600
rect 191557 253542 193660 253544
rect 66989 253539 67055 253542
rect 191557 253539 191623 253542
rect 100845 253330 100911 253333
rect 98716 253328 100911 253330
rect 98716 253272 100850 253328
rect 100906 253272 100911 253328
rect 98716 253270 100911 253272
rect 100845 253267 100911 253270
rect 252878 253197 252938 253300
rect 252829 253192 252938 253197
rect 252829 253136 252834 253192
rect 252890 253136 252938 253192
rect 252829 253134 252938 253136
rect 252829 253131 252895 253134
rect 255405 252922 255471 252925
rect 253460 252920 255471 252922
rect 253460 252864 255410 252920
rect 255466 252864 255471 252920
rect 253460 252862 255471 252864
rect 255405 252859 255471 252862
rect 62113 252786 62179 252789
rect 63401 252786 63467 252789
rect 62113 252784 68908 252786
rect 62113 252728 62118 252784
rect 62174 252728 63406 252784
rect 63462 252728 68908 252784
rect 62113 252726 68908 252728
rect 62113 252723 62179 252726
rect 63401 252723 63467 252726
rect 191649 252650 191715 252653
rect 191649 252648 193660 252650
rect 191649 252592 191654 252648
rect 191710 252592 193660 252648
rect 191649 252590 193660 252592
rect 191649 252587 191715 252590
rect 269062 252588 269068 252652
rect 269132 252650 269138 252652
rect 269389 252650 269455 252653
rect 269132 252648 269455 252650
rect 269132 252592 269394 252648
rect 269450 252592 269455 252648
rect 269132 252590 269455 252592
rect 269132 252588 269138 252590
rect 269389 252587 269455 252590
rect 100702 252514 100708 252516
rect 98716 252454 100708 252514
rect 100702 252452 100708 252454
rect 100772 252514 100778 252516
rect 101673 252514 101739 252517
rect 255405 252514 255471 252517
rect 100772 252512 101739 252514
rect 100772 252456 101678 252512
rect 101734 252456 101739 252512
rect 100772 252454 101739 252456
rect 253460 252512 255471 252514
rect 253460 252456 255410 252512
rect 255466 252456 255471 252512
rect 253460 252454 255471 252456
rect 100772 252452 100778 252454
rect 101673 252451 101739 252454
rect 255405 252451 255471 252454
rect 255497 252106 255563 252109
rect 253460 252104 255563 252106
rect 253460 252048 255502 252104
rect 255558 252048 255563 252104
rect 253460 252046 255563 252048
rect 255497 252043 255563 252046
rect 66805 251970 66871 251973
rect 66805 251968 68908 251970
rect 66805 251912 66810 251968
rect 66866 251912 68908 251968
rect 66805 251910 68908 251912
rect 66805 251907 66871 251910
rect 182909 251834 182975 251837
rect 193254 251834 193260 251836
rect 182909 251832 193260 251834
rect 182909 251776 182914 251832
rect 182970 251776 193260 251832
rect 182909 251774 193260 251776
rect 182909 251771 182975 251774
rect 193254 251772 193260 251774
rect 193324 251772 193330 251836
rect 98686 251290 98746 251668
rect 98686 251230 100034 251290
rect 99974 251157 100034 251230
rect 177246 251228 177252 251292
rect 177316 251290 177322 251292
rect 193630 251290 193690 251668
rect 258533 251562 258599 251565
rect 253460 251560 258599 251562
rect 253460 251504 258538 251560
rect 258594 251504 258599 251560
rect 253460 251502 258599 251504
rect 258533 251499 258599 251502
rect 177316 251230 193690 251290
rect 177316 251228 177322 251230
rect 66437 251156 66503 251157
rect 66437 251154 66484 251156
rect 66356 251152 66484 251154
rect 66548 251154 66554 251156
rect 99974 251154 100083 251157
rect 137461 251154 137527 251157
rect 255497 251154 255563 251157
rect 66356 251096 66442 251152
rect 66356 251094 66484 251096
rect 66437 251092 66484 251094
rect 66548 251094 68908 251154
rect 99974 251152 137527 251154
rect 99974 251096 100022 251152
rect 100078 251096 137466 251152
rect 137522 251096 137527 251152
rect 99974 251094 137527 251096
rect 253460 251152 255563 251154
rect 253460 251096 255502 251152
rect 255558 251096 255563 251152
rect 253460 251094 255563 251096
rect 66548 251092 66554 251094
rect 66437 251091 66503 251092
rect 100017 251091 100083 251094
rect 137461 251091 137527 251094
rect 255497 251091 255563 251094
rect 271965 251154 272031 251157
rect 272558 251154 272564 251156
rect 271965 251152 272564 251154
rect 271965 251096 271970 251152
rect 272026 251096 272564 251152
rect 271965 251094 272564 251096
rect 271965 251091 272031 251094
rect 272558 251092 272564 251094
rect 272628 251092 272634 251156
rect 100845 250882 100911 250885
rect 98716 250880 100911 250882
rect 98716 250824 100850 250880
rect 100906 250824 100911 250880
rect 98716 250822 100911 250824
rect 100845 250819 100911 250822
rect 190637 250746 190703 250749
rect 272149 250746 272215 250749
rect 190637 250744 193660 250746
rect 190637 250688 190642 250744
rect 190698 250688 193660 250744
rect 190637 250686 193660 250688
rect 253460 250744 277410 250746
rect 253460 250688 272154 250744
rect 272210 250688 277410 250744
rect 253460 250686 277410 250688
rect 190637 250683 190703 250686
rect 272149 250683 272215 250686
rect 271965 250610 272031 250613
rect 253430 250608 272031 250610
rect 253430 250552 271970 250608
rect 272026 250552 272031 250608
rect 253430 250550 272031 250552
rect 66805 250338 66871 250341
rect 66805 250336 68908 250338
rect 66805 250280 66810 250336
rect 66866 250280 68908 250336
rect 253430 250308 253490 250550
rect 271965 250547 272031 250550
rect 277350 250474 277410 250686
rect 582557 250474 582623 250477
rect 277350 250472 582623 250474
rect 277350 250416 582562 250472
rect 582618 250416 582623 250472
rect 277350 250414 582623 250416
rect 582557 250411 582623 250414
rect 66805 250278 68908 250280
rect 66805 250275 66871 250278
rect 101949 250066 102015 250069
rect 98716 250064 102015 250066
rect 98716 250008 101954 250064
rect 102010 250008 102015 250064
rect 98716 250006 102015 250008
rect 101949 250003 102015 250006
rect 255865 249930 255931 249933
rect 253460 249928 255931 249930
rect 253460 249872 255870 249928
rect 255926 249872 255931 249928
rect 253460 249870 255931 249872
rect 255865 249867 255931 249870
rect 262070 249732 262076 249796
rect 262140 249794 262146 249796
rect 262438 249794 262444 249796
rect 262140 249734 262444 249794
rect 262140 249732 262146 249734
rect 262438 249732 262444 249734
rect 262508 249732 262514 249796
rect 190821 249658 190887 249661
rect 190821 249656 193660 249658
rect 190821 249600 190826 249656
rect 190882 249600 193660 249656
rect 190821 249598 193660 249600
rect 190821 249595 190887 249598
rect 66621 249522 66687 249525
rect 253933 249522 253999 249525
rect 254945 249522 255011 249525
rect 66621 249520 68908 249522
rect 66621 249464 66626 249520
rect 66682 249464 68908 249520
rect 66621 249462 68908 249464
rect 253460 249520 255011 249522
rect 253460 249464 253938 249520
rect 253994 249464 254950 249520
rect 255006 249464 255011 249520
rect 253460 249462 255011 249464
rect 66621 249459 66687 249462
rect 253933 249459 253999 249462
rect 254945 249459 255011 249462
rect 100845 249250 100911 249253
rect 98716 249248 100911 249250
rect 98716 249192 100850 249248
rect 100906 249192 100911 249248
rect 98716 249190 100911 249192
rect 100845 249187 100911 249190
rect 255405 249114 255471 249117
rect 253460 249112 255471 249114
rect 253460 249056 255410 249112
rect 255466 249056 255471 249112
rect 253460 249054 255471 249056
rect 255405 249051 255471 249054
rect 66161 248706 66227 248709
rect 254577 248706 254643 248709
rect 66161 248704 68908 248706
rect 66161 248648 66166 248704
rect 66222 248648 68908 248704
rect 253460 248704 254643 248706
rect 66161 248646 68908 248648
rect 66161 248643 66227 248646
rect 99189 248434 99255 248437
rect 98348 248432 99255 248434
rect 98348 248430 99194 248432
rect 98318 248376 99194 248430
rect 99250 248376 99255 248432
rect 98318 248374 99255 248376
rect 98318 248301 98378 248374
rect 99189 248371 99255 248374
rect 188521 248434 188587 248437
rect 193630 248434 193690 248676
rect 253460 248648 254582 248704
rect 254638 248648 254643 248704
rect 253460 248646 254643 248648
rect 254577 248643 254643 248646
rect 188521 248432 193690 248434
rect 188521 248376 188526 248432
rect 188582 248376 193690 248432
rect 188521 248374 193690 248376
rect 188521 248371 188587 248374
rect 267774 248372 267780 248436
rect 267844 248434 267850 248436
rect 269021 248434 269087 248437
rect 267844 248432 269087 248434
rect 267844 248376 269026 248432
rect 269082 248376 269087 248432
rect 267844 248374 269087 248376
rect 267844 248372 267850 248374
rect 269021 248371 269087 248374
rect 98269 248296 98378 248301
rect 98269 248240 98274 248296
rect 98330 248240 98378 248296
rect 98269 248238 98378 248240
rect 98269 248235 98335 248238
rect 252878 248164 252938 248268
rect 252870 248100 252876 248164
rect 252940 248100 252946 248164
rect 262673 247890 262739 247893
rect 262806 247890 262812 247892
rect 262673 247888 262812 247890
rect 68878 247346 68938 247860
rect 191649 247754 191715 247757
rect 253430 247754 253490 247860
rect 262673 247832 262678 247888
rect 262734 247832 262812 247888
rect 262673 247830 262812 247832
rect 262673 247827 262739 247830
rect 262806 247828 262812 247830
rect 262876 247890 262882 247892
rect 266302 247890 266308 247892
rect 262876 247830 266308 247890
rect 262876 247828 262882 247830
rect 266302 247828 266308 247830
rect 266372 247828 266378 247892
rect 283005 247754 283071 247757
rect 191649 247752 193660 247754
rect 191649 247696 191654 247752
rect 191710 247696 193660 247752
rect 191649 247694 193660 247696
rect 253430 247752 283071 247754
rect 253430 247696 283010 247752
rect 283066 247696 283071 247752
rect 253430 247694 283071 247696
rect 191649 247691 191715 247694
rect 283005 247691 283071 247694
rect 100201 247618 100267 247621
rect 98716 247616 100267 247618
rect 98716 247560 100206 247616
rect 100262 247560 100267 247616
rect 98716 247558 100267 247560
rect 100201 247555 100267 247558
rect 254209 247482 254275 247485
rect 253460 247480 254275 247482
rect 253460 247424 254214 247480
rect 254270 247424 254275 247480
rect 253460 247422 254275 247424
rect 254209 247419 254275 247422
rect 64830 247286 68938 247346
rect 57830 247148 57836 247212
rect 57900 247210 57906 247212
rect 64830 247210 64890 247286
rect 57900 247150 64890 247210
rect 57900 247148 57906 247150
rect 67449 247074 67515 247077
rect 255497 247074 255563 247077
rect 67449 247072 68908 247074
rect 67449 247016 67454 247072
rect 67510 247016 68908 247072
rect 67449 247014 68908 247016
rect 253460 247072 255563 247074
rect 253460 247016 255502 247072
rect 255558 247016 255563 247072
rect 253460 247014 255563 247016
rect 67449 247011 67515 247014
rect 255497 247011 255563 247014
rect 100845 246802 100911 246805
rect 98716 246800 100911 246802
rect 98716 246744 100850 246800
rect 100906 246744 100911 246800
rect 98716 246742 100911 246744
rect 100845 246739 100911 246742
rect 67357 246258 67423 246261
rect 67357 246256 68908 246258
rect 67357 246200 67362 246256
rect 67418 246200 68908 246256
rect 67357 246198 68908 246200
rect 67357 246195 67423 246198
rect 160686 246196 160692 246260
rect 160756 246258 160762 246260
rect 181529 246258 181595 246261
rect 160756 246256 181595 246258
rect 160756 246200 181534 246256
rect 181590 246200 181595 246256
rect 160756 246198 181595 246200
rect 160756 246196 160762 246198
rect 181529 246195 181595 246198
rect 192017 246258 192083 246261
rect 193630 246258 193690 246772
rect 255405 246666 255471 246669
rect 253460 246664 255471 246666
rect 253460 246608 255410 246664
rect 255466 246608 255471 246664
rect 253460 246606 255471 246608
rect 255405 246603 255471 246606
rect 255681 246258 255747 246261
rect 192017 246256 193690 246258
rect 192017 246200 192022 246256
rect 192078 246200 193690 246256
rect 192017 246198 193690 246200
rect 253460 246256 255747 246258
rect 253460 246200 255686 246256
rect 255742 246200 255747 246256
rect 253460 246198 255747 246200
rect 192017 246195 192083 246198
rect 255681 246195 255747 246198
rect 100845 245986 100911 245989
rect 98716 245984 100911 245986
rect 98716 245928 100850 245984
rect 100906 245928 100911 245984
rect 98716 245926 100911 245928
rect 100845 245923 100911 245926
rect 189717 245850 189783 245853
rect 255405 245850 255471 245853
rect 189717 245848 193660 245850
rect 189717 245792 189722 245848
rect 189778 245792 193660 245848
rect 189717 245790 193660 245792
rect 253460 245848 255471 245850
rect 253460 245792 255410 245848
rect 255466 245792 255471 245848
rect 253460 245790 255471 245792
rect 189717 245787 189783 245790
rect 255405 245787 255471 245790
rect 184238 245652 184244 245716
rect 184308 245714 184314 245716
rect 192017 245714 192083 245717
rect 184308 245712 192083 245714
rect 184308 245656 192022 245712
rect 192078 245656 192083 245712
rect 184308 245654 192083 245656
rect 184308 245652 184314 245654
rect 192017 245651 192083 245654
rect 582373 245578 582439 245581
rect 583520 245578 584960 245668
rect 582373 245576 584960 245578
rect 582373 245520 582378 245576
rect 582434 245520 584960 245576
rect 582373 245518 584960 245520
rect 582373 245515 582439 245518
rect 255405 245442 255471 245445
rect 253460 245440 255471 245442
rect 68878 244898 68938 245412
rect 253460 245384 255410 245440
rect 255466 245384 255471 245440
rect 583520 245428 584960 245518
rect 253460 245382 255471 245384
rect 255405 245379 255471 245382
rect 100845 245170 100911 245173
rect 98716 245168 100911 245170
rect 98716 245112 100850 245168
rect 100906 245112 100911 245168
rect 98716 245110 100911 245112
rect 100845 245107 100911 245110
rect 255589 245034 255655 245037
rect 253460 245032 255655 245034
rect 253460 244976 255594 245032
rect 255650 244976 255655 245032
rect 253460 244974 255655 244976
rect 255589 244971 255655 244974
rect 64830 244838 68938 244898
rect 191649 244898 191715 244901
rect 191649 244896 193660 244898
rect 191649 244840 191654 244896
rect 191710 244840 193660 244896
rect 191649 244838 193660 244840
rect 64638 244428 64644 244492
rect 64708 244490 64714 244492
rect 64830 244490 64890 244838
rect 191649 244835 191715 244838
rect 66805 244626 66871 244629
rect 255497 244626 255563 244629
rect 66805 244624 68908 244626
rect 66805 244568 66810 244624
rect 66866 244568 68908 244624
rect 66805 244566 68908 244568
rect 253460 244624 255563 244626
rect 253460 244568 255502 244624
rect 255558 244568 255563 244624
rect 253460 244566 255563 244568
rect 66805 244563 66871 244566
rect 255497 244563 255563 244566
rect 64708 244430 64890 244490
rect 64708 244428 64714 244430
rect 100937 244354 101003 244357
rect 98716 244352 101003 244354
rect 98716 244296 100942 244352
rect 100998 244296 101003 244352
rect 98716 244294 101003 244296
rect 100937 244291 101003 244294
rect 255405 244218 255471 244221
rect 253460 244216 255471 244218
rect 253460 244160 255410 244216
rect 255466 244160 255471 244216
rect 253460 244158 255471 244160
rect 255405 244155 255471 244158
rect 191649 243946 191715 243949
rect 191649 243944 193660 243946
rect 191649 243888 191654 243944
rect 191710 243888 193660 243944
rect 191649 243886 193660 243888
rect 191649 243883 191715 243886
rect 66621 243810 66687 243813
rect 255497 243810 255563 243813
rect 66621 243808 68908 243810
rect 66621 243752 66626 243808
rect 66682 243752 68908 243808
rect 66621 243750 68908 243752
rect 253460 243808 255563 243810
rect 253460 243752 255502 243808
rect 255558 243752 255563 243808
rect 253460 243750 255563 243752
rect 66621 243747 66687 243750
rect 255497 243747 255563 243750
rect 100845 243538 100911 243541
rect 98716 243536 100911 243538
rect 98716 243480 100850 243536
rect 100906 243480 100911 243536
rect 98716 243478 100911 243480
rect 100845 243475 100911 243478
rect 253430 243266 253490 243372
rect 253430 243206 258090 243266
rect 66805 242994 66871 242997
rect 189993 242994 190059 242997
rect 258030 242994 258090 243206
rect 66805 242992 68908 242994
rect 66805 242936 66810 242992
rect 66866 242936 68908 242992
rect 66805 242934 68908 242936
rect 189993 242992 193660 242994
rect 189993 242936 189998 242992
rect 190054 242936 193660 242992
rect 189993 242934 193660 242936
rect 66805 242931 66871 242934
rect 189993 242931 190059 242934
rect 252878 242861 252938 242964
rect 258030 242934 265082 242994
rect 193254 242796 193260 242860
rect 193324 242858 193330 242860
rect 193673 242858 193739 242861
rect 193324 242856 193739 242858
rect 193324 242800 193678 242856
rect 193734 242800 193739 242856
rect 193324 242798 193739 242800
rect 193324 242796 193330 242798
rect 193673 242795 193739 242798
rect 252829 242856 252938 242861
rect 252829 242800 252834 242856
rect 252890 242800 252938 242856
rect 252829 242798 252938 242800
rect 265022 242858 265082 242934
rect 265617 242858 265683 242861
rect 273294 242858 273300 242860
rect 265022 242856 273300 242858
rect 265022 242800 265622 242856
rect 265678 242800 273300 242856
rect 265022 242798 273300 242800
rect 252829 242795 252895 242798
rect 265617 242795 265683 242798
rect 273294 242796 273300 242798
rect 273364 242796 273370 242860
rect 284385 242858 284451 242861
rect 284569 242858 284635 242861
rect 284385 242856 284635 242858
rect 284385 242800 284390 242856
rect 284446 242800 284574 242856
rect 284630 242800 284635 242856
rect 284385 242798 284635 242800
rect 284385 242795 284451 242798
rect 284569 242795 284635 242798
rect 102317 242722 102383 242725
rect 98716 242720 102383 242722
rect 98716 242664 102322 242720
rect 102378 242664 102383 242720
rect 98716 242662 102383 242664
rect 102317 242659 102383 242662
rect 252878 242453 252938 242556
rect 252878 242448 252987 242453
rect 252878 242392 252926 242448
rect 252982 242392 252987 242448
rect 252878 242390 252987 242392
rect 252921 242387 252987 242390
rect 255589 242314 255655 242317
rect 259678 242314 259684 242316
rect 255589 242312 259684 242314
rect 255589 242256 255594 242312
rect 255650 242256 259684 242312
rect 255589 242254 259684 242256
rect 255589 242251 255655 242254
rect 259678 242252 259684 242254
rect 259748 242314 259754 242316
rect 277158 242314 277164 242316
rect 259748 242254 277164 242314
rect 259748 242252 259754 242254
rect 277158 242252 277164 242254
rect 277228 242252 277234 242316
rect 57697 242178 57763 242181
rect 66294 242178 66300 242180
rect 57697 242176 66300 242178
rect 57697 242120 57702 242176
rect 57758 242120 66300 242176
rect 57697 242118 66300 242120
rect 57697 242115 57763 242118
rect 66294 242116 66300 242118
rect 66364 242178 66370 242180
rect 256049 242178 256115 242181
rect 284385 242178 284451 242181
rect 66364 242118 68908 242178
rect 253460 242176 256115 242178
rect 253460 242120 256054 242176
rect 256110 242120 256115 242176
rect 253460 242118 256115 242120
rect 66364 242116 66370 242118
rect 256049 242115 256115 242118
rect 258030 242176 284451 242178
rect 258030 242120 284390 242176
rect 284446 242120 284451 242176
rect 258030 242118 284451 242120
rect 258030 242042 258090 242118
rect 284385 242115 284451 242118
rect 104249 241906 104315 241909
rect 98716 241904 104315 241906
rect 98716 241848 104254 241904
rect 104310 241848 104315 241904
rect 98716 241846 104315 241848
rect 104249 241843 104315 241846
rect 68686 241708 68692 241772
rect 68756 241770 68762 241772
rect 69473 241770 69539 241773
rect 72693 241772 72759 241773
rect 73245 241772 73311 241773
rect 72693 241770 72740 241772
rect 68756 241768 69539 241770
rect 68756 241712 69478 241768
rect 69534 241712 69539 241768
rect 68756 241710 69539 241712
rect 72648 241768 72740 241770
rect 72648 241712 72698 241768
rect 72648 241710 72740 241712
rect 68756 241708 68762 241710
rect 69473 241707 69539 241710
rect 72693 241708 72740 241710
rect 72804 241708 72810 241772
rect 73245 241770 73292 241772
rect 73164 241768 73292 241770
rect 73356 241770 73362 241772
rect 73797 241770 73863 241773
rect 73356 241768 73863 241770
rect 73164 241712 73250 241768
rect 73356 241712 73802 241768
rect 73858 241712 73863 241768
rect 73164 241710 73292 241712
rect 73245 241708 73292 241710
rect 73356 241710 73863 241712
rect 73356 241708 73362 241710
rect 72693 241707 72759 241708
rect 73245 241707 73311 241708
rect 73797 241707 73863 241710
rect 83733 241770 83799 241773
rect 84694 241770 84700 241772
rect 83733 241768 84700 241770
rect 83733 241712 83738 241768
rect 83794 241712 84700 241768
rect 83733 241710 84700 241712
rect 83733 241707 83799 241710
rect 84694 241708 84700 241710
rect 84764 241708 84770 241772
rect 86585 241770 86651 241773
rect 87137 241772 87203 241773
rect 86718 241770 86724 241772
rect 86585 241768 86724 241770
rect 86585 241712 86590 241768
rect 86646 241712 86724 241768
rect 86585 241710 86724 241712
rect 86585 241707 86651 241710
rect 86718 241708 86724 241710
rect 86788 241708 86794 241772
rect 87086 241708 87092 241772
rect 87156 241770 87203 241772
rect 90357 241770 90423 241773
rect 91553 241772 91619 241773
rect 90950 241770 90956 241772
rect 87156 241768 87248 241770
rect 87198 241712 87248 241768
rect 87156 241710 87248 241712
rect 90357 241768 90956 241770
rect 90357 241712 90362 241768
rect 90418 241712 90956 241768
rect 90357 241710 90956 241712
rect 87156 241708 87203 241710
rect 87137 241707 87203 241708
rect 90357 241707 90423 241710
rect 90950 241708 90956 241710
rect 91020 241708 91026 241772
rect 91502 241708 91508 241772
rect 91572 241770 91619 241772
rect 93761 241770 93827 241773
rect 93894 241770 93900 241772
rect 91572 241768 91664 241770
rect 91614 241712 91664 241768
rect 91572 241710 91664 241712
rect 93761 241768 93900 241770
rect 93761 241712 93766 241768
rect 93822 241712 93900 241768
rect 93761 241710 93900 241712
rect 91572 241708 91619 241710
rect 91553 241707 91619 241708
rect 93761 241707 93827 241710
rect 93894 241708 93900 241710
rect 93964 241708 93970 241772
rect 85941 241634 86007 241637
rect 87454 241634 87460 241636
rect 85941 241632 87460 241634
rect 85941 241576 85946 241632
rect 86002 241576 87460 241632
rect 85941 241574 87460 241576
rect 85941 241571 86007 241574
rect 86910 241501 86970 241574
rect 87454 241572 87460 241574
rect 87524 241572 87530 241636
rect 97717 241634 97783 241637
rect 102225 241634 102291 241637
rect 97717 241632 102291 241634
rect 97717 241576 97722 241632
rect 97778 241576 102230 241632
rect 102286 241576 102291 241632
rect 97717 241574 102291 241576
rect 97717 241571 97783 241574
rect 102225 241571 102291 241574
rect 188286 241572 188292 241636
rect 188356 241634 188362 241636
rect 193630 241634 193690 242012
rect 253430 241982 258090 242042
rect 253430 241740 253490 241982
rect 188356 241574 193690 241634
rect 188356 241572 188362 241574
rect 69657 241498 69723 241501
rect 70301 241500 70367 241501
rect 86585 241500 86651 241501
rect 70301 241498 70348 241500
rect 69657 241496 70348 241498
rect 69657 241440 69662 241496
rect 69718 241440 70306 241496
rect 69657 241438 70348 241440
rect 69657 241435 69723 241438
rect 70301 241436 70348 241438
rect 70412 241436 70418 241500
rect 86534 241436 86540 241500
rect 86604 241498 86651 241500
rect 86604 241496 86696 241498
rect 86646 241440 86696 241496
rect 86604 241438 86696 241440
rect 86861 241496 86970 241501
rect 86861 241440 86866 241496
rect 86922 241440 86970 241496
rect 86861 241438 86970 241440
rect 88057 241498 88123 241501
rect 187049 241498 187115 241501
rect 187601 241498 187667 241501
rect 201585 241500 201651 241501
rect 208393 241500 208459 241501
rect 215201 241500 215267 241501
rect 88057 241496 180810 241498
rect 88057 241440 88062 241496
rect 88118 241440 180810 241496
rect 88057 241438 180810 241440
rect 86604 241436 86651 241438
rect 70301 241435 70367 241436
rect 86585 241435 86651 241436
rect 86861 241435 86927 241438
rect 88057 241435 88123 241438
rect 68870 241300 68876 241364
rect 68940 241362 68946 241364
rect 70807 241362 70873 241365
rect 68940 241360 70873 241362
rect 68940 241304 70812 241360
rect 70868 241304 70873 241360
rect 68940 241302 70873 241304
rect 68940 241300 68946 241302
rect 70807 241299 70873 241302
rect 71313 241362 71379 241365
rect 106917 241362 106983 241365
rect 71313 241360 106983 241362
rect 71313 241304 71318 241360
rect 71374 241304 106922 241360
rect 106978 241304 106983 241360
rect 71313 241302 106983 241304
rect 71313 241299 71379 241302
rect 106917 241299 106983 241302
rect 84101 241226 84167 241229
rect 88057 241226 88123 241229
rect 84101 241224 88123 241226
rect -960 241090 480 241180
rect 84101 241168 84106 241224
rect 84162 241168 88062 241224
rect 88118 241168 88123 241224
rect 84101 241166 88123 241168
rect 84101 241163 84167 241166
rect 88057 241163 88123 241166
rect 89621 241226 89687 241229
rect 93761 241226 93827 241229
rect 89621 241224 93827 241226
rect 89621 241168 89626 241224
rect 89682 241168 93766 241224
rect 93822 241168 93827 241224
rect 89621 241166 93827 241168
rect 89621 241163 89687 241166
rect 93761 241163 93827 241166
rect 3509 241090 3575 241093
rect -960 241088 3575 241090
rect -960 241032 3514 241088
rect 3570 241032 3575 241088
rect -960 241030 3575 241032
rect 180750 241090 180810 241438
rect 187049 241496 187667 241498
rect 187049 241440 187054 241496
rect 187110 241440 187606 241496
rect 187662 241440 187667 241496
rect 187049 241438 187667 241440
rect 187049 241435 187115 241438
rect 187601 241435 187667 241438
rect 201534 241436 201540 241500
rect 201604 241498 201651 241500
rect 201604 241496 201696 241498
rect 201646 241440 201696 241496
rect 201604 241438 201696 241440
rect 201604 241436 201651 241438
rect 208342 241436 208348 241500
rect 208412 241498 208459 241500
rect 208412 241496 208504 241498
rect 208454 241440 208504 241496
rect 208412 241438 208504 241440
rect 208412 241436 208459 241438
rect 215150 241436 215156 241500
rect 215220 241498 215267 241500
rect 218605 241500 218671 241501
rect 218605 241498 218652 241500
rect 215220 241496 215312 241498
rect 215262 241440 215312 241496
rect 215220 241438 215312 241440
rect 218560 241496 218652 241498
rect 218560 241440 218610 241496
rect 218560 241438 218652 241440
rect 215220 241436 215267 241438
rect 201585 241435 201651 241436
rect 208393 241435 208459 241436
rect 215201 241435 215267 241436
rect 218605 241436 218652 241438
rect 218716 241436 218722 241500
rect 220905 241498 220971 241501
rect 221222 241498 221228 241500
rect 220905 241496 221228 241498
rect 220905 241440 220910 241496
rect 220966 241440 221228 241496
rect 220905 241438 221228 241440
rect 218605 241435 218671 241436
rect 220905 241435 220971 241438
rect 221222 241436 221228 241438
rect 221292 241498 221298 241500
rect 221549 241498 221615 241501
rect 221292 241496 221615 241498
rect 221292 241440 221554 241496
rect 221610 241440 221615 241496
rect 221292 241438 221615 241440
rect 221292 241436 221298 241438
rect 221549 241435 221615 241438
rect 225505 241498 225571 241501
rect 226190 241498 226196 241500
rect 225505 241496 226196 241498
rect 225505 241440 225510 241496
rect 225566 241440 226196 241496
rect 225505 241438 226196 241440
rect 225505 241435 225571 241438
rect 226190 241436 226196 241438
rect 226260 241436 226266 241500
rect 235441 241498 235507 241501
rect 236494 241498 236500 241500
rect 235441 241496 236500 241498
rect 235441 241440 235446 241496
rect 235502 241440 236500 241496
rect 235441 241438 236500 241440
rect 235441 241435 235507 241438
rect 236494 241436 236500 241438
rect 236564 241436 236570 241500
rect 238661 241498 238727 241501
rect 238886 241498 238892 241500
rect 238661 241496 238892 241498
rect 238661 241440 238666 241496
rect 238722 241440 238892 241496
rect 238661 241438 238892 241440
rect 238661 241435 238727 241438
rect 238886 241436 238892 241438
rect 238956 241436 238962 241500
rect 242249 241498 242315 241501
rect 242750 241498 242756 241500
rect 242249 241496 242756 241498
rect 242249 241440 242254 241496
rect 242310 241440 242756 241496
rect 242249 241438 242756 241440
rect 242249 241435 242315 241438
rect 242750 241436 242756 241438
rect 242820 241436 242826 241500
rect 245510 241436 245516 241500
rect 245580 241498 245586 241500
rect 245653 241498 245719 241501
rect 245580 241496 245719 241498
rect 245580 241440 245658 241496
rect 245714 241440 245719 241496
rect 245580 241438 245719 241440
rect 245580 241436 245586 241438
rect 245653 241435 245719 241438
rect 188981 241090 189047 241093
rect 238753 241090 238819 241093
rect 258257 241090 258323 241093
rect 180750 241088 190470 241090
rect 180750 241032 188986 241088
rect 189042 241032 190470 241088
rect 180750 241030 190470 241032
rect -960 240940 480 241030
rect 3509 241027 3575 241030
rect 188981 241027 189047 241030
rect 173249 240954 173315 240957
rect 187693 240954 187759 240957
rect 173249 240952 187759 240954
rect 173249 240896 173254 240952
rect 173310 240896 187698 240952
rect 187754 240896 187759 240952
rect 173249 240894 187759 240896
rect 190410 240954 190470 241030
rect 238753 241088 258323 241090
rect 238753 241032 238758 241088
rect 238814 241032 258262 241088
rect 258318 241032 258323 241088
rect 238753 241030 258323 241032
rect 238753 241027 238819 241030
rect 258257 241027 258323 241030
rect 210366 240954 210372 240956
rect 190410 240894 210372 240954
rect 173249 240891 173315 240894
rect 187693 240891 187759 240894
rect 210366 240892 210372 240894
rect 210436 240954 210442 240956
rect 255405 240954 255471 240957
rect 259729 240954 259795 240957
rect 210436 240894 248430 240954
rect 210436 240892 210442 240894
rect 187601 240818 187667 240821
rect 244273 240818 244339 240821
rect 187601 240816 244339 240818
rect 187601 240760 187606 240816
rect 187662 240760 244278 240816
rect 244334 240760 244339 240816
rect 187601 240758 244339 240760
rect 248370 240818 248430 240894
rect 255405 240952 259795 240954
rect 255405 240896 255410 240952
rect 255466 240896 259734 240952
rect 259790 240896 259795 240952
rect 255405 240894 259795 240896
rect 255405 240891 255471 240894
rect 259729 240891 259795 240894
rect 255589 240818 255655 240821
rect 248370 240816 255655 240818
rect 248370 240760 255594 240816
rect 255650 240760 255655 240816
rect 248370 240758 255655 240760
rect 187601 240755 187667 240758
rect 244273 240755 244339 240758
rect 255589 240755 255655 240758
rect 257337 240818 257403 240821
rect 262070 240818 262076 240820
rect 257337 240816 262076 240818
rect 257337 240760 257342 240816
rect 257398 240760 262076 240816
rect 257337 240758 262076 240760
rect 257337 240755 257403 240758
rect 262070 240756 262076 240758
rect 262140 240756 262146 240820
rect 62021 240274 62087 240277
rect 66294 240274 66300 240276
rect 62021 240272 66300 240274
rect 62021 240216 62026 240272
rect 62082 240216 66300 240272
rect 62021 240214 66300 240216
rect 62021 240211 62087 240214
rect 66294 240212 66300 240214
rect 66364 240212 66370 240276
rect 91001 240274 91067 240277
rect 93894 240274 93900 240276
rect 91001 240272 93900 240274
rect 91001 240216 91006 240272
rect 91062 240216 93900 240272
rect 91001 240214 93900 240216
rect 91001 240211 91067 240214
rect 93894 240212 93900 240214
rect 93964 240212 93970 240276
rect 70894 240076 70900 240140
rect 70964 240138 70970 240140
rect 71313 240138 71379 240141
rect 70964 240136 71379 240138
rect 70964 240080 71318 240136
rect 71374 240080 71379 240136
rect 70964 240078 71379 240080
rect 70964 240076 70970 240078
rect 71313 240075 71379 240078
rect 72233 240138 72299 240141
rect 72734 240138 72740 240140
rect 72233 240136 72740 240138
rect 72233 240080 72238 240136
rect 72294 240080 72740 240136
rect 72233 240078 72740 240080
rect 72233 240075 72299 240078
rect 72734 240076 72740 240078
rect 72804 240076 72810 240140
rect 74901 240138 74967 240141
rect 74490 240136 74967 240138
rect 74490 240080 74906 240136
rect 74962 240080 74967 240136
rect 74490 240078 74967 240080
rect 69197 240002 69263 240005
rect 74490 240002 74550 240078
rect 74901 240075 74967 240078
rect 88241 240138 88307 240141
rect 88701 240138 88767 240141
rect 88241 240136 88767 240138
rect 88241 240080 88246 240136
rect 88302 240080 88706 240136
rect 88762 240080 88767 240136
rect 88241 240078 88767 240080
rect 88241 240075 88307 240078
rect 88701 240075 88767 240078
rect 96889 240138 96955 240141
rect 97758 240138 97764 240140
rect 96889 240136 97764 240138
rect 96889 240080 96894 240136
rect 96950 240080 97764 240136
rect 96889 240078 97764 240080
rect 96889 240075 96955 240078
rect 97758 240076 97764 240078
rect 97828 240076 97834 240140
rect 98729 240138 98795 240141
rect 104801 240138 104867 240141
rect 177941 240138 178007 240141
rect 98729 240136 180810 240138
rect 98729 240080 98734 240136
rect 98790 240080 104806 240136
rect 104862 240080 177946 240136
rect 178002 240080 180810 240136
rect 98729 240078 180810 240080
rect 98729 240075 98795 240078
rect 104801 240075 104867 240078
rect 177941 240075 178007 240078
rect 69197 240000 74550 240002
rect 69197 239944 69202 240000
rect 69258 239944 74550 240000
rect 69197 239942 74550 239944
rect 87505 240002 87571 240005
rect 88149 240002 88215 240005
rect 87505 240000 88215 240002
rect 87505 239944 87510 240000
rect 87566 239944 88154 240000
rect 88210 239944 88215 240000
rect 87505 239942 88215 239944
rect 180750 240002 180810 240078
rect 188838 240076 188844 240140
rect 188908 240138 188914 240140
rect 188981 240138 189047 240141
rect 203006 240138 203012 240140
rect 188908 240136 189047 240138
rect 188908 240080 188986 240136
rect 189042 240080 189047 240136
rect 188908 240078 189047 240080
rect 188908 240076 188914 240078
rect 188981 240075 189047 240078
rect 200070 240078 203012 240138
rect 197997 240002 198063 240005
rect 180750 240000 198063 240002
rect 180750 239944 198002 240000
rect 198058 239944 198063 240000
rect 180750 239942 198063 239944
rect 69197 239939 69263 239942
rect 87505 239939 87571 239942
rect 88149 239939 88215 239942
rect 197997 239939 198063 239942
rect 65977 239866 66043 239869
rect 74809 239866 74875 239869
rect 75453 239866 75519 239869
rect 65977 239864 75519 239866
rect 65977 239808 65982 239864
rect 66038 239808 74814 239864
rect 74870 239808 75458 239864
rect 75514 239808 75519 239864
rect 65977 239806 75519 239808
rect 65977 239803 66043 239806
rect 74809 239803 74875 239806
rect 75453 239803 75519 239806
rect 86769 239866 86835 239869
rect 88977 239866 89043 239869
rect 86769 239864 89043 239866
rect 86769 239808 86774 239864
rect 86830 239808 88982 239864
rect 89038 239808 89043 239864
rect 86769 239806 89043 239808
rect 86769 239803 86835 239806
rect 88977 239803 89043 239806
rect 188337 239866 188403 239869
rect 200070 239866 200130 240078
rect 203006 240076 203012 240078
rect 203076 240138 203082 240140
rect 204253 240138 204319 240141
rect 203076 240136 204319 240138
rect 203076 240080 204258 240136
rect 204314 240080 204319 240136
rect 203076 240078 204319 240080
rect 203076 240076 203082 240078
rect 204253 240075 204319 240078
rect 209773 240138 209839 240141
rect 210550 240138 210556 240140
rect 209773 240136 210556 240138
rect 209773 240080 209778 240136
rect 209834 240080 210556 240136
rect 209773 240078 210556 240080
rect 209773 240075 209839 240078
rect 210550 240076 210556 240078
rect 210620 240076 210626 240140
rect 229093 240138 229159 240141
rect 229686 240138 229692 240140
rect 229093 240136 229692 240138
rect 229093 240080 229098 240136
rect 229154 240080 229692 240136
rect 229093 240078 229692 240080
rect 229093 240075 229159 240078
rect 229686 240076 229692 240078
rect 229756 240076 229762 240140
rect 234613 240138 234679 240141
rect 234838 240138 234844 240140
rect 234613 240136 234844 240138
rect 234613 240080 234618 240136
rect 234674 240080 234844 240136
rect 234613 240078 234844 240080
rect 234613 240075 234679 240078
rect 234838 240076 234844 240078
rect 234908 240076 234914 240140
rect 238886 240076 238892 240140
rect 238956 240138 238962 240140
rect 241605 240138 241671 240141
rect 238956 240136 241671 240138
rect 238956 240080 241610 240136
rect 241666 240080 241671 240136
rect 238956 240078 241671 240080
rect 238956 240076 238962 240078
rect 241605 240075 241671 240078
rect 250437 240138 250503 240141
rect 263726 240138 263732 240140
rect 250437 240136 263732 240138
rect 250437 240080 250442 240136
rect 250498 240080 263732 240136
rect 250437 240078 263732 240080
rect 250437 240075 250503 240078
rect 263726 240076 263732 240078
rect 263796 240076 263802 240140
rect 216438 239940 216444 240004
rect 216508 240002 216514 240004
rect 252737 240002 252803 240005
rect 216508 240000 252803 240002
rect 216508 239944 252742 240000
rect 252798 239944 252803 240000
rect 216508 239942 252803 239944
rect 216508 239940 216514 239942
rect 252737 239939 252803 239942
rect 188337 239864 200130 239866
rect 188337 239808 188342 239864
rect 188398 239808 200130 239864
rect 188337 239806 200130 239808
rect 188337 239803 188403 239806
rect 224166 239804 224172 239868
rect 224236 239866 224242 239868
rect 251265 239866 251331 239869
rect 224236 239864 251331 239866
rect 224236 239808 251270 239864
rect 251326 239808 251331 239864
rect 224236 239806 251331 239808
rect 224236 239804 224242 239806
rect 251265 239803 251331 239806
rect 178861 239730 178927 239733
rect 218697 239730 218763 239733
rect 178861 239728 218763 239730
rect 178861 239672 178866 239728
rect 178922 239672 218702 239728
rect 218758 239672 218763 239728
rect 178861 239670 218763 239672
rect 178861 239667 178927 239670
rect 218697 239667 218763 239670
rect 248413 239730 248479 239733
rect 257245 239730 257311 239733
rect 248413 239728 257311 239730
rect 248413 239672 248418 239728
rect 248474 239672 257250 239728
rect 257306 239672 257311 239728
rect 248413 239670 257311 239672
rect 248413 239667 248479 239670
rect 257245 239667 257311 239670
rect 204253 239458 204319 239461
rect 228541 239458 228607 239461
rect 204253 239456 228607 239458
rect 204253 239400 204258 239456
rect 204314 239400 228546 239456
rect 228602 239400 228607 239456
rect 204253 239398 228607 239400
rect 204253 239395 204319 239398
rect 228541 239395 228607 239398
rect 82169 238914 82235 238917
rect 84837 238914 84903 238917
rect 82169 238912 84903 238914
rect 82169 238856 82174 238912
rect 82230 238856 84842 238912
rect 84898 238856 84903 238912
rect 82169 238854 84903 238856
rect 82169 238851 82235 238854
rect 84837 238851 84903 238854
rect 84101 238778 84167 238781
rect 84694 238778 84700 238780
rect 84101 238776 84700 238778
rect 84101 238720 84106 238776
rect 84162 238720 84700 238776
rect 84101 238718 84700 238720
rect 84101 238715 84167 238718
rect 84694 238716 84700 238718
rect 84764 238716 84770 238780
rect 230238 238716 230244 238780
rect 230308 238778 230314 238780
rect 233877 238778 233943 238781
rect 230308 238776 233943 238778
rect 230308 238720 233882 238776
rect 233938 238720 233943 238776
rect 230308 238718 233943 238720
rect 230308 238716 230314 238718
rect 233877 238715 233943 238718
rect 78765 238642 78831 238645
rect 102777 238642 102843 238645
rect 78765 238640 102843 238642
rect 78765 238584 78770 238640
rect 78826 238584 102782 238640
rect 102838 238584 102843 238640
rect 78765 238582 102843 238584
rect 78765 238579 78831 238582
rect 102777 238579 102843 238582
rect 182081 238642 182147 238645
rect 254526 238642 254532 238644
rect 182081 238640 254532 238642
rect 182081 238584 182086 238640
rect 182142 238584 254532 238640
rect 182081 238582 254532 238584
rect 182081 238579 182147 238582
rect 254526 238580 254532 238582
rect 254596 238580 254602 238644
rect 95141 238098 95207 238101
rect 115289 238098 115355 238101
rect 95141 238096 115355 238098
rect 95141 238040 95146 238096
rect 95202 238040 115294 238096
rect 115350 238040 115355 238096
rect 95141 238038 115355 238040
rect 95141 238035 95207 238038
rect 115289 238035 115355 238038
rect 166533 238098 166599 238101
rect 216438 238098 216444 238100
rect 166533 238096 216444 238098
rect 166533 238040 166538 238096
rect 166594 238040 216444 238096
rect 166533 238038 216444 238040
rect 166533 238035 166599 238038
rect 216438 238036 216444 238038
rect 216508 238036 216514 238100
rect 111558 237900 111564 237964
rect 111628 237962 111634 237964
rect 188429 237962 188495 237965
rect 111628 237960 188495 237962
rect 111628 237904 188434 237960
rect 188490 237904 188495 237960
rect 111628 237902 188495 237904
rect 111628 237900 111634 237902
rect 188429 237899 188495 237902
rect 192477 237962 192543 237965
rect 201534 237962 201540 237964
rect 192477 237960 201540 237962
rect 192477 237904 192482 237960
rect 192538 237904 201540 237960
rect 192477 237902 201540 237904
rect 192477 237899 192543 237902
rect 201534 237900 201540 237902
rect 201604 237900 201610 237964
rect 205398 237900 205404 237964
rect 205468 237962 205474 237964
rect 245694 237962 245700 237964
rect 205468 237902 245700 237962
rect 205468 237900 205474 237902
rect 245694 237900 245700 237902
rect 245764 237900 245770 237964
rect 246389 237962 246455 237965
rect 265750 237962 265756 237964
rect 246389 237960 265756 237962
rect 246389 237904 246394 237960
rect 246450 237904 265756 237960
rect 246389 237902 265756 237904
rect 246389 237899 246455 237902
rect 265750 237900 265756 237902
rect 265820 237900 265826 237964
rect 71681 237554 71747 237557
rect 73102 237554 73108 237556
rect 71681 237552 73108 237554
rect 71681 237496 71686 237552
rect 71742 237496 73108 237552
rect 71681 237494 73108 237496
rect 71681 237491 71747 237494
rect 73102 237492 73108 237494
rect 73172 237492 73178 237556
rect 93710 237492 93716 237556
rect 93780 237554 93786 237556
rect 94221 237554 94287 237557
rect 93780 237552 94287 237554
rect 93780 237496 94226 237552
rect 94282 237496 94287 237552
rect 93780 237494 94287 237496
rect 93780 237492 93786 237494
rect 94221 237491 94287 237494
rect 53465 237418 53531 237421
rect 53649 237418 53715 237421
rect 166533 237418 166599 237421
rect 166901 237418 166967 237421
rect 53465 237416 166967 237418
rect 53465 237360 53470 237416
rect 53526 237360 53654 237416
rect 53710 237360 166538 237416
rect 166594 237360 166906 237416
rect 166962 237360 166967 237416
rect 53465 237358 166967 237360
rect 53465 237355 53531 237358
rect 53649 237355 53715 237358
rect 166533 237355 166599 237358
rect 166901 237355 166967 237358
rect 184289 236874 184355 236877
rect 202229 236874 202295 236877
rect 184289 236872 202295 236874
rect 184289 236816 184294 236872
rect 184350 236816 202234 236872
rect 202290 236816 202295 236872
rect 184289 236814 202295 236816
rect 184289 236811 184355 236814
rect 202229 236811 202295 236814
rect 77569 236738 77635 236741
rect 104709 236738 104775 236741
rect 106365 236738 106431 236741
rect 77569 236736 106431 236738
rect 77569 236680 77574 236736
rect 77630 236680 104714 236736
rect 104770 236680 106370 236736
rect 106426 236680 106431 236736
rect 77569 236678 106431 236680
rect 77569 236675 77635 236678
rect 104709 236675 104775 236678
rect 106365 236675 106431 236678
rect 175181 236738 175247 236741
rect 258390 236738 258396 236740
rect 175181 236736 258396 236738
rect 175181 236680 175186 236736
rect 175242 236680 258396 236736
rect 175181 236678 258396 236680
rect 175181 236675 175247 236678
rect 258390 236676 258396 236678
rect 258460 236676 258466 236740
rect 15101 236602 15167 236605
rect 189993 236602 190059 236605
rect 15101 236600 190059 236602
rect 15101 236544 15106 236600
rect 15162 236544 189998 236600
rect 190054 236544 190059 236600
rect 15101 236542 190059 236544
rect 15101 236539 15167 236542
rect 189993 236539 190059 236542
rect 228449 236602 228515 236605
rect 255405 236602 255471 236605
rect 228449 236600 255471 236602
rect 228449 236544 228454 236600
rect 228510 236544 255410 236600
rect 255466 236544 255471 236600
rect 228449 236542 255471 236544
rect 228449 236539 228515 236542
rect 255405 236539 255471 236542
rect 104157 236058 104223 236061
rect 106549 236058 106615 236061
rect 104157 236056 106615 236058
rect 104157 236000 104162 236056
rect 104218 236000 106554 236056
rect 106610 236000 106615 236056
rect 104157 235998 106615 236000
rect 104157 235995 104223 235998
rect 106549 235995 106615 235998
rect 80329 235922 80395 235925
rect 103513 235922 103579 235925
rect 107653 235922 107719 235925
rect 80329 235920 107719 235922
rect 80329 235864 80334 235920
rect 80390 235864 103518 235920
rect 103574 235864 107658 235920
rect 107714 235864 107719 235920
rect 80329 235862 107719 235864
rect 80329 235859 80395 235862
rect 103513 235859 103579 235862
rect 107653 235859 107719 235862
rect 177941 235922 178007 235925
rect 238753 235922 238819 235925
rect 177941 235920 238819 235922
rect 177941 235864 177946 235920
rect 178002 235864 238758 235920
rect 238814 235864 238819 235920
rect 177941 235862 238819 235864
rect 177941 235859 178007 235862
rect 238753 235859 238819 235862
rect 196617 235786 196683 235789
rect 200614 235786 200620 235788
rect 196617 235784 200620 235786
rect 196617 235728 196622 235784
rect 196678 235728 200620 235784
rect 196617 235726 200620 235728
rect 196617 235723 196683 235726
rect 200614 235724 200620 235726
rect 200684 235724 200690 235788
rect 202229 235786 202295 235789
rect 202781 235786 202847 235789
rect 263542 235786 263548 235788
rect 202229 235784 263548 235786
rect 202229 235728 202234 235784
rect 202290 235728 202786 235784
rect 202842 235728 263548 235784
rect 202229 235726 263548 235728
rect 202229 235723 202295 235726
rect 202781 235723 202847 235726
rect 263542 235724 263548 235726
rect 263612 235724 263618 235788
rect 172605 235650 172671 235653
rect 229870 235650 229876 235652
rect 172605 235648 229876 235650
rect 172605 235592 172610 235648
rect 172666 235592 229876 235648
rect 172605 235590 229876 235592
rect 172605 235587 172671 235590
rect 229870 235588 229876 235590
rect 229940 235588 229946 235652
rect 64781 235378 64847 235381
rect 158069 235378 158135 235381
rect 64781 235376 158135 235378
rect 64781 235320 64786 235376
rect 64842 235320 158074 235376
rect 158130 235320 158135 235376
rect 64781 235318 158135 235320
rect 64781 235315 64847 235318
rect 158069 235315 158135 235318
rect 39941 235242 40007 235245
rect 188521 235242 188587 235245
rect 39941 235240 188587 235242
rect 39941 235184 39946 235240
rect 40002 235184 188526 235240
rect 188582 235184 188587 235240
rect 39941 235182 188587 235184
rect 39941 235179 40007 235182
rect 188521 235179 188587 235182
rect 231761 235242 231827 235245
rect 256785 235242 256851 235245
rect 231761 235240 256851 235242
rect 231761 235184 231766 235240
rect 231822 235184 256790 235240
rect 256846 235184 256851 235240
rect 231761 235182 256851 235184
rect 231761 235179 231827 235182
rect 256785 235179 256851 235182
rect 184473 234562 184539 234565
rect 273345 234562 273411 234565
rect 184473 234560 273411 234562
rect 184473 234504 184478 234560
rect 184534 234504 273350 234560
rect 273406 234504 273411 234560
rect 184473 234502 273411 234504
rect 184473 234499 184539 234502
rect 273345 234499 273411 234502
rect 94129 234018 94195 234021
rect 119337 234018 119403 234021
rect 126329 234018 126395 234021
rect 94129 234016 126395 234018
rect 94129 233960 94134 234016
rect 94190 233960 119342 234016
rect 119398 233960 126334 234016
rect 126390 233960 126395 234016
rect 94129 233958 126395 233960
rect 94129 233955 94195 233958
rect 119337 233955 119403 233958
rect 126329 233955 126395 233958
rect 153929 234018 153995 234021
rect 229829 234018 229895 234021
rect 153929 234016 229895 234018
rect 153929 233960 153934 234016
rect 153990 233960 229834 234016
rect 229890 233960 229895 234016
rect 153929 233958 229895 233960
rect 153929 233955 153995 233958
rect 229829 233955 229895 233958
rect 24761 233882 24827 233885
rect 187141 233882 187207 233885
rect 24761 233880 187207 233882
rect 24761 233824 24766 233880
rect 24822 233824 187146 233880
rect 187202 233824 187207 233880
rect 24761 233822 187207 233824
rect 24761 233819 24827 233822
rect 187141 233819 187207 233822
rect 229829 233202 229895 233205
rect 284661 233202 284727 233205
rect 229829 233200 284727 233202
rect 229829 233144 229834 233200
rect 229890 233144 284666 233200
rect 284722 233144 284727 233200
rect 229829 233142 284727 233144
rect 229829 233139 229895 233142
rect 284661 233139 284727 233142
rect 184289 232658 184355 232661
rect 250345 232658 250411 232661
rect 184289 232656 250411 232658
rect 184289 232600 184294 232656
rect 184350 232600 250350 232656
rect 250406 232600 250411 232656
rect 184289 232598 250411 232600
rect 184289 232595 184355 232598
rect 250345 232595 250411 232598
rect 6821 232522 6887 232525
rect 189809 232522 189875 232525
rect 6821 232520 189875 232522
rect 6821 232464 6826 232520
rect 6882 232464 189814 232520
rect 189870 232464 189875 232520
rect 6821 232462 189875 232464
rect 6821 232459 6887 232462
rect 189809 232459 189875 232462
rect 193029 232522 193095 232525
rect 208342 232522 208348 232524
rect 193029 232520 208348 232522
rect 193029 232464 193034 232520
rect 193090 232464 208348 232520
rect 193029 232462 208348 232464
rect 193029 232459 193095 232462
rect 208342 232460 208348 232462
rect 208412 232460 208418 232524
rect 580165 232386 580231 232389
rect 583520 232386 584960 232476
rect 580165 232384 584960 232386
rect 580165 232328 580170 232384
rect 580226 232328 584960 232384
rect 580165 232326 584960 232328
rect 580165 232323 580231 232326
rect 583520 232236 584960 232326
rect 181529 231842 181595 231845
rect 259494 231842 259500 231844
rect 181529 231840 259500 231842
rect 181529 231784 181534 231840
rect 181590 231784 259500 231840
rect 181529 231782 259500 231784
rect 181529 231779 181595 231782
rect 259494 231780 259500 231782
rect 259564 231780 259570 231844
rect 106917 231162 106983 231165
rect 236678 231162 236684 231164
rect 106917 231160 236684 231162
rect 106917 231104 106922 231160
rect 106978 231104 236684 231160
rect 106917 231102 236684 231104
rect 106917 231099 106983 231102
rect 236678 231100 236684 231102
rect 236748 231100 236754 231164
rect 180241 230482 180307 230485
rect 251909 230482 251975 230485
rect 180241 230480 251975 230482
rect 180241 230424 180246 230480
rect 180302 230424 251914 230480
rect 251970 230424 251975 230480
rect 180241 230422 251975 230424
rect 180241 230419 180307 230422
rect 251909 230419 251975 230422
rect 222285 230346 222351 230349
rect 222694 230346 222700 230348
rect 222285 230344 222700 230346
rect 222285 230288 222290 230344
rect 222346 230288 222700 230344
rect 222285 230286 222700 230288
rect 222285 230283 222351 230286
rect 222694 230284 222700 230286
rect 222764 230284 222770 230348
rect 223430 229876 223436 229940
rect 223500 229938 223506 229940
rect 252645 229938 252711 229941
rect 223500 229936 252711 229938
rect 223500 229880 252650 229936
rect 252706 229880 252711 229936
rect 223500 229878 252711 229880
rect 223500 229876 223506 229878
rect 252645 229875 252711 229878
rect 49601 229802 49667 229805
rect 226558 229802 226564 229804
rect 49601 229800 226564 229802
rect 49601 229744 49606 229800
rect 49662 229744 226564 229800
rect 49601 229742 226564 229744
rect 49601 229739 49667 229742
rect 226558 229740 226564 229742
rect 226628 229740 226634 229804
rect 206369 229122 206435 229125
rect 211654 229122 211660 229124
rect 206369 229120 211660 229122
rect 206369 229064 206374 229120
rect 206430 229064 211660 229120
rect 206369 229062 211660 229064
rect 206369 229059 206435 229062
rect 211654 229060 211660 229062
rect 211724 229060 211730 229124
rect 61878 228924 61884 228988
rect 61948 228986 61954 228988
rect 179321 228986 179387 228989
rect 184289 228986 184355 228989
rect 61948 228984 184355 228986
rect 61948 228928 179326 228984
rect 179382 228928 184294 228984
rect 184350 228928 184355 228984
rect 61948 228926 184355 228928
rect 61948 228924 61954 228926
rect 179321 228923 179387 228926
rect 184289 228923 184355 228926
rect 220077 228986 220143 228989
rect 250437 228986 250503 228989
rect 220077 228984 250503 228986
rect 220077 228928 220082 228984
rect 220138 228928 250442 228984
rect 250498 228928 250503 228984
rect 220077 228926 250503 228928
rect 220077 228923 220143 228926
rect 250437 228923 250503 228926
rect 198641 228442 198707 228445
rect 206134 228442 206140 228444
rect 198641 228440 206140 228442
rect 198641 228384 198646 228440
rect 198702 228384 206140 228440
rect 198641 228382 206140 228384
rect 198641 228379 198707 228382
rect 206134 228380 206140 228382
rect 206204 228380 206210 228444
rect 240041 228442 240107 228445
rect 262254 228442 262260 228444
rect 240041 228440 262260 228442
rect 240041 228384 240046 228440
rect 240102 228384 262260 228440
rect 240041 228382 262260 228384
rect 240041 228379 240107 228382
rect 262254 228380 262260 228382
rect 262324 228380 262330 228444
rect 180057 228306 180123 228309
rect 198733 228306 198799 228309
rect 266486 228306 266492 228308
rect 180057 228304 266492 228306
rect 180057 228248 180062 228304
rect 180118 228248 198738 228304
rect 198794 228248 266492 228304
rect 180057 228246 266492 228248
rect 180057 228243 180123 228246
rect 198733 228243 198799 228246
rect 266486 228244 266492 228246
rect 266556 228244 266562 228308
rect -960 227884 480 228124
rect 184054 227700 184060 227764
rect 184124 227762 184130 227764
rect 184289 227762 184355 227765
rect 184124 227760 184355 227762
rect 184124 227704 184294 227760
rect 184350 227704 184355 227760
rect 184124 227702 184355 227704
rect 184124 227700 184130 227702
rect 184289 227699 184355 227702
rect 220077 227762 220143 227765
rect 220670 227762 220676 227764
rect 220077 227760 220676 227762
rect 220077 227704 220082 227760
rect 220138 227704 220676 227760
rect 220077 227702 220676 227704
rect 220077 227699 220143 227702
rect 220670 227700 220676 227702
rect 220740 227700 220746 227764
rect 237373 227082 237439 227085
rect 266629 227082 266695 227085
rect 237373 227080 266695 227082
rect 237373 227024 237378 227080
rect 237434 227024 266634 227080
rect 266690 227024 266695 227080
rect 237373 227022 266695 227024
rect 237373 227019 237439 227022
rect 266629 227019 266695 227022
rect 110321 226946 110387 226949
rect 237598 226946 237604 226948
rect 110321 226944 237604 226946
rect 110321 226888 110326 226944
rect 110382 226888 237604 226944
rect 110321 226886 237604 226888
rect 110321 226883 110387 226886
rect 237598 226884 237604 226886
rect 237668 226884 237674 226948
rect 240726 226884 240732 226948
rect 240796 226946 240802 226948
rect 248413 226946 248479 226949
rect 240796 226944 248479 226946
rect 240796 226888 248418 226944
rect 248474 226888 248479 226944
rect 240796 226886 248479 226888
rect 240796 226884 240802 226886
rect 248413 226883 248479 226886
rect 65793 226402 65859 226405
rect 66110 226402 66116 226404
rect 65793 226400 66116 226402
rect 65793 226344 65798 226400
rect 65854 226344 66116 226400
rect 65793 226342 66116 226344
rect 65793 226339 65859 226342
rect 66110 226340 66116 226342
rect 66180 226340 66186 226404
rect 180057 226266 180123 226269
rect 180609 226266 180675 226269
rect 246297 226266 246363 226269
rect 180057 226264 246363 226266
rect 180057 226208 180062 226264
rect 180118 226208 180614 226264
rect 180670 226208 246302 226264
rect 246358 226208 246363 226264
rect 180057 226206 246363 226208
rect 180057 226203 180123 226206
rect 180609 226203 180675 226206
rect 246297 226203 246363 226206
rect 119981 225722 120047 225725
rect 238518 225722 238524 225724
rect 119981 225720 238524 225722
rect 119981 225664 119986 225720
rect 120042 225664 238524 225720
rect 119981 225662 238524 225664
rect 119981 225659 120047 225662
rect 238518 225660 238524 225662
rect 238588 225660 238594 225724
rect 48221 225586 48287 225589
rect 207054 225586 207060 225588
rect 48221 225584 207060 225586
rect 48221 225528 48226 225584
rect 48282 225528 207060 225584
rect 48221 225526 207060 225528
rect 48221 225523 48287 225526
rect 207054 225524 207060 225526
rect 207124 225524 207130 225588
rect 115197 224906 115263 224909
rect 240225 224906 240291 224909
rect 115197 224904 240291 224906
rect 115197 224848 115202 224904
rect 115258 224848 240230 224904
rect 240286 224848 240291 224904
rect 115197 224846 240291 224848
rect 115197 224843 115263 224846
rect 240225 224843 240291 224846
rect 189901 224770 189967 224773
rect 253054 224770 253060 224772
rect 189901 224768 253060 224770
rect 189901 224712 189906 224768
rect 189962 224712 253060 224768
rect 189901 224710 253060 224712
rect 189901 224707 189967 224710
rect 253054 224708 253060 224710
rect 253124 224708 253130 224772
rect 38561 224226 38627 224229
rect 220854 224226 220860 224228
rect 38561 224224 220860 224226
rect 38561 224168 38566 224224
rect 38622 224168 220860 224224
rect 38561 224166 220860 224168
rect 38561 224163 38627 224166
rect 220854 224164 220860 224166
rect 220924 224164 220930 224228
rect 222101 223002 222167 223005
rect 259678 223002 259684 223004
rect 222101 223000 259684 223002
rect 222101 222944 222106 223000
rect 222162 222944 259684 223000
rect 222101 222942 259684 222944
rect 222101 222939 222167 222942
rect 259678 222940 259684 222942
rect 259748 222940 259754 223004
rect 115197 222866 115263 222869
rect 237373 222866 237439 222869
rect 238661 222866 238727 222869
rect 262806 222866 262812 222868
rect 115197 222864 219450 222866
rect 115197 222808 115202 222864
rect 115258 222808 219450 222864
rect 115197 222806 219450 222808
rect 115197 222803 115263 222806
rect 219390 222730 219450 222806
rect 237373 222864 262812 222866
rect 237373 222808 237378 222864
rect 237434 222808 238666 222864
rect 238722 222808 262812 222864
rect 237373 222806 262812 222808
rect 237373 222803 237439 222806
rect 238661 222803 238727 222806
rect 262806 222804 262812 222806
rect 262876 222804 262882 222868
rect 237782 222730 237788 222732
rect 219390 222670 237788 222730
rect 237782 222668 237788 222670
rect 237852 222668 237858 222732
rect 105537 221642 105603 221645
rect 211153 221642 211219 221645
rect 105537 221640 211219 221642
rect 105537 221584 105542 221640
rect 105598 221584 211158 221640
rect 211214 221584 211219 221640
rect 105537 221582 211219 221584
rect 105537 221579 105603 221582
rect 211153 221579 211219 221582
rect 19241 221506 19307 221509
rect 222285 221506 222351 221509
rect 19241 221504 222351 221506
rect 19241 221448 19246 221504
rect 19302 221448 222290 221504
rect 222346 221448 222351 221504
rect 19241 221446 222351 221448
rect 19241 221443 19307 221446
rect 222285 221443 222351 221446
rect 173249 220282 173315 220285
rect 273529 220282 273595 220285
rect 173249 220280 273595 220282
rect 173249 220224 173254 220280
rect 173310 220224 273534 220280
rect 273590 220224 273595 220280
rect 173249 220222 273595 220224
rect 173249 220219 173315 220222
rect 273529 220219 273595 220222
rect 4061 220146 4127 220149
rect 186814 220146 186820 220148
rect 4061 220144 186820 220146
rect 4061 220088 4066 220144
rect 4122 220088 186820 220144
rect 4061 220086 186820 220088
rect 4061 220083 4127 220086
rect 186814 220084 186820 220086
rect 186884 220084 186890 220148
rect 211153 219330 211219 219333
rect 212441 219330 212507 219333
rect 270718 219330 270724 219332
rect 211153 219328 270724 219330
rect 211153 219272 211158 219328
rect 211214 219272 212446 219328
rect 212502 219272 270724 219328
rect 211153 219270 270724 219272
rect 211153 219267 211219 219270
rect 212441 219267 212507 219270
rect 270718 219268 270724 219270
rect 270788 219268 270794 219332
rect 107009 219194 107075 219197
rect 213177 219194 213243 219197
rect 107009 219192 213243 219194
rect 107009 219136 107014 219192
rect 107070 219136 213182 219192
rect 213238 219136 213243 219192
rect 107009 219134 213243 219136
rect 107009 219131 107075 219134
rect 213177 219131 213243 219134
rect 253054 219132 253060 219196
rect 253124 219194 253130 219196
rect 288433 219194 288499 219197
rect 253124 219192 288499 219194
rect 253124 219136 288438 219192
rect 288494 219136 288499 219192
rect 253124 219134 288499 219136
rect 253124 219132 253130 219134
rect 288433 219131 288499 219134
rect 579889 219058 579955 219061
rect 583520 219058 584960 219148
rect 579889 219056 584960 219058
rect 579889 219000 579894 219056
rect 579950 219000 584960 219056
rect 579889 218998 584960 219000
rect 579889 218995 579955 218998
rect 583520 218908 584960 218998
rect 212574 218044 212580 218108
rect 212644 218106 212650 218108
rect 213177 218106 213243 218109
rect 212644 218104 213243 218106
rect 212644 218048 213182 218104
rect 213238 218048 213243 218104
rect 212644 218046 213243 218048
rect 212644 218044 212650 218046
rect 213177 218043 213243 218046
rect 159449 217970 159515 217973
rect 267774 217970 267780 217972
rect 159449 217968 267780 217970
rect 159449 217912 159454 217968
rect 159510 217912 267780 217968
rect 159449 217910 267780 217912
rect 159449 217907 159515 217910
rect 267774 217908 267780 217910
rect 267844 217908 267850 217972
rect 78029 217290 78095 217293
rect 105537 217290 105603 217293
rect 78029 217288 105603 217290
rect 78029 217232 78034 217288
rect 78090 217232 105542 217288
rect 105598 217232 105603 217288
rect 78029 217230 105603 217232
rect 78029 217227 78095 217230
rect 105537 217227 105603 217230
rect 114461 217290 114527 217293
rect 180149 217290 180215 217293
rect 114461 217288 180215 217290
rect 114461 217232 114466 217288
rect 114522 217232 180154 217288
rect 180210 217232 180215 217288
rect 114461 217230 180215 217232
rect 114461 217227 114527 217230
rect 180149 217227 180215 217230
rect 192702 217228 192708 217292
rect 192772 217290 192778 217292
rect 223757 217290 223823 217293
rect 192772 217288 223823 217290
rect 192772 217232 223762 217288
rect 223818 217232 223823 217288
rect 192772 217230 223823 217232
rect 192772 217228 192778 217230
rect 223757 217227 223823 217230
rect 76649 216066 76715 216069
rect 187693 216066 187759 216069
rect 76649 216064 187759 216066
rect 76649 216008 76654 216064
rect 76710 216008 187698 216064
rect 187754 216008 187759 216064
rect 76649 216006 187759 216008
rect 76649 216003 76715 216006
rect 187693 216003 187759 216006
rect 57830 215868 57836 215932
rect 57900 215930 57906 215932
rect 180057 215930 180123 215933
rect 57900 215928 180123 215930
rect 57900 215872 180062 215928
rect 180118 215872 180123 215928
rect 57900 215870 180123 215872
rect 57900 215868 57906 215870
rect 180057 215867 180123 215870
rect 190310 215868 190316 215932
rect 190380 215930 190386 215932
rect 582373 215930 582439 215933
rect 190380 215928 582439 215930
rect 190380 215872 582378 215928
rect 582434 215872 582439 215928
rect 190380 215870 582439 215872
rect 190380 215868 190386 215870
rect 582373 215867 582439 215870
rect 75913 215386 75979 215389
rect 76649 215386 76715 215389
rect 75913 215384 76715 215386
rect 75913 215328 75918 215384
rect 75974 215328 76654 215384
rect 76710 215328 76715 215384
rect 75913 215326 76715 215328
rect 75913 215323 75979 215326
rect 76649 215323 76715 215326
rect 187693 215386 187759 215389
rect 188337 215386 188403 215389
rect 187693 215384 188403 215386
rect 187693 215328 187698 215384
rect 187754 215328 188342 215384
rect 188398 215328 188403 215384
rect 187693 215326 188403 215328
rect 187693 215323 187759 215326
rect 188337 215323 188403 215326
rect -960 214978 480 215068
rect 3417 214978 3483 214981
rect -960 214976 3483 214978
rect -960 214920 3422 214976
rect 3478 214920 3483 214976
rect -960 214918 3483 214920
rect -960 214828 480 214918
rect 3417 214915 3483 214918
rect 195237 214706 195303 214709
rect 203006 214706 203012 214708
rect 195237 214704 203012 214706
rect 195237 214648 195242 214704
rect 195298 214648 203012 214704
rect 195237 214646 203012 214648
rect 195237 214643 195303 214646
rect 203006 214644 203012 214646
rect 203076 214644 203082 214708
rect 37089 214570 37155 214573
rect 183001 214570 183067 214573
rect 37089 214568 183067 214570
rect 37089 214512 37094 214568
rect 37150 214512 183006 214568
rect 183062 214512 183067 214568
rect 37089 214510 183067 214512
rect 37089 214507 37155 214510
rect 183001 214507 183067 214510
rect 198089 214570 198155 214573
rect 255262 214570 255268 214572
rect 198089 214568 255268 214570
rect 198089 214512 198094 214568
rect 198150 214512 255268 214568
rect 198089 214510 255268 214512
rect 198089 214507 198155 214510
rect 255262 214508 255268 214510
rect 255332 214508 255338 214572
rect 255957 214570 256023 214573
rect 276238 214570 276244 214572
rect 255957 214568 276244 214570
rect 255957 214512 255962 214568
rect 256018 214512 276244 214568
rect 255957 214510 276244 214512
rect 255957 214507 256023 214510
rect 276238 214508 276244 214510
rect 276308 214508 276314 214572
rect 78673 213210 78739 213213
rect 113817 213210 113883 213213
rect 258073 213210 258139 213213
rect 78673 213208 258139 213210
rect 78673 213152 78678 213208
rect 78734 213152 113822 213208
rect 113878 213152 258078 213208
rect 258134 213152 258139 213208
rect 78673 213150 258139 213152
rect 78673 213147 78739 213150
rect 113817 213147 113883 213150
rect 258073 213147 258139 213150
rect 72734 212468 72740 212532
rect 72804 212530 72810 212532
rect 258717 212530 258783 212533
rect 72804 212528 258783 212530
rect 72804 212472 258722 212528
rect 258778 212472 258783 212528
rect 72804 212470 258783 212472
rect 72804 212468 72810 212470
rect 258717 212467 258783 212470
rect 200849 211986 200915 211989
rect 254526 211986 254532 211988
rect 200849 211984 254532 211986
rect 200849 211928 200854 211984
rect 200910 211928 254532 211984
rect 200849 211926 254532 211928
rect 200849 211923 200915 211926
rect 254526 211924 254532 211926
rect 254596 211924 254602 211988
rect 104801 211850 104867 211853
rect 215886 211850 215892 211852
rect 104801 211848 215892 211850
rect 104801 211792 104806 211848
rect 104862 211792 215892 211848
rect 104801 211790 215892 211792
rect 104801 211787 104867 211790
rect 215886 211788 215892 211790
rect 215956 211788 215962 211852
rect 64638 210292 64644 210356
rect 64708 210354 64714 210356
rect 181529 210354 181595 210357
rect 64708 210352 181595 210354
rect 64708 210296 181534 210352
rect 181590 210296 181595 210352
rect 64708 210294 181595 210296
rect 64708 210292 64714 210294
rect 181529 210291 181595 210294
rect 193121 210354 193187 210357
rect 215334 210354 215340 210356
rect 193121 210352 215340 210354
rect 193121 210296 193126 210352
rect 193182 210296 215340 210352
rect 193121 210294 215340 210296
rect 193121 210291 193187 210294
rect 215334 210292 215340 210294
rect 215404 210292 215410 210356
rect 52361 209674 52427 209677
rect 175181 209674 175247 209677
rect 52361 209672 175247 209674
rect 52361 209616 52366 209672
rect 52422 209616 175186 209672
rect 175242 209616 175247 209672
rect 52361 209614 175247 209616
rect 52361 209611 52427 209614
rect 175181 209611 175247 209614
rect 113081 208994 113147 208997
rect 229093 208994 229159 208997
rect 113081 208992 229159 208994
rect 113081 208936 113086 208992
rect 113142 208936 229098 208992
rect 229154 208936 229159 208992
rect 113081 208934 229159 208936
rect 113081 208931 113147 208934
rect 229093 208931 229159 208934
rect 256049 207634 256115 207637
rect 262305 207634 262371 207637
rect 256049 207632 262371 207634
rect 256049 207576 256054 207632
rect 256110 207576 262310 207632
rect 262366 207576 262371 207632
rect 256049 207574 262371 207576
rect 256049 207571 256115 207574
rect 262305 207571 262371 207574
rect 207657 206274 207723 206277
rect 253054 206274 253060 206276
rect 207657 206272 253060 206274
rect 207657 206216 207662 206272
rect 207718 206216 253060 206272
rect 207657 206214 253060 206216
rect 207657 206211 207723 206214
rect 253054 206212 253060 206214
rect 253124 206212 253130 206276
rect 580257 205730 580323 205733
rect 583520 205730 584960 205820
rect 580257 205728 584960 205730
rect 580257 205672 580262 205728
rect 580318 205672 584960 205728
rect 580257 205670 584960 205672
rect 580257 205667 580323 205670
rect 583520 205580 584960 205670
rect 97206 204988 97212 205052
rect 97276 205050 97282 205052
rect 255313 205050 255379 205053
rect 255957 205050 256023 205053
rect 97276 205048 256023 205050
rect 97276 204992 255318 205048
rect 255374 204992 255962 205048
rect 256018 204992 256023 205048
rect 97276 204990 256023 204992
rect 97276 204988 97282 204990
rect 255313 204987 255379 204990
rect 255957 204987 256023 204990
rect 45461 204914 45527 204917
rect 226742 204914 226748 204916
rect 45461 204912 226748 204914
rect 45461 204856 45466 204912
rect 45522 204856 226748 204912
rect 45461 204854 226748 204856
rect 45461 204851 45527 204854
rect 226742 204852 226748 204854
rect 226812 204852 226818 204916
rect 23381 203554 23447 203557
rect 222326 203554 222332 203556
rect 23381 203552 222332 203554
rect 23381 203496 23386 203552
rect 23442 203496 222332 203552
rect 23381 203494 222332 203496
rect 23381 203491 23447 203494
rect 222326 203492 222332 203494
rect 222396 203492 222402 203556
rect 34421 202194 34487 202197
rect 204294 202194 204300 202196
rect 34421 202192 204300 202194
rect 34421 202136 34426 202192
rect 34482 202136 204300 202192
rect 34421 202134 204300 202136
rect 34421 202131 34487 202134
rect 204294 202132 204300 202134
rect 204364 202132 204370 202196
rect -960 201922 480 202012
rect 3233 201922 3299 201925
rect -960 201920 3299 201922
rect -960 201864 3238 201920
rect 3294 201864 3299 201920
rect -960 201862 3299 201864
rect -960 201772 480 201862
rect 3233 201859 3299 201862
rect 188889 201380 188955 201381
rect 188838 201378 188844 201380
rect 188798 201318 188844 201378
rect 188908 201376 188955 201380
rect 188950 201320 188955 201376
rect 188838 201316 188844 201318
rect 188908 201316 188955 201320
rect 188889 201315 188955 201316
rect 31661 200698 31727 200701
rect 223614 200698 223620 200700
rect 31661 200696 223620 200698
rect 31661 200640 31666 200696
rect 31722 200640 223620 200696
rect 31661 200638 223620 200640
rect 31661 200635 31727 200638
rect 223614 200636 223620 200638
rect 223684 200636 223690 200700
rect 42701 197978 42767 197981
rect 224902 197978 224908 197980
rect 42701 197976 224908 197978
rect 42701 197920 42706 197976
rect 42762 197920 224908 197976
rect 42701 197918 224908 197920
rect 42701 197915 42767 197918
rect 224902 197916 224908 197918
rect 224972 197916 224978 197980
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect 55121 189682 55187 189685
rect 227662 189682 227668 189684
rect 55121 189680 227668 189682
rect 55121 189624 55126 189680
rect 55182 189624 227668 189680
rect 55121 189622 227668 189624
rect 55121 189619 55187 189622
rect 227662 189620 227668 189622
rect 227732 189620 227738 189684
rect 228214 189620 228220 189684
rect 228284 189682 228290 189684
rect 265065 189682 265131 189685
rect 228284 189680 265131 189682
rect 228284 189624 265070 189680
rect 265126 189624 265131 189680
rect 228284 189622 265131 189624
rect 228284 189620 228290 189622
rect 265065 189619 265131 189622
rect -960 188866 480 188956
rect 3417 188866 3483 188869
rect -960 188864 3483 188866
rect -960 188808 3422 188864
rect 3478 188808 3483 188864
rect -960 188806 3483 188808
rect -960 188716 480 188806
rect 3417 188803 3483 188806
rect 203517 184242 203583 184245
rect 258390 184242 258396 184244
rect 203517 184240 258396 184242
rect 203517 184184 203522 184240
rect 203578 184184 258396 184240
rect 203517 184182 258396 184184
rect 203517 184179 203583 184182
rect 258390 184180 258396 184182
rect 258460 184180 258466 184244
rect 187550 182820 187556 182884
rect 187620 182882 187626 182884
rect 252737 182882 252803 182885
rect 187620 182880 252803 182882
rect 187620 182824 252742 182880
rect 252798 182824 252803 182880
rect 187620 182822 252803 182824
rect 187620 182820 187626 182822
rect 252737 182819 252803 182822
rect 86718 181324 86724 181388
rect 86788 181386 86794 181388
rect 115933 181386 115999 181389
rect 86788 181384 115999 181386
rect 86788 181328 115938 181384
rect 115994 181328 115999 181384
rect 86788 181326 115999 181328
rect 86788 181324 86794 181326
rect 115933 181323 115999 181326
rect 197353 181386 197419 181389
rect 269062 181386 269068 181388
rect 197353 181384 269068 181386
rect 197353 181328 197358 181384
rect 197414 181328 269068 181384
rect 197353 181326 269068 181328
rect 197353 181323 197419 181326
rect 269062 181324 269068 181326
rect 269132 181324 269138 181388
rect 169109 180026 169175 180029
rect 214414 180026 214420 180028
rect 169109 180024 214420 180026
rect 169109 179968 169114 180024
rect 169170 179968 214420 180024
rect 169109 179966 214420 179968
rect 169109 179963 169175 179966
rect 214414 179964 214420 179966
rect 214484 179964 214490 180028
rect 97942 179420 97948 179484
rect 98012 179482 98018 179484
rect 99189 179482 99255 179485
rect 98012 179480 99255 179482
rect 98012 179424 99194 179480
rect 99250 179424 99255 179480
rect 98012 179422 99255 179424
rect 98012 179420 98018 179422
rect 99189 179419 99255 179422
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect 193213 178666 193279 178669
rect 242934 178666 242940 178668
rect 193213 178664 242940 178666
rect 193213 178608 193218 178664
rect 193274 178608 242940 178664
rect 193213 178606 242940 178608
rect 193213 178603 193279 178606
rect 242934 178604 242940 178606
rect 243004 178604 243010 178668
rect 219709 177442 219775 177445
rect 220486 177442 220492 177444
rect 219709 177440 220492 177442
rect 219709 177384 219714 177440
rect 219770 177384 220492 177440
rect 219709 177382 220492 177384
rect 219709 177379 219775 177382
rect 220486 177380 220492 177382
rect 220556 177380 220562 177444
rect -960 175796 480 176036
rect 88977 175946 89043 175949
rect 89478 175946 89484 175948
rect 88977 175944 89484 175946
rect 88977 175888 88982 175944
rect 89038 175888 89484 175944
rect 88977 175886 89484 175888
rect 88977 175883 89043 175886
rect 89478 175884 89484 175886
rect 89548 175946 89554 175948
rect 212625 175946 212691 175949
rect 213177 175946 213243 175949
rect 89548 175944 213243 175946
rect 89548 175888 212630 175944
rect 212686 175888 213182 175944
rect 213238 175888 213243 175944
rect 89548 175886 213243 175888
rect 89548 175884 89554 175886
rect 212625 175883 212691 175886
rect 213177 175883 213243 175886
rect 207013 175266 207079 175269
rect 207657 175266 207723 175269
rect 207013 175264 207723 175266
rect 207013 175208 207018 175264
rect 207074 175208 207662 175264
rect 207718 175208 207723 175264
rect 207013 175206 207723 175208
rect 207013 175203 207079 175206
rect 207657 175203 207723 175206
rect 84837 174042 84903 174045
rect 207013 174042 207079 174045
rect 84837 174040 207079 174042
rect 84837 173984 84842 174040
rect 84898 173984 207018 174040
rect 207074 173984 207079 174040
rect 84837 173982 207079 173984
rect 84837 173979 84903 173982
rect 207013 173979 207079 173982
rect 88926 172484 88932 172548
rect 88996 172546 89002 172548
rect 213913 172546 213979 172549
rect 88996 172544 213979 172546
rect 88996 172488 213918 172544
rect 213974 172488 213979 172544
rect 88996 172486 213979 172488
rect 88996 172484 89002 172486
rect 213913 172483 213979 172486
rect 92473 169826 92539 169829
rect 222193 169826 222259 169829
rect 222837 169826 222903 169829
rect 92473 169824 222903 169826
rect 92473 169768 92478 169824
rect 92534 169768 222198 169824
rect 222254 169768 222842 169824
rect 222898 169768 222903 169824
rect 92473 169766 222903 169768
rect 92473 169763 92539 169766
rect 222193 169763 222259 169766
rect 222837 169763 222903 169766
rect 89805 168466 89871 168469
rect 220813 168466 220879 168469
rect 89805 168464 220879 168466
rect 89805 168408 89810 168464
rect 89866 168408 220818 168464
rect 220874 168408 220879 168464
rect 89805 168406 220879 168408
rect 89805 168403 89871 168406
rect 220813 168403 220879 168406
rect 60641 167650 60707 167653
rect 213678 167650 213684 167652
rect 60641 167648 213684 167650
rect 60641 167592 60646 167648
rect 60702 167592 213684 167648
rect 60641 167590 213684 167592
rect 60641 167587 60707 167590
rect 213678 167588 213684 167590
rect 213748 167588 213754 167652
rect 582833 165882 582899 165885
rect 583520 165882 584960 165972
rect 582833 165880 584960 165882
rect 582833 165824 582838 165880
rect 582894 165824 584960 165880
rect 582833 165822 584960 165824
rect 582833 165819 582899 165822
rect 86953 165746 87019 165749
rect 215293 165746 215359 165749
rect 86953 165744 215359 165746
rect 86953 165688 86958 165744
rect 87014 165688 215298 165744
rect 215354 165688 215359 165744
rect 583520 165732 584960 165822
rect 86953 165686 215359 165688
rect 86953 165683 87019 165686
rect 215293 165683 215359 165686
rect 74533 164386 74599 164389
rect 147029 164386 147095 164389
rect 238845 164386 238911 164389
rect 74533 164384 142170 164386
rect 74533 164328 74538 164384
rect 74594 164328 142170 164384
rect 74533 164326 142170 164328
rect 74533 164323 74599 164326
rect 142110 164250 142170 164326
rect 147029 164384 238911 164386
rect 147029 164328 147034 164384
rect 147090 164328 238850 164384
rect 238906 164328 238911 164384
rect 147029 164326 238911 164328
rect 147029 164323 147095 164326
rect 238845 164323 238911 164326
rect 200205 164250 200271 164253
rect 200849 164250 200915 164253
rect 142110 164248 200915 164250
rect 142110 164192 200210 164248
rect 200266 164192 200854 164248
rect 200910 164192 200915 164248
rect 142110 164190 200915 164192
rect 200205 164187 200271 164190
rect 200849 164187 200915 164190
rect 195973 163434 196039 163437
rect 284477 163434 284543 163437
rect 303613 163434 303679 163437
rect 195973 163432 303679 163434
rect 195973 163376 195978 163432
rect 196034 163376 284482 163432
rect 284538 163376 303618 163432
rect 303674 163376 303679 163432
rect 195973 163374 303679 163376
rect 195973 163371 196039 163374
rect 284477 163371 284543 163374
rect 303613 163371 303679 163374
rect -960 162890 480 162980
rect 3417 162890 3483 162893
rect -960 162888 3483 162890
rect -960 162832 3422 162888
rect 3478 162832 3483 162888
rect -960 162830 3483 162832
rect -960 162740 480 162830
rect 3417 162827 3483 162830
rect 61837 162890 61903 162893
rect 189717 162890 189783 162893
rect 61837 162888 189783 162890
rect 61837 162832 61842 162888
rect 61898 162832 189722 162888
rect 189778 162832 189783 162888
rect 61837 162830 189783 162832
rect 61837 162827 61903 162830
rect 189717 162827 189783 162830
rect 63217 161666 63283 161669
rect 190310 161666 190316 161668
rect 63217 161664 190316 161666
rect 63217 161608 63222 161664
rect 63278 161608 190316 161664
rect 63217 161606 190316 161608
rect 63217 161603 63283 161606
rect 190310 161604 190316 161606
rect 190380 161666 190386 161668
rect 198089 161666 198155 161669
rect 199377 161668 199443 161669
rect 190380 161664 198155 161666
rect 190380 161608 198094 161664
rect 198150 161608 198155 161664
rect 190380 161606 198155 161608
rect 190380 161604 190386 161606
rect 198089 161603 198155 161606
rect 199326 161604 199332 161668
rect 199396 161666 199443 161668
rect 199396 161664 199488 161666
rect 199438 161608 199488 161664
rect 199396 161606 199488 161608
rect 199396 161604 199443 161606
rect 199377 161603 199443 161604
rect 107009 161530 107075 161533
rect 236085 161530 236151 161533
rect 107009 161528 236151 161530
rect 107009 161472 107014 161528
rect 107070 161472 236090 161528
rect 236146 161472 236151 161528
rect 107009 161470 236151 161472
rect 107009 161467 107075 161470
rect 236085 161467 236151 161470
rect 109677 160306 109743 160309
rect 231853 160306 231919 160309
rect 109677 160304 231919 160306
rect 109677 160248 109682 160304
rect 109738 160248 231858 160304
rect 231914 160248 231919 160304
rect 109677 160246 231919 160248
rect 109677 160243 109743 160246
rect 231853 160243 231919 160246
rect 87137 160170 87203 160173
rect 215385 160170 215451 160173
rect 87137 160168 215451 160170
rect 87137 160112 87142 160168
rect 87198 160112 215390 160168
rect 215446 160112 215451 160168
rect 87137 160110 215451 160112
rect 87137 160107 87203 160110
rect 215385 160107 215451 160110
rect 203517 159354 203583 159357
rect 190410 159352 203583 159354
rect 190410 159296 203522 159352
rect 203578 159296 203583 159352
rect 190410 159294 203583 159296
rect 53465 158810 53531 158813
rect 53741 158810 53807 158813
rect 188889 158810 188955 158813
rect 190410 158810 190470 159294
rect 203517 159291 203583 159294
rect 53465 158808 190470 158810
rect 53465 158752 53470 158808
rect 53526 158752 53746 158808
rect 53802 158752 188894 158808
rect 188950 158752 190470 158808
rect 53465 158750 190470 158752
rect 53465 158747 53531 158750
rect 53741 158747 53807 158750
rect 188889 158747 188955 158750
rect 151261 157586 151327 157589
rect 224217 157586 224283 157589
rect 151261 157584 224283 157586
rect 151261 157528 151266 157584
rect 151322 157528 224222 157584
rect 224278 157528 224283 157584
rect 151261 157526 224283 157528
rect 151261 157523 151327 157526
rect 224217 157523 224283 157526
rect 75177 157450 75243 157453
rect 200297 157450 200363 157453
rect 75177 157448 200363 157450
rect 75177 157392 75182 157448
rect 75238 157392 200302 157448
rect 200358 157392 200363 157448
rect 75177 157390 200363 157392
rect 75177 157387 75243 157390
rect 200297 157387 200363 157390
rect 72877 156500 72943 156501
rect 72877 156496 72924 156500
rect 72988 156498 72994 156500
rect 72877 156440 72882 156496
rect 72877 156436 72924 156440
rect 72988 156438 73034 156498
rect 72988 156436 72994 156438
rect 72877 156435 72943 156436
rect 144177 156226 144243 156229
rect 224902 156226 224908 156228
rect 144177 156224 224908 156226
rect 144177 156168 144182 156224
rect 144238 156168 224908 156224
rect 144177 156166 224908 156168
rect 144177 156163 144243 156166
rect 224902 156164 224908 156166
rect 224972 156164 224978 156228
rect 83457 156090 83523 156093
rect 209129 156090 209195 156093
rect 83457 156088 209195 156090
rect 83457 156032 83462 156088
rect 83518 156032 209134 156088
rect 209190 156032 209195 156088
rect 83457 156030 209195 156032
rect 83457 156027 83523 156030
rect 209129 156027 209195 156030
rect 211797 155954 211863 155957
rect 212441 155954 212507 155957
rect 211797 155952 212507 155954
rect 211797 155896 211802 155952
rect 211858 155896 212446 155952
rect 212502 155896 212507 155952
rect 211797 155894 212507 155896
rect 211797 155891 211863 155894
rect 212441 155891 212507 155894
rect 195830 155212 195836 155276
rect 195900 155274 195906 155276
rect 217542 155274 217548 155276
rect 195900 155214 217548 155274
rect 195900 155212 195906 155214
rect 217542 155212 217548 155214
rect 217612 155274 217618 155276
rect 335353 155274 335419 155277
rect 217612 155272 335419 155274
rect 217612 155216 335358 155272
rect 335414 155216 335419 155272
rect 217612 155214 335419 155216
rect 217612 155212 217618 155214
rect 335353 155211 335419 155214
rect 152549 154730 152615 154733
rect 238017 154730 238083 154733
rect 152549 154728 238083 154730
rect 152549 154672 152554 154728
rect 152610 154672 238022 154728
rect 238078 154672 238083 154728
rect 152549 154670 238083 154672
rect 152549 154667 152615 154670
rect 238017 154667 238083 154670
rect 86217 154594 86283 154597
rect 209221 154594 209287 154597
rect 86217 154592 209287 154594
rect 86217 154536 86222 154592
rect 86278 154536 209226 154592
rect 209282 154536 209287 154592
rect 86217 154534 209287 154536
rect 86217 154531 86283 154534
rect 209221 154531 209287 154534
rect 211797 154594 211863 154597
rect 226374 154594 226380 154596
rect 211797 154592 226380 154594
rect 211797 154536 211802 154592
rect 211858 154536 226380 154592
rect 211797 154534 226380 154536
rect 211797 154531 211863 154534
rect 226374 154532 226380 154534
rect 226444 154532 226450 154596
rect 237373 154458 237439 154461
rect 237557 154458 237623 154461
rect 237373 154456 237623 154458
rect 237373 154400 237378 154456
rect 237434 154400 237562 154456
rect 237618 154400 237623 154456
rect 237373 154398 237623 154400
rect 237373 154395 237439 154398
rect 237557 154395 237623 154398
rect 149789 153370 149855 153373
rect 237557 153370 237623 153373
rect 149789 153368 237623 153370
rect 149789 153312 149794 153368
rect 149850 153312 237562 153368
rect 237618 153312 237623 153368
rect 149789 153310 237623 153312
rect 149789 153307 149855 153310
rect 237557 153307 237623 153310
rect 124949 153234 125015 153237
rect 229093 153234 229159 153237
rect 124949 153232 229159 153234
rect 124949 153176 124954 153232
rect 125010 153176 229098 153232
rect 229154 153176 229159 153232
rect 124949 153174 229159 153176
rect 124949 153171 125015 153174
rect 229093 153171 229159 153174
rect 192477 153098 192543 153101
rect 193806 153098 193812 153100
rect 192477 153096 193812 153098
rect 192477 153040 192482 153096
rect 192538 153040 193812 153096
rect 192477 153038 193812 153040
rect 192477 153035 192543 153038
rect 193806 153036 193812 153038
rect 193876 153036 193882 153100
rect 200297 153098 200363 153101
rect 256049 153098 256115 153101
rect 200297 153096 256115 153098
rect 200297 153040 200302 153096
rect 200358 153040 256054 153096
rect 256110 153040 256115 153096
rect 200297 153038 256115 153040
rect 200297 153035 200363 153038
rect 256049 153035 256115 153038
rect 193806 152628 193812 152692
rect 193876 152690 193882 152692
rect 218697 152690 218763 152693
rect 193876 152688 218763 152690
rect 193876 152632 218702 152688
rect 218758 152632 218763 152688
rect 193876 152630 218763 152632
rect 193876 152628 193882 152630
rect 218697 152627 218763 152630
rect 582557 152690 582623 152693
rect 583520 152690 584960 152780
rect 582557 152688 584960 152690
rect 582557 152632 582562 152688
rect 582618 152632 584960 152688
rect 582557 152630 584960 152632
rect 582557 152627 582623 152630
rect 83549 152554 83615 152557
rect 168281 152554 168347 152557
rect 201585 152554 201651 152557
rect 83549 152552 201651 152554
rect 83549 152496 83554 152552
rect 83610 152496 168286 152552
rect 168342 152496 201590 152552
rect 201646 152496 201651 152552
rect 583520 152540 584960 152630
rect 83549 152494 201651 152496
rect 83549 152491 83615 152494
rect 168281 152491 168347 152494
rect 201585 152491 201651 152494
rect 33041 152418 33107 152421
rect 184238 152418 184244 152420
rect 33041 152416 184244 152418
rect 33041 152360 33046 152416
rect 33102 152360 184244 152416
rect 33041 152358 184244 152360
rect 33041 152355 33107 152358
rect 184238 152356 184244 152358
rect 184308 152356 184314 152420
rect 202045 152418 202111 152421
rect 238753 152418 238819 152421
rect 202045 152416 238819 152418
rect 202045 152360 202050 152416
rect 202106 152360 238758 152416
rect 238814 152360 238819 152416
rect 202045 152358 238819 152360
rect 202045 152355 202111 152358
rect 238753 152355 238819 152358
rect 209221 151738 209287 151741
rect 270493 151738 270559 151741
rect 209221 151736 270559 151738
rect 209221 151680 209226 151736
rect 209282 151680 270498 151736
rect 270554 151680 270559 151736
rect 209221 151678 270559 151680
rect 209221 151675 209287 151678
rect 270493 151675 270559 151678
rect 56409 151194 56475 151197
rect 156689 151194 156755 151197
rect 185761 151194 185827 151197
rect 56409 151192 185827 151194
rect 56409 151136 56414 151192
rect 56470 151136 156694 151192
rect 156750 151136 185766 151192
rect 185822 151136 185827 151192
rect 56409 151134 185827 151136
rect 56409 151131 56475 151134
rect 156689 151131 156755 151134
rect 185761 151131 185827 151134
rect 50705 151058 50771 151061
rect 177246 151058 177252 151060
rect 50705 151056 177252 151058
rect 50705 151000 50710 151056
rect 50766 151000 177252 151056
rect 50705 150998 177252 151000
rect 50705 150995 50771 150998
rect 177246 150996 177252 150998
rect 177316 150996 177322 151060
rect 204253 151058 204319 151061
rect 213269 151058 213335 151061
rect 204253 151056 213335 151058
rect 204253 151000 204258 151056
rect 204314 151000 213274 151056
rect 213330 151000 213335 151056
rect 204253 150998 213335 151000
rect 204253 150995 204319 150998
rect 213269 150995 213335 150998
rect 184381 150514 184447 150517
rect 230473 150514 230539 150517
rect 184381 150512 230539 150514
rect 184381 150456 184386 150512
rect 184442 150456 230478 150512
rect 230534 150456 230539 150512
rect 184381 150454 230539 150456
rect 184381 150451 184447 150454
rect 230473 150451 230539 150454
rect -960 149834 480 149924
rect 3325 149834 3391 149837
rect -960 149832 3391 149834
rect -960 149776 3330 149832
rect 3386 149776 3391 149832
rect -960 149774 3391 149776
rect -960 149684 480 149774
rect 3325 149771 3391 149774
rect 155309 149426 155375 149429
rect 240225 149426 240291 149429
rect 155309 149424 240291 149426
rect 155309 149368 155314 149424
rect 155370 149368 240230 149424
rect 240286 149368 240291 149424
rect 155309 149366 240291 149368
rect 155309 149363 155375 149366
rect 240225 149363 240291 149366
rect 82997 149290 83063 149293
rect 102777 149290 102843 149293
rect 227662 149290 227668 149292
rect 82997 149288 84210 149290
rect 82997 149232 83002 149288
rect 83058 149232 84210 149288
rect 82997 149230 84210 149232
rect 82997 149227 83063 149230
rect 66662 149092 66668 149156
rect 66732 149154 66738 149156
rect 67541 149154 67607 149157
rect 66732 149152 67607 149154
rect 66732 149096 67546 149152
rect 67602 149096 67607 149152
rect 66732 149094 67607 149096
rect 66732 149092 66738 149094
rect 67541 149091 67607 149094
rect 81341 149154 81407 149157
rect 83406 149154 83412 149156
rect 81341 149152 83412 149154
rect 81341 149096 81346 149152
rect 81402 149096 83412 149152
rect 81341 149094 83412 149096
rect 81341 149091 81407 149094
rect 83406 149092 83412 149094
rect 83476 149092 83482 149156
rect 84150 149154 84210 149230
rect 102777 149288 227668 149290
rect 102777 149232 102782 149288
rect 102838 149232 227668 149288
rect 102777 149230 227668 149232
rect 102777 149227 102843 149230
rect 227662 149228 227668 149230
rect 227732 149228 227738 149292
rect 211153 149154 211219 149157
rect 212441 149154 212507 149157
rect 84150 149152 212507 149154
rect 84150 149096 211158 149152
rect 211214 149096 212446 149152
rect 212502 149096 212507 149152
rect 84150 149094 212507 149096
rect 211153 149091 211219 149094
rect 212441 149091 212507 149094
rect 53741 148338 53807 148341
rect 185669 148338 185735 148341
rect 53741 148336 185735 148338
rect 53741 148280 53746 148336
rect 53802 148280 185674 148336
rect 185730 148280 185735 148336
rect 53741 148278 185735 148280
rect 53741 148275 53807 148278
rect 185669 148275 185735 148278
rect 187693 147930 187759 147933
rect 229185 147930 229251 147933
rect 229829 147930 229895 147933
rect 187693 147928 229895 147930
rect 187693 147872 187698 147928
rect 187754 147872 229190 147928
rect 229246 147872 229834 147928
rect 229890 147872 229895 147928
rect 187693 147870 229895 147872
rect 187693 147867 187759 147870
rect 229185 147867 229251 147870
rect 229829 147867 229895 147870
rect 126329 147794 126395 147797
rect 223614 147794 223620 147796
rect 126329 147792 223620 147794
rect 126329 147736 126334 147792
rect 126390 147736 223620 147792
rect 126329 147734 223620 147736
rect 126329 147731 126395 147734
rect 223614 147732 223620 147734
rect 223684 147732 223690 147796
rect 183001 147114 183067 147117
rect 219198 147114 219204 147116
rect 183001 147112 219204 147114
rect 183001 147056 183006 147112
rect 183062 147056 219204 147112
rect 183001 147054 219204 147056
rect 183001 147051 183067 147054
rect 219198 147052 219204 147054
rect 219268 147114 219274 147116
rect 226333 147114 226399 147117
rect 219268 147112 226399 147114
rect 219268 147056 226338 147112
rect 226394 147056 226399 147112
rect 219268 147054 226399 147056
rect 219268 147052 219274 147054
rect 226333 147051 226399 147054
rect 10961 146978 11027 146981
rect 188286 146978 188292 146980
rect 10961 146976 188292 146978
rect 10961 146920 10966 146976
rect 11022 146920 188292 146976
rect 10961 146918 188292 146920
rect 10961 146915 11027 146918
rect 188286 146916 188292 146918
rect 188356 146916 188362 146980
rect 210049 146978 210115 146981
rect 285949 146978 286015 146981
rect 210049 146976 286015 146978
rect 210049 146920 210054 146976
rect 210110 146920 285954 146976
rect 286010 146920 286015 146976
rect 210049 146918 286015 146920
rect 210049 146915 210115 146918
rect 285949 146915 286015 146918
rect 188429 146434 188495 146437
rect 188429 146432 226442 146434
rect 188429 146376 188434 146432
rect 188490 146376 226442 146432
rect 188429 146374 226442 146376
rect 188429 146371 188495 146374
rect 226382 146298 226442 146374
rect 226926 146298 226932 146300
rect 226382 146238 226932 146298
rect 226926 146236 226932 146238
rect 226996 146298 227002 146300
rect 278865 146298 278931 146301
rect 226996 146296 278931 146298
rect 226996 146240 278870 146296
rect 278926 146240 278931 146296
rect 226996 146238 278931 146240
rect 226996 146236 227002 146238
rect 278865 146235 278931 146238
rect 245653 146162 245719 146165
rect 246481 146162 246547 146165
rect 245653 146160 246547 146162
rect 245653 146104 245658 146160
rect 245714 146104 246486 146160
rect 246542 146104 246547 146160
rect 245653 146102 246547 146104
rect 245653 146099 245719 146102
rect 246481 146099 246547 146102
rect 159541 145754 159607 145757
rect 193397 145754 193463 145757
rect 159541 145752 193463 145754
rect 159541 145696 159546 145752
rect 159602 145696 193402 145752
rect 193458 145696 193463 145752
rect 159541 145694 193463 145696
rect 159541 145691 159607 145694
rect 193397 145691 193463 145694
rect 108297 145618 108363 145621
rect 187693 145618 187759 145621
rect 108297 145616 187759 145618
rect 108297 145560 108302 145616
rect 108358 145560 187698 145616
rect 187754 145560 187759 145616
rect 108297 145558 187759 145560
rect 108297 145555 108363 145558
rect 187693 145555 187759 145558
rect 185577 145074 185643 145077
rect 217225 145074 217291 145077
rect 185577 145072 217291 145074
rect 185577 145016 185582 145072
rect 185638 145016 217230 145072
rect 217286 145016 217291 145072
rect 185577 145014 217291 145016
rect 185577 145011 185643 145014
rect 217225 145011 217291 145014
rect 65793 144938 65859 144941
rect 177389 144938 177455 144941
rect 65793 144936 177455 144938
rect 65793 144880 65798 144936
rect 65854 144880 177394 144936
rect 177450 144880 177455 144936
rect 65793 144878 177455 144880
rect 65793 144875 65859 144878
rect 177389 144875 177455 144878
rect 192569 144938 192635 144941
rect 246481 144938 246547 144941
rect 192569 144936 246547 144938
rect 192569 144880 192574 144936
rect 192630 144880 246486 144936
rect 246542 144880 246547 144936
rect 192569 144878 246547 144880
rect 192569 144875 192635 144878
rect 246481 144875 246547 144878
rect 91502 144740 91508 144804
rect 91572 144802 91578 144804
rect 93117 144802 93183 144805
rect 91572 144800 93183 144802
rect 91572 144744 93122 144800
rect 93178 144744 93183 144800
rect 91572 144742 93183 144744
rect 91572 144740 91578 144742
rect 93117 144739 93183 144742
rect 155953 144802 156019 144805
rect 156689 144802 156755 144805
rect 155953 144800 156755 144802
rect 155953 144744 155958 144800
rect 156014 144744 156694 144800
rect 156750 144744 156755 144800
rect 155953 144742 156755 144744
rect 155953 144739 156019 144742
rect 156689 144739 156755 144742
rect 173341 144258 173407 144261
rect 202137 144258 202203 144261
rect 173341 144256 202203 144258
rect 173341 144200 173346 144256
rect 173402 144200 202142 144256
rect 202198 144200 202203 144256
rect 173341 144198 202203 144200
rect 173341 144195 173407 144198
rect 202137 144195 202203 144198
rect 81985 144122 82051 144125
rect 106549 144122 106615 144125
rect 81985 144120 106615 144122
rect 81985 144064 81990 144120
rect 82046 144064 106554 144120
rect 106610 144064 106615 144120
rect 81985 144062 106615 144064
rect 81985 144059 82051 144062
rect 106549 144059 106615 144062
rect 107561 144122 107627 144125
rect 186957 144122 187023 144125
rect 107561 144120 187023 144122
rect 107561 144064 107566 144120
rect 107622 144064 186962 144120
rect 187018 144064 187023 144120
rect 107561 144062 187023 144064
rect 107561 144059 107627 144062
rect 186957 144059 187023 144062
rect 208117 144122 208183 144125
rect 295425 144122 295491 144125
rect 302233 144122 302299 144125
rect 208117 144120 302299 144122
rect 208117 144064 208122 144120
rect 208178 144064 295430 144120
rect 295486 144064 302238 144120
rect 302294 144064 302299 144120
rect 208117 144062 302299 144064
rect 208117 144059 208183 144062
rect 295425 144059 295491 144062
rect 302233 144059 302299 144062
rect 209037 143850 209103 143853
rect 211654 143850 211660 143852
rect 209037 143848 211660 143850
rect 209037 143792 209042 143848
rect 209098 143792 211660 143848
rect 209037 143790 211660 143792
rect 209037 143787 209103 143790
rect 211654 143788 211660 143790
rect 211724 143788 211730 143852
rect 211245 143714 211311 143717
rect 231945 143714 232011 143717
rect 211245 143712 232011 143714
rect 211245 143656 211250 143712
rect 211306 143656 231950 143712
rect 232006 143656 232011 143712
rect 211245 143654 232011 143656
rect 211245 143651 211311 143654
rect 231945 143651 232011 143654
rect 67766 143516 67772 143580
rect 67836 143578 67842 143580
rect 156689 143578 156755 143581
rect 67836 143576 156755 143578
rect 67836 143520 156694 143576
rect 156750 143520 156755 143576
rect 67836 143518 156755 143520
rect 67836 143516 67842 143518
rect 156689 143515 156755 143518
rect 181529 143578 181595 143581
rect 223389 143578 223455 143581
rect 181529 143576 223455 143578
rect 181529 143520 181534 143576
rect 181590 143520 223394 143576
rect 223450 143520 223455 143576
rect 181529 143518 223455 143520
rect 181529 143515 181595 143518
rect 223389 143515 223455 143518
rect 104893 143442 104959 143445
rect 206277 143442 206343 143445
rect 206829 143442 206895 143445
rect 103470 143440 206895 143442
rect 103470 143384 104898 143440
rect 104954 143384 206282 143440
rect 206338 143384 206834 143440
rect 206890 143384 206895 143440
rect 103470 143382 206895 143384
rect 80053 142898 80119 142901
rect 103470 142898 103530 143382
rect 104893 143379 104959 143382
rect 206277 143379 206343 143382
rect 206829 143379 206895 143382
rect 212625 143442 212691 143445
rect 213453 143442 213519 143445
rect 212625 143440 213519 143442
rect 212625 143384 212630 143440
rect 212686 143384 213458 143440
rect 213514 143384 213519 143440
rect 212625 143382 213519 143384
rect 212625 143379 212691 143382
rect 213453 143379 213519 143382
rect 122833 143306 122899 143309
rect 206461 143306 206527 143309
rect 122833 143304 206527 143306
rect 122833 143248 122838 143304
rect 122894 143248 206466 143304
rect 206522 143248 206527 143304
rect 122833 143246 206527 143248
rect 122833 143243 122899 143246
rect 206461 143243 206527 143246
rect 197854 143108 197860 143172
rect 197924 143170 197930 143172
rect 198641 143170 198707 143173
rect 197924 143168 198707 143170
rect 197924 143112 198646 143168
rect 198702 143112 198707 143168
rect 197924 143110 198707 143112
rect 197924 143108 197930 143110
rect 198641 143107 198707 143110
rect 80053 142896 103530 142898
rect 80053 142840 80058 142896
rect 80114 142840 103530 142896
rect 80053 142838 103530 142840
rect 80053 142835 80119 142838
rect 66110 142700 66116 142764
rect 66180 142762 66186 142764
rect 76189 142762 76255 142765
rect 66180 142760 76255 142762
rect 66180 142704 76194 142760
rect 76250 142704 76255 142760
rect 66180 142702 76255 142704
rect 66180 142700 66186 142702
rect 76189 142699 76255 142702
rect 78673 142762 78739 142765
rect 122833 142762 122899 142765
rect 78673 142760 122899 142762
rect 78673 142704 78678 142760
rect 78734 142704 122838 142760
rect 122894 142704 122899 142760
rect 78673 142702 122899 142704
rect 78673 142699 78739 142702
rect 122833 142699 122899 142702
rect 224217 142354 224283 142357
rect 224217 142352 229110 142354
rect 224217 142296 224222 142352
rect 224278 142296 229110 142352
rect 224217 142294 229110 142296
rect 224217 142291 224283 142294
rect 189073 142218 189139 142221
rect 196617 142218 196683 142221
rect 189073 142216 196683 142218
rect 189073 142160 189078 142216
rect 189134 142160 196622 142216
rect 196678 142160 196683 142216
rect 189073 142158 196683 142160
rect 189073 142155 189139 142158
rect 196617 142155 196683 142158
rect 204989 142218 205055 142221
rect 219433 142218 219499 142221
rect 204989 142216 219499 142218
rect 204989 142160 204994 142216
rect 205050 142160 219438 142216
rect 219494 142160 219499 142216
rect 204989 142158 219499 142160
rect 204989 142155 205055 142158
rect 219433 142155 219499 142158
rect 221917 142218 221983 142221
rect 224718 142218 224724 142220
rect 221917 142216 224724 142218
rect 221917 142160 221922 142216
rect 221978 142160 224724 142216
rect 221917 142158 224724 142160
rect 221917 142155 221983 142158
rect 224718 142156 224724 142158
rect 224788 142156 224794 142220
rect 229050 142218 229110 142294
rect 229829 142218 229895 142221
rect 229050 142216 229895 142218
rect 229050 142160 229834 142216
rect 229890 142160 229895 142216
rect 229050 142158 229895 142160
rect 229829 142155 229895 142158
rect 83406 141476 83412 141540
rect 83476 141538 83482 141540
rect 104249 141538 104315 141541
rect 83476 141536 104315 141538
rect 83476 141480 104254 141536
rect 104310 141480 104315 141536
rect 83476 141478 104315 141480
rect 83476 141476 83482 141478
rect 104249 141475 104315 141478
rect 81341 141402 81407 141405
rect 208117 141402 208183 141405
rect 81341 141400 208183 141402
rect 81341 141344 81346 141400
rect 81402 141344 208122 141400
rect 208178 141344 208183 141400
rect 81341 141342 208183 141344
rect 81341 141339 81407 141342
rect 208117 141339 208183 141342
rect 209957 140994 210023 140997
rect 236637 140994 236703 140997
rect 209957 140992 236703 140994
rect 209957 140936 209962 140992
rect 210018 140936 236642 140992
rect 236698 140936 236703 140992
rect 209957 140934 236703 140936
rect 209957 140931 210023 140934
rect 236637 140931 236703 140934
rect 80605 140858 80671 140861
rect 81341 140858 81407 140861
rect 80605 140856 81407 140858
rect 80605 140800 80610 140856
rect 80666 140800 81346 140856
rect 81402 140800 81407 140856
rect 80605 140798 81407 140800
rect 80605 140795 80671 140798
rect 81341 140795 81407 140798
rect 214281 140858 214347 140861
rect 583017 140858 583083 140861
rect 214281 140856 583083 140858
rect 214281 140800 214286 140856
rect 214342 140800 583022 140856
rect 583078 140800 583083 140856
rect 214281 140798 583083 140800
rect 214281 140795 214347 140798
rect 583017 140795 583083 140798
rect 194593 140586 194659 140589
rect 197854 140586 197860 140588
rect 180750 140584 197860 140586
rect 180750 140528 194598 140584
rect 194654 140528 197860 140584
rect 180750 140526 197860 140528
rect 69974 140116 69980 140180
rect 70044 140178 70050 140180
rect 180750 140178 180810 140526
rect 194593 140523 194659 140526
rect 197854 140524 197860 140526
rect 197924 140524 197930 140588
rect 196566 140388 196572 140452
rect 196636 140450 196642 140452
rect 196801 140450 196867 140453
rect 196636 140448 196867 140450
rect 196636 140392 196806 140448
rect 196862 140392 196867 140448
rect 196636 140390 196867 140392
rect 196636 140388 196642 140390
rect 196801 140387 196867 140390
rect 223389 140450 223455 140453
rect 226793 140450 226859 140453
rect 223389 140448 226859 140450
rect 223389 140392 223394 140448
rect 223450 140392 226798 140448
rect 226854 140392 226859 140448
rect 223389 140390 226859 140392
rect 223389 140387 223455 140390
rect 226793 140387 226859 140390
rect 70044 140118 180810 140178
rect 70044 140116 70050 140118
rect 253289 140042 253355 140045
rect 229050 140040 253355 140042
rect 229050 139984 253294 140040
rect 253350 139984 253355 140040
rect 229050 139982 253355 139984
rect 191649 139906 191715 139909
rect 226333 139906 226399 139909
rect 229050 139906 229110 139982
rect 253289 139979 253355 139982
rect 191649 139904 193660 139906
rect 191649 139848 191654 139904
rect 191710 139848 193660 139904
rect 191649 139846 193660 139848
rect 224940 139904 229110 139906
rect 224940 139848 226338 139904
rect 226394 139848 229110 139904
rect 224940 139846 229110 139848
rect 191649 139843 191715 139846
rect 226333 139843 226399 139846
rect 64689 139634 64755 139637
rect 94814 139634 94820 139636
rect 64689 139632 94820 139634
rect 64689 139576 64694 139632
rect 64750 139576 94820 139632
rect 64689 139574 94820 139576
rect 64689 139571 64755 139574
rect 94814 139572 94820 139574
rect 94884 139572 94890 139636
rect 69289 139498 69355 139501
rect 69974 139498 69980 139500
rect 69289 139496 69980 139498
rect 69289 139440 69294 139496
rect 69350 139440 69980 139496
rect 69289 139438 69980 139440
rect 69289 139435 69355 139438
rect 69974 139436 69980 139438
rect 70044 139436 70050 139500
rect 71681 139362 71747 139365
rect 189073 139362 189139 139365
rect 71681 139360 189139 139362
rect 71681 139304 71686 139360
rect 71742 139304 189078 139360
rect 189134 139304 189139 139360
rect 71681 139302 189139 139304
rect 71681 139299 71747 139302
rect 189073 139299 189139 139302
rect 582741 139362 582807 139365
rect 583520 139362 584960 139452
rect 582741 139360 584960 139362
rect 582741 139304 582746 139360
rect 582802 139304 584960 139360
rect 582741 139302 584960 139304
rect 582741 139299 582807 139302
rect 583520 139212 584960 139302
rect 71630 138756 71636 138820
rect 71700 138818 71706 138820
rect 81433 138818 81499 138821
rect 71700 138816 81499 138818
rect 71700 138760 81438 138816
rect 81494 138760 81499 138816
rect 71700 138758 81499 138760
rect 71700 138756 71706 138758
rect 81433 138755 81499 138758
rect 81433 138682 81499 138685
rect 157977 138682 158043 138685
rect 81433 138680 158043 138682
rect 81433 138624 81438 138680
rect 81494 138624 157982 138680
rect 158038 138624 158043 138680
rect 81433 138622 158043 138624
rect 81433 138619 81499 138622
rect 157977 138619 158043 138622
rect 71129 138546 71195 138549
rect 71681 138546 71747 138549
rect 71129 138544 71747 138546
rect 71129 138488 71134 138544
rect 71190 138488 71686 138544
rect 71742 138488 71747 138544
rect 71129 138486 71747 138488
rect 71129 138483 71195 138486
rect 71681 138483 71747 138486
rect 190361 138546 190427 138549
rect 193630 138546 193690 139060
rect 190361 138544 193690 138546
rect 190361 138488 190366 138544
rect 190422 138488 193690 138544
rect 190361 138486 193690 138488
rect 224910 138546 224970 139060
rect 236085 138546 236151 138549
rect 224910 138544 236151 138546
rect 224910 138488 236090 138544
rect 236146 138488 236151 138544
rect 224910 138486 236151 138488
rect 190361 138483 190427 138486
rect 236085 138483 236151 138486
rect 69422 138348 69428 138412
rect 69492 138410 69498 138412
rect 71037 138410 71103 138413
rect 69492 138408 71103 138410
rect 69492 138352 71042 138408
rect 71098 138352 71103 138408
rect 69492 138350 71103 138352
rect 69492 138348 69498 138350
rect 71037 138347 71103 138350
rect 70025 138274 70091 138277
rect 70158 138274 70164 138276
rect 70025 138272 70164 138274
rect 70025 138216 70030 138272
rect 70086 138216 70164 138272
rect 70025 138214 70164 138216
rect 70025 138211 70091 138214
rect 70158 138212 70164 138214
rect 70228 138212 70234 138276
rect 192661 138274 192727 138277
rect 192937 138274 193003 138277
rect 226609 138274 226675 138277
rect 192661 138272 193660 138274
rect 192661 138216 192666 138272
rect 192722 138216 192942 138272
rect 192998 138216 193660 138272
rect 192661 138214 193660 138216
rect 224940 138272 226675 138274
rect 224940 138216 226614 138272
rect 226670 138216 226675 138272
rect 224940 138214 226675 138216
rect 192661 138211 192727 138214
rect 192937 138211 193003 138214
rect 226609 138211 226675 138214
rect 59169 138138 59235 138141
rect 96286 138138 96292 138140
rect 59169 138136 96292 138138
rect 59169 138080 59174 138136
rect 59230 138080 96292 138136
rect 59169 138078 96292 138080
rect 59169 138075 59235 138078
rect 96286 138076 96292 138078
rect 96356 138076 96362 138140
rect 79869 138002 79935 138005
rect 84837 138002 84903 138005
rect 79869 138000 84903 138002
rect 79869 137944 79874 138000
rect 79930 137944 84842 138000
rect 84898 137944 84903 138000
rect 79869 137942 84903 137944
rect 79869 137939 79935 137942
rect 84837 137939 84903 137942
rect 75545 137730 75611 137733
rect 83641 137730 83707 137733
rect 75545 137728 83707 137730
rect 75545 137672 75550 137728
rect 75606 137672 83646 137728
rect 83702 137672 83707 137728
rect 75545 137670 83707 137672
rect 75545 137667 75611 137670
rect 83641 137667 83707 137670
rect 194174 137668 194180 137732
rect 194244 137668 194250 137732
rect 194182 137428 194242 137668
rect 69841 137322 69907 137325
rect 80697 137322 80763 137325
rect 69841 137320 80763 137322
rect 69841 137264 69846 137320
rect 69902 137264 80702 137320
rect 80758 137264 80763 137320
rect 69841 137262 80763 137264
rect 69841 137259 69907 137262
rect 80697 137259 80763 137262
rect 89161 137322 89227 137325
rect 192477 137322 192543 137325
rect 89161 137320 192543 137322
rect 89161 137264 89166 137320
rect 89222 137264 192482 137320
rect 192538 137264 192543 137320
rect 89161 137262 192543 137264
rect 89161 137259 89227 137262
rect 192477 137259 192543 137262
rect 226609 137186 226675 137189
rect 224940 137184 226675 137186
rect 224940 137128 226614 137184
rect 226670 137128 226675 137184
rect 224940 137126 226675 137128
rect 226609 137123 226675 137126
rect 81341 136914 81407 136917
rect 86217 136914 86283 136917
rect 81341 136912 86283 136914
rect -960 136778 480 136868
rect 81341 136856 81346 136912
rect 81402 136856 86222 136912
rect 86278 136856 86283 136912
rect 81341 136854 86283 136856
rect 81341 136851 81407 136854
rect 86217 136851 86283 136854
rect 3233 136778 3299 136781
rect -960 136776 3299 136778
rect -960 136720 3238 136776
rect 3294 136720 3299 136776
rect -960 136718 3299 136720
rect -960 136628 480 136718
rect 3233 136715 3299 136718
rect 57237 136778 57303 136781
rect 75821 136778 75887 136781
rect 57237 136776 75887 136778
rect 57237 136720 57242 136776
rect 57298 136720 75826 136776
rect 75882 136720 75887 136776
rect 57237 136718 75887 136720
rect 57237 136715 57303 136718
rect 75821 136715 75887 136718
rect 82905 136778 82971 136781
rect 83406 136778 83412 136780
rect 82905 136776 83412 136778
rect 82905 136720 82910 136776
rect 82966 136720 83412 136776
rect 82905 136718 83412 136720
rect 82905 136715 82971 136718
rect 83406 136716 83412 136718
rect 83476 136716 83482 136780
rect 85481 136778 85547 136781
rect 88926 136778 88932 136780
rect 85481 136776 88932 136778
rect 85481 136720 85486 136776
rect 85542 136720 88932 136776
rect 85481 136718 88932 136720
rect 85481 136715 85547 136718
rect 88926 136716 88932 136718
rect 88996 136716 89002 136780
rect 191649 136370 191715 136373
rect 226926 136370 226932 136372
rect 191649 136368 193660 136370
rect 191649 136312 191654 136368
rect 191710 136312 193660 136368
rect 191649 136310 193660 136312
rect 224940 136310 226932 136370
rect 191649 136307 191715 136310
rect 226926 136308 226932 136310
rect 226996 136308 227002 136372
rect 96705 135962 96771 135965
rect 107009 135962 107075 135965
rect 96705 135960 107075 135962
rect 96705 135904 96710 135960
rect 96766 135904 107014 135960
rect 107070 135904 107075 135960
rect 96705 135902 107075 135904
rect 96705 135899 96771 135902
rect 107009 135899 107075 135902
rect 152641 135962 152707 135965
rect 186865 135962 186931 135965
rect 152641 135960 186931 135962
rect 152641 135904 152646 135960
rect 152702 135904 186870 135960
rect 186926 135904 186931 135960
rect 152641 135902 186931 135904
rect 152641 135899 152707 135902
rect 186865 135899 186931 135902
rect 224718 135900 224724 135964
rect 224788 135962 224794 135964
rect 276013 135962 276079 135965
rect 224788 135960 276079 135962
rect 224788 135904 276018 135960
rect 276074 135904 276079 135960
rect 224788 135902 276079 135904
rect 224788 135900 224794 135902
rect 276013 135899 276079 135902
rect 90950 135492 90956 135556
rect 91020 135554 91026 135556
rect 95233 135554 95299 135557
rect 91020 135552 95299 135554
rect 91020 135496 95238 135552
rect 95294 135496 95299 135552
rect 91020 135494 95299 135496
rect 91020 135492 91026 135494
rect 95233 135491 95299 135494
rect 191649 135554 191715 135557
rect 227662 135554 227668 135556
rect 191649 135552 193660 135554
rect 191649 135496 191654 135552
rect 191710 135496 193660 135552
rect 191649 135494 193660 135496
rect 224940 135494 227668 135554
rect 191649 135491 191715 135494
rect 227662 135492 227668 135494
rect 227732 135492 227738 135556
rect 58617 135418 58683 135421
rect 91737 135418 91803 135421
rect 58617 135416 91803 135418
rect 58617 135360 58622 135416
rect 58678 135360 91742 135416
rect 91798 135360 91803 135416
rect 58617 135358 91803 135360
rect 58617 135355 58683 135358
rect 91737 135355 91803 135358
rect 92289 135418 92355 135421
rect 95182 135418 95188 135420
rect 92289 135416 95188 135418
rect 92289 135360 92294 135416
rect 92350 135360 95188 135416
rect 92289 135358 95188 135360
rect 92289 135355 92355 135358
rect 95182 135356 95188 135358
rect 95252 135356 95258 135420
rect 69238 135220 69244 135284
rect 69308 135282 69314 135284
rect 172513 135282 172579 135285
rect 173801 135282 173867 135285
rect 69308 135280 173867 135282
rect 69308 135224 172518 135280
rect 172574 135224 173806 135280
rect 173862 135224 173867 135280
rect 69308 135222 173867 135224
rect 69308 135220 69314 135222
rect 172513 135219 172579 135222
rect 173801 135219 173867 135222
rect 188838 135084 188844 135148
rect 188908 135146 188914 135148
rect 189809 135146 189875 135149
rect 188908 135144 189875 135146
rect 188908 135088 189814 135144
rect 189870 135088 189875 135144
rect 188908 135086 189875 135088
rect 188908 135084 188914 135086
rect 189809 135083 189875 135086
rect 69565 135010 69631 135013
rect 69430 135008 69631 135010
rect 69430 134952 69570 135008
rect 69626 134952 69631 135008
rect 69430 134950 69631 134952
rect 69430 134436 69490 134950
rect 69565 134947 69631 134950
rect 72366 134676 72372 134740
rect 72436 134738 72442 134740
rect 73061 134738 73127 134741
rect 72436 134736 73127 134738
rect 72436 134680 73066 134736
rect 73122 134680 73127 134736
rect 72436 134678 73127 134680
rect 72436 134676 72442 134678
rect 73061 134675 73127 134678
rect 192477 134738 192543 134741
rect 226793 134738 226859 134741
rect 192477 134736 193660 134738
rect 192477 134680 192482 134736
rect 192538 134680 193660 134736
rect 192477 134678 193660 134680
rect 224940 134736 226859 134738
rect 224940 134680 226798 134736
rect 226854 134680 226859 134736
rect 224940 134678 226859 134680
rect 192477 134675 192543 134678
rect 226793 134675 226859 134678
rect 183001 133922 183067 133925
rect 94668 133920 183067 133922
rect 94668 133864 183006 133920
rect 183062 133864 183067 133920
rect 94668 133862 183067 133864
rect 183001 133859 183067 133862
rect 189901 133922 189967 133925
rect 189901 133920 193660 133922
rect 189901 133864 189906 133920
rect 189962 133864 193660 133920
rect 189901 133862 193660 133864
rect 189901 133859 189967 133862
rect 226609 133650 226675 133653
rect 224940 133648 226675 133650
rect 69430 133516 69490 133620
rect 224940 133592 226614 133648
rect 226670 133592 226675 133648
rect 224940 133590 226675 133592
rect 226609 133587 226675 133590
rect 69422 133452 69428 133516
rect 69492 133452 69498 133516
rect 96705 133106 96771 133109
rect 94668 133104 96771 133106
rect 94668 133048 96710 133104
rect 96766 133048 96771 133104
rect 94668 133046 96771 133048
rect 96705 133043 96771 133046
rect 67817 132834 67883 132837
rect 226517 132834 226583 132837
rect 67817 132832 68908 132834
rect 67817 132776 67822 132832
rect 67878 132776 68908 132832
rect 224940 132832 226583 132834
rect 67817 132774 68908 132776
rect 67817 132771 67883 132774
rect 189717 132562 189783 132565
rect 193630 132562 193690 132804
rect 224940 132776 226522 132832
rect 226578 132776 226583 132832
rect 224940 132774 226583 132776
rect 226517 132771 226583 132774
rect 189717 132560 193690 132562
rect 189717 132504 189722 132560
rect 189778 132504 193690 132560
rect 189717 132502 193690 132504
rect 189717 132499 189783 132502
rect 96613 132290 96679 132293
rect 94668 132288 96679 132290
rect 94668 132232 96618 132288
rect 96674 132232 96679 132288
rect 94668 132230 96679 132232
rect 96613 132227 96679 132230
rect 94814 132092 94820 132156
rect 94884 132154 94890 132156
rect 192569 132154 192635 132157
rect 94884 132152 192635 132154
rect 94884 132096 192574 132152
rect 192630 132096 192635 132152
rect 94884 132094 192635 132096
rect 94884 132092 94890 132094
rect 192569 132091 192635 132094
rect 66253 132018 66319 132021
rect 191189 132018 191255 132021
rect 226333 132018 226399 132021
rect 66253 132016 68908 132018
rect 66253 131960 66258 132016
rect 66314 131960 68908 132016
rect 66253 131958 68908 131960
rect 191189 132016 193660 132018
rect 191189 131960 191194 132016
rect 191250 131960 193660 132016
rect 191189 131958 193660 131960
rect 224940 132016 226399 132018
rect 224940 131960 226338 132016
rect 226394 131960 226399 132016
rect 224940 131958 226399 131960
rect 66253 131955 66319 131958
rect 191189 131955 191255 131958
rect 226333 131955 226399 131958
rect 96705 131474 96771 131477
rect 94668 131472 96771 131474
rect 94668 131416 96710 131472
rect 96766 131416 96771 131472
rect 94668 131414 96771 131416
rect 96705 131411 96771 131414
rect 66345 131202 66411 131205
rect 66345 131200 68908 131202
rect 66345 131144 66350 131200
rect 66406 131144 68908 131200
rect 66345 131142 68908 131144
rect 66345 131139 66411 131142
rect 190310 131140 190316 131204
rect 190380 131202 190386 131204
rect 190380 131142 193660 131202
rect 190380 131140 190386 131142
rect 96705 130930 96771 130933
rect 225597 130930 225663 130933
rect 94668 130928 96771 130930
rect 94668 130872 96710 130928
rect 96766 130872 96771 130928
rect 94668 130870 96771 130872
rect 224940 130928 225663 130930
rect 224940 130872 225602 130928
rect 225658 130872 225663 130928
rect 224940 130870 225663 130872
rect 96705 130867 96771 130870
rect 225597 130867 225663 130870
rect 66253 130658 66319 130661
rect 66253 130656 68908 130658
rect 66253 130600 66258 130656
rect 66314 130600 68908 130656
rect 66253 130598 68908 130600
rect 66253 130595 66319 130598
rect 224902 130596 224908 130660
rect 224972 130596 224978 130660
rect 96613 130114 96679 130117
rect 94668 130112 96679 130114
rect 94668 130056 96618 130112
rect 96674 130056 96679 130112
rect 94668 130054 96679 130056
rect 96613 130051 96679 130054
rect 190821 130114 190887 130117
rect 224910 130114 224970 130596
rect 226333 130114 226399 130117
rect 190821 130112 193660 130114
rect 190821 130056 190826 130112
rect 190882 130056 193660 130112
rect 224910 130112 226399 130114
rect 224910 130084 226338 130112
rect 190821 130054 193660 130056
rect 224940 130056 226338 130084
rect 226394 130056 226399 130112
rect 224940 130054 226399 130056
rect 190821 130051 190887 130054
rect 226333 130051 226399 130054
rect 67173 129842 67239 129845
rect 67173 129840 68908 129842
rect 67173 129784 67178 129840
rect 67234 129784 68908 129840
rect 67173 129782 68908 129784
rect 67173 129779 67239 129782
rect 225045 129570 225111 129573
rect 224910 129568 225111 129570
rect 224910 129512 225050 129568
rect 225106 129512 225111 129568
rect 224910 129510 225111 129512
rect 96705 129298 96771 129301
rect 94668 129296 96771 129298
rect 94668 129240 96710 129296
rect 96766 129240 96771 129296
rect 94668 129238 96771 129240
rect 96705 129235 96771 129238
rect 191414 129236 191420 129300
rect 191484 129298 191490 129300
rect 191649 129298 191715 129301
rect 224910 129298 224970 129510
rect 225045 129507 225111 129510
rect 225321 129298 225387 129301
rect 191484 129296 193660 129298
rect 191484 129240 191654 129296
rect 191710 129240 193660 129296
rect 224910 129296 225387 129298
rect 224910 129268 225326 129296
rect 191484 129238 193660 129240
rect 224940 129240 225326 129268
rect 225382 129240 225387 129296
rect 224940 129238 225387 129240
rect 191484 129236 191490 129238
rect 191649 129235 191715 129238
rect 225321 129235 225387 129238
rect 66253 129026 66319 129029
rect 66253 129024 68908 129026
rect 66253 128968 66258 129024
rect 66314 128968 68908 129024
rect 66253 128966 68908 128968
rect 66253 128963 66319 128966
rect 69238 128420 69244 128484
rect 69308 128420 69314 128484
rect 108297 128482 108363 128485
rect 94668 128480 108363 128482
rect 94668 128424 108302 128480
rect 108358 128424 108363 128480
rect 94668 128422 108363 128424
rect 69246 128180 69306 128420
rect 108297 128419 108363 128422
rect 188889 128482 188955 128485
rect 192702 128482 192708 128484
rect 188889 128480 192708 128482
rect 188889 128424 188894 128480
rect 188950 128424 192708 128480
rect 188889 128422 192708 128424
rect 188889 128419 188955 128422
rect 192702 128420 192708 128422
rect 192772 128482 192778 128484
rect 227069 128482 227135 128485
rect 192772 128422 193660 128482
rect 224940 128480 227135 128482
rect 224940 128424 227074 128480
rect 227130 128424 227135 128480
rect 224940 128422 227135 128424
rect 192772 128420 192778 128422
rect 227069 128419 227135 128422
rect 66897 127666 66963 127669
rect 95417 127666 95483 127669
rect 66897 127664 68908 127666
rect 66897 127608 66902 127664
rect 66958 127608 68908 127664
rect 66897 127606 68908 127608
rect 94668 127664 95483 127666
rect 94668 127608 95422 127664
rect 95478 127608 95483 127664
rect 94668 127606 95483 127608
rect 66897 127603 66963 127606
rect 95417 127603 95483 127606
rect 191649 127666 191715 127669
rect 191649 127664 193660 127666
rect 191649 127608 191654 127664
rect 191710 127608 193660 127664
rect 191649 127606 193660 127608
rect 191649 127603 191715 127606
rect 226793 127394 226859 127397
rect 224940 127392 226859 127394
rect 224940 127336 226798 127392
rect 226854 127336 226859 127392
rect 224940 127334 226859 127336
rect 226793 127331 226859 127334
rect 97625 127122 97691 127125
rect 94668 127120 97691 127122
rect 94668 127064 97630 127120
rect 97686 127064 97691 127120
rect 94668 127062 97691 127064
rect 97625 127059 97691 127062
rect 66805 126850 66871 126853
rect 66805 126848 68908 126850
rect 66805 126792 66810 126848
rect 66866 126792 68908 126848
rect 66805 126790 68908 126792
rect 66805 126787 66871 126790
rect 193121 126578 193187 126581
rect 226517 126578 226583 126581
rect 193121 126576 193660 126578
rect 193121 126520 193126 126576
rect 193182 126520 193660 126576
rect 193121 126518 193660 126520
rect 224940 126576 226583 126578
rect 224940 126520 226522 126576
rect 226578 126520 226583 126576
rect 224940 126518 226583 126520
rect 193121 126515 193187 126518
rect 226517 126515 226583 126518
rect 97901 126306 97967 126309
rect 94668 126304 97967 126306
rect 94668 126248 97906 126304
rect 97962 126248 97967 126304
rect 94668 126246 97967 126248
rect 97901 126243 97967 126246
rect 66897 126034 66963 126037
rect 582925 126034 582991 126037
rect 583520 126034 584960 126124
rect 66897 126032 68908 126034
rect 66897 125976 66902 126032
rect 66958 125976 68908 126032
rect 66897 125974 68908 125976
rect 582925 126032 584960 126034
rect 582925 125976 582930 126032
rect 582986 125976 584960 126032
rect 582925 125974 584960 125976
rect 66897 125971 66963 125974
rect 582925 125971 582991 125974
rect 583520 125884 584960 125974
rect 191005 125762 191071 125765
rect 226609 125762 226675 125765
rect 191005 125760 193660 125762
rect 191005 125704 191010 125760
rect 191066 125704 193660 125760
rect 191005 125702 193660 125704
rect 224940 125760 226675 125762
rect 224940 125704 226614 125760
rect 226670 125704 226675 125760
rect 224940 125702 226675 125704
rect 191005 125699 191071 125702
rect 226609 125699 226675 125702
rect 96705 125490 96771 125493
rect 97901 125490 97967 125493
rect 94668 125488 97967 125490
rect 94668 125432 96710 125488
rect 96766 125432 97906 125488
rect 97962 125432 97967 125488
rect 94668 125430 97967 125432
rect 96705 125427 96771 125430
rect 97901 125427 97967 125430
rect 66805 125218 66871 125221
rect 66805 125216 68908 125218
rect 66805 125160 66810 125216
rect 66866 125160 68908 125216
rect 66805 125158 68908 125160
rect 66805 125155 66871 125158
rect 97809 124674 97875 124677
rect 94668 124672 97875 124674
rect 94668 124616 97814 124672
rect 97870 124616 97875 124672
rect 94668 124614 97875 124616
rect 97809 124611 97875 124614
rect 67766 124340 67772 124404
rect 67836 124402 67842 124404
rect 67836 124342 68908 124402
rect 67836 124340 67842 124342
rect 189717 124266 189783 124269
rect 193630 124266 193690 124916
rect 226793 124674 226859 124677
rect 224940 124672 226859 124674
rect 224940 124616 226798 124672
rect 226854 124616 226859 124672
rect 224940 124614 226859 124616
rect 226793 124611 226859 124614
rect 189717 124264 193690 124266
rect 189717 124208 189722 124264
rect 189778 124208 193690 124264
rect 189717 124206 193690 124208
rect 189717 124203 189783 124206
rect 97901 124130 97967 124133
rect 94668 124128 97967 124130
rect 94668 124072 97906 124128
rect 97962 124072 97967 124128
rect 94668 124070 97967 124072
rect 97901 124067 97967 124070
rect 224350 124068 224356 124132
rect 224420 124068 224426 124132
rect 66069 123858 66135 123861
rect 193029 123858 193095 123861
rect 66069 123856 68908 123858
rect -960 123572 480 123812
rect 66069 123800 66074 123856
rect 66130 123800 68908 123856
rect 66069 123798 68908 123800
rect 193029 123856 193660 123858
rect 193029 123800 193034 123856
rect 193090 123800 193660 123856
rect 224358 123828 224418 124068
rect 193029 123798 193660 123800
rect 66069 123795 66135 123798
rect 193029 123795 193095 123798
rect 97717 123450 97783 123453
rect 173341 123450 173407 123453
rect 97717 123448 173407 123450
rect 97717 123392 97722 123448
rect 97778 123392 173346 123448
rect 173402 123392 173407 123448
rect 97717 123390 173407 123392
rect 97717 123387 97783 123390
rect 173341 123387 173407 123390
rect 97441 123314 97507 123317
rect 94668 123312 97507 123314
rect 94668 123256 97446 123312
rect 97502 123256 97507 123312
rect 94668 123254 97507 123256
rect 97441 123251 97507 123254
rect 66805 123042 66871 123045
rect 226609 123042 226675 123045
rect 66805 123040 68908 123042
rect 66805 122984 66810 123040
rect 66866 122984 68908 123040
rect 224940 123040 226675 123042
rect 66805 122982 68908 122984
rect 66805 122979 66871 122982
rect 185761 122906 185827 122909
rect 193630 122906 193690 123012
rect 224940 122984 226614 123040
rect 226670 122984 226675 123040
rect 224940 122982 226675 122984
rect 226609 122979 226675 122982
rect 185761 122904 193690 122906
rect 185761 122848 185766 122904
rect 185822 122848 193690 122904
rect 185761 122846 193690 122848
rect 185761 122843 185827 122846
rect 97901 122498 97967 122501
rect 94668 122496 97967 122498
rect 94668 122440 97906 122496
rect 97962 122440 97967 122496
rect 94668 122438 97967 122440
rect 97901 122435 97967 122438
rect 66345 122226 66411 122229
rect 191557 122226 191623 122229
rect 226609 122226 226675 122229
rect 66345 122224 68908 122226
rect 66345 122168 66350 122224
rect 66406 122168 68908 122224
rect 66345 122166 68908 122168
rect 191557 122224 193660 122226
rect 191557 122168 191562 122224
rect 191618 122168 193660 122224
rect 191557 122166 193660 122168
rect 224940 122224 226675 122226
rect 224940 122168 226614 122224
rect 226670 122168 226675 122224
rect 224940 122166 226675 122168
rect 66345 122163 66411 122166
rect 191557 122163 191623 122166
rect 226609 122163 226675 122166
rect 97441 121682 97507 121685
rect 94668 121680 97507 121682
rect 94668 121624 97446 121680
rect 97502 121624 97507 121680
rect 94668 121622 97507 121624
rect 97441 121619 97507 121622
rect 66805 121410 66871 121413
rect 190821 121410 190887 121413
rect 66805 121408 68908 121410
rect 66805 121352 66810 121408
rect 66866 121352 68908 121408
rect 66805 121350 68908 121352
rect 190821 121408 193660 121410
rect 190821 121352 190826 121408
rect 190882 121352 193660 121408
rect 190821 121350 193660 121352
rect 66805 121347 66871 121350
rect 190821 121347 190887 121350
rect 97625 120866 97691 120869
rect 94668 120864 97691 120866
rect 94668 120808 97630 120864
rect 97686 120808 97691 120864
rect 94668 120806 97691 120808
rect 97625 120803 97691 120806
rect 66897 120594 66963 120597
rect 224910 120594 224970 121108
rect 66897 120592 68908 120594
rect 66897 120536 66902 120592
rect 66958 120536 68908 120592
rect 66897 120534 68908 120536
rect 224910 120534 229110 120594
rect 66897 120531 66963 120534
rect 95325 120322 95391 120325
rect 97533 120322 97599 120325
rect 94668 120320 97599 120322
rect 94668 120264 95330 120320
rect 95386 120264 97538 120320
rect 97594 120264 97599 120320
rect 94668 120262 97599 120264
rect 95325 120259 95391 120262
rect 97533 120259 97599 120262
rect 190453 120322 190519 120325
rect 226609 120322 226675 120325
rect 190453 120320 193660 120322
rect 190453 120264 190458 120320
rect 190514 120264 193660 120320
rect 190453 120262 193660 120264
rect 224940 120320 226675 120322
rect 224940 120264 226614 120320
rect 226670 120264 226675 120320
rect 224940 120262 226675 120264
rect 229050 120322 229110 120534
rect 240225 120322 240291 120325
rect 229050 120320 240291 120322
rect 229050 120264 240230 120320
rect 240286 120264 240291 120320
rect 229050 120262 240291 120264
rect 190453 120259 190519 120262
rect 226609 120259 226675 120262
rect 240225 120259 240291 120262
rect 66805 120050 66871 120053
rect 66805 120048 68908 120050
rect 66805 119992 66810 120048
rect 66866 119992 68908 120048
rect 66805 119990 68908 119992
rect 66805 119987 66871 119990
rect 96286 119988 96292 120052
rect 96356 120050 96362 120052
rect 182357 120050 182423 120053
rect 183001 120050 183067 120053
rect 96356 120048 183067 120050
rect 96356 119992 182362 120048
rect 182418 119992 183006 120048
rect 183062 119992 183067 120048
rect 96356 119990 183067 119992
rect 96356 119988 96362 119990
rect 182357 119987 182423 119990
rect 183001 119987 183067 119990
rect 97165 119506 97231 119509
rect 94668 119504 97231 119506
rect 94668 119448 97170 119504
rect 97226 119448 97231 119504
rect 94668 119446 97231 119448
rect 97165 119443 97231 119446
rect 191557 119506 191623 119509
rect 226609 119506 226675 119509
rect 191557 119504 193660 119506
rect 191557 119448 191562 119504
rect 191618 119448 193660 119504
rect 191557 119446 193660 119448
rect 224940 119504 226675 119506
rect 224940 119448 226614 119504
rect 226670 119448 226675 119504
rect 224940 119446 226675 119448
rect 191557 119443 191623 119446
rect 226609 119443 226675 119446
rect 66897 119234 66963 119237
rect 66897 119232 68908 119234
rect 66897 119176 66902 119232
rect 66958 119176 68908 119232
rect 66897 119174 68908 119176
rect 66897 119171 66963 119174
rect 97901 118690 97967 118693
rect 94668 118688 97967 118690
rect 94668 118632 97906 118688
rect 97962 118632 97967 118688
rect 94668 118630 97967 118632
rect 97901 118627 97967 118630
rect 191557 118690 191623 118693
rect 191557 118688 193660 118690
rect 191557 118632 191562 118688
rect 191618 118632 193660 118688
rect 191557 118630 193660 118632
rect 191557 118627 191623 118630
rect 66897 118418 66963 118421
rect 226793 118418 226859 118421
rect 66897 118416 68908 118418
rect 66897 118360 66902 118416
rect 66958 118360 68908 118416
rect 66897 118358 68908 118360
rect 224940 118416 226859 118418
rect 224940 118360 226798 118416
rect 226854 118360 226859 118416
rect 224940 118358 226859 118360
rect 66897 118355 66963 118358
rect 226793 118355 226859 118358
rect 190821 118010 190887 118013
rect 191598 118010 191604 118012
rect 190821 118008 191604 118010
rect 190821 117952 190826 118008
rect 190882 117952 191604 118008
rect 190821 117950 191604 117952
rect 190821 117947 190887 117950
rect 191598 117948 191604 117950
rect 191668 118010 191674 118012
rect 191668 117950 193690 118010
rect 191668 117948 191674 117950
rect 97809 117874 97875 117877
rect 94668 117872 97875 117874
rect 94668 117816 97814 117872
rect 97870 117816 97875 117872
rect 94668 117814 97875 117816
rect 97809 117811 97875 117814
rect 66805 117602 66871 117605
rect 66805 117600 68908 117602
rect 66805 117544 66810 117600
rect 66866 117544 68908 117600
rect 193630 117572 193690 117950
rect 226609 117602 226675 117605
rect 224940 117600 226675 117602
rect 66805 117542 68908 117544
rect 224940 117544 226614 117600
rect 226670 117544 226675 117600
rect 224940 117542 226675 117544
rect 66805 117539 66871 117542
rect 226609 117539 226675 117542
rect 66110 116996 66116 117060
rect 66180 117058 66186 117060
rect 97901 117058 97967 117061
rect 66180 116998 68908 117058
rect 94668 117056 97967 117058
rect 94668 117000 97906 117056
rect 97962 117000 97967 117056
rect 94668 116998 97967 117000
rect 66180 116996 66186 116998
rect 97901 116995 97967 116998
rect 191557 116786 191623 116789
rect 225229 116786 225295 116789
rect 191557 116784 193660 116786
rect 191557 116728 191562 116784
rect 191618 116728 193660 116784
rect 191557 116726 193660 116728
rect 224940 116784 225295 116786
rect 224940 116728 225234 116784
rect 225290 116728 225295 116784
rect 224940 116726 225295 116728
rect 191557 116723 191623 116726
rect 225229 116723 225295 116726
rect 97349 116650 97415 116653
rect 100886 116650 100892 116652
rect 97349 116648 100892 116650
rect 97349 116592 97354 116648
rect 97410 116592 100892 116648
rect 97349 116590 100892 116592
rect 97349 116587 97415 116590
rect 100886 116588 100892 116590
rect 100956 116588 100962 116652
rect 97717 116514 97783 116517
rect 94668 116512 97783 116514
rect 94668 116456 97722 116512
rect 97778 116456 97783 116512
rect 94668 116454 97783 116456
rect 97717 116451 97783 116454
rect 66621 116242 66687 116245
rect 66621 116240 68908 116242
rect 66621 116184 66626 116240
rect 66682 116184 68908 116240
rect 66621 116182 68908 116184
rect 66621 116179 66687 116182
rect 191373 115970 191439 115973
rect 226609 115970 226675 115973
rect 191373 115968 193660 115970
rect 191373 115912 191378 115968
rect 191434 115912 193660 115968
rect 191373 115910 193660 115912
rect 224940 115968 226675 115970
rect 224940 115912 226614 115968
rect 226670 115912 226675 115968
rect 224940 115910 226675 115912
rect 191373 115907 191439 115910
rect 226609 115907 226675 115910
rect 97165 115698 97231 115701
rect 94668 115696 97231 115698
rect 94668 115640 97170 115696
rect 97226 115640 97231 115696
rect 94668 115638 97231 115640
rect 97165 115635 97231 115638
rect 66805 115426 66871 115429
rect 66805 115424 68908 115426
rect 66805 115368 66810 115424
rect 66866 115368 68908 115424
rect 66805 115366 68908 115368
rect 66805 115363 66871 115366
rect 191005 115154 191071 115157
rect 191005 115152 193660 115154
rect 191005 115096 191010 115152
rect 191066 115096 193660 115152
rect 191005 115094 193660 115096
rect 191005 115091 191071 115094
rect 97533 114882 97599 114885
rect 227989 114882 228055 114885
rect 94668 114880 97599 114882
rect 94668 114824 97538 114880
rect 97594 114824 97599 114880
rect 94668 114822 97599 114824
rect 224940 114880 228055 114882
rect 224940 114824 227994 114880
rect 228050 114824 228055 114880
rect 224940 114822 228055 114824
rect 97533 114819 97599 114822
rect 227989 114819 228055 114822
rect 66897 114610 66963 114613
rect 66897 114608 68908 114610
rect 66897 114552 66902 114608
rect 66958 114552 68908 114608
rect 66897 114550 68908 114552
rect 66897 114547 66963 114550
rect 97349 114066 97415 114069
rect 94668 114064 97415 114066
rect 94668 114008 97354 114064
rect 97410 114008 97415 114064
rect 94668 114006 97415 114008
rect 97349 114003 97415 114006
rect 190821 114066 190887 114069
rect 227805 114066 227871 114069
rect 190821 114064 193660 114066
rect 190821 114008 190826 114064
rect 190882 114008 193660 114064
rect 190821 114006 193660 114008
rect 224940 114064 227871 114066
rect 224940 114008 227810 114064
rect 227866 114008 227871 114064
rect 224940 114006 227871 114008
rect 190821 114003 190887 114006
rect 227805 114003 227871 114006
rect 66805 113794 66871 113797
rect 66805 113792 68908 113794
rect 66805 113736 66810 113792
rect 66866 113736 68908 113792
rect 66805 113734 68908 113736
rect 66805 113731 66871 113734
rect 97533 113522 97599 113525
rect 94668 113520 97599 113522
rect 94668 113464 97538 113520
rect 97594 113464 97599 113520
rect 94668 113462 97599 113464
rect 97533 113459 97599 113462
rect 66897 113250 66963 113253
rect 191557 113250 191623 113253
rect 226517 113250 226583 113253
rect 66897 113248 68908 113250
rect 66897 113192 66902 113248
rect 66958 113192 68908 113248
rect 66897 113190 68908 113192
rect 191557 113248 193660 113250
rect 191557 113192 191562 113248
rect 191618 113192 193660 113248
rect 191557 113190 193660 113192
rect 224940 113248 226583 113250
rect 224940 113192 226522 113248
rect 226578 113192 226583 113248
rect 224940 113190 226583 113192
rect 66897 113187 66963 113190
rect 191557 113187 191623 113190
rect 226517 113187 226583 113190
rect 582649 112842 582715 112845
rect 583520 112842 584960 112932
rect 582649 112840 584960 112842
rect 582649 112784 582654 112840
rect 582710 112784 584960 112840
rect 582649 112782 584960 112784
rect 582649 112779 582715 112782
rect 97901 112706 97967 112709
rect 94668 112704 97967 112706
rect 94668 112648 97906 112704
rect 97962 112648 97967 112704
rect 583520 112692 584960 112782
rect 94668 112646 97967 112648
rect 97901 112643 97967 112646
rect 67725 112434 67791 112437
rect 191557 112434 191623 112437
rect 67725 112432 68908 112434
rect 67725 112376 67730 112432
rect 67786 112376 68908 112432
rect 67725 112374 68908 112376
rect 191557 112432 193660 112434
rect 191557 112376 191562 112432
rect 191618 112376 193660 112432
rect 191557 112374 193660 112376
rect 67725 112371 67791 112374
rect 191557 112371 191623 112374
rect 226609 112162 226675 112165
rect 224940 112160 226675 112162
rect 224940 112104 226614 112160
rect 226670 112104 226675 112160
rect 224940 112102 226675 112104
rect 226609 112099 226675 112102
rect 96705 111890 96771 111893
rect 94668 111888 96771 111890
rect 94668 111832 96710 111888
rect 96766 111832 96771 111888
rect 94668 111830 96771 111832
rect 96705 111827 96771 111830
rect 66897 111618 66963 111621
rect 66897 111616 68908 111618
rect 66897 111560 66902 111616
rect 66958 111560 68908 111616
rect 66897 111558 68908 111560
rect 66897 111555 66963 111558
rect 226977 111346 227043 111349
rect 224940 111344 227043 111346
rect 96705 111074 96771 111077
rect 94668 111072 96771 111074
rect 94668 111016 96710 111072
rect 96766 111016 96771 111072
rect 94668 111014 96771 111016
rect 96705 111011 96771 111014
rect 67173 110802 67239 110805
rect 67725 110802 67791 110805
rect 190269 110802 190335 110805
rect 193630 110802 193690 111316
rect 224940 111288 226982 111344
rect 227038 111288 227043 111344
rect 224940 111286 227043 111288
rect 226977 111283 227043 111286
rect 67173 110800 68908 110802
rect -960 110666 480 110756
rect 67173 110744 67178 110800
rect 67234 110744 67730 110800
rect 67786 110744 68908 110800
rect 67173 110742 68908 110744
rect 190269 110800 193690 110802
rect 190269 110744 190274 110800
rect 190330 110744 193690 110800
rect 190269 110742 193690 110744
rect 67173 110739 67239 110742
rect 67725 110739 67791 110742
rect 190269 110739 190335 110742
rect 3417 110666 3483 110669
rect -960 110664 3483 110666
rect -960 110608 3422 110664
rect 3478 110608 3483 110664
rect -960 110606 3483 110608
rect -960 110516 480 110606
rect 3417 110603 3483 110606
rect 191189 110530 191255 110533
rect 226701 110530 226767 110533
rect 191189 110528 193660 110530
rect 191189 110472 191194 110528
rect 191250 110472 193660 110528
rect 191189 110470 193660 110472
rect 224940 110528 226767 110530
rect 224940 110472 226706 110528
rect 226762 110472 226767 110528
rect 224940 110470 226767 110472
rect 191189 110467 191255 110470
rect 226701 110467 226767 110470
rect 65977 110258 66043 110261
rect 97073 110258 97139 110261
rect 65977 110256 68908 110258
rect 65977 110200 65982 110256
rect 66038 110200 68908 110256
rect 65977 110198 68908 110200
rect 94668 110256 97139 110258
rect 94668 110200 97078 110256
rect 97134 110200 97139 110256
rect 94668 110198 97139 110200
rect 65977 110195 66043 110198
rect 97073 110195 97139 110198
rect 97901 109714 97967 109717
rect 94668 109712 97967 109714
rect 94668 109656 97906 109712
rect 97962 109656 97967 109712
rect 94668 109654 97967 109656
rect 97901 109651 97967 109654
rect 191005 109714 191071 109717
rect 226425 109714 226491 109717
rect 191005 109712 193660 109714
rect 191005 109656 191010 109712
rect 191066 109656 193660 109712
rect 191005 109654 193660 109656
rect 224940 109712 226491 109714
rect 224940 109656 226430 109712
rect 226486 109656 226491 109712
rect 224940 109654 226491 109656
rect 191005 109651 191071 109654
rect 226425 109651 226491 109654
rect 66805 109442 66871 109445
rect 66805 109440 68908 109442
rect 66805 109384 66810 109440
rect 66866 109384 68908 109440
rect 66805 109382 68908 109384
rect 66805 109379 66871 109382
rect 94638 108762 94698 108868
rect 94773 108762 94839 108765
rect 94638 108760 94839 108762
rect 94638 108704 94778 108760
rect 94834 108704 94839 108760
rect 94638 108702 94839 108704
rect 94773 108699 94839 108702
rect 66478 108564 66484 108628
rect 66548 108626 66554 108628
rect 66548 108566 68908 108626
rect 66548 108564 66554 108566
rect 98494 108292 98500 108356
rect 98564 108354 98570 108356
rect 111885 108354 111951 108357
rect 98564 108352 111951 108354
rect 98564 108296 111890 108352
rect 111946 108296 111951 108352
rect 98564 108294 111951 108296
rect 98564 108292 98570 108294
rect 111885 108291 111951 108294
rect 97942 108082 97948 108084
rect 94668 108022 97948 108082
rect 97942 108020 97948 108022
rect 98012 108020 98018 108084
rect 184054 108020 184060 108084
rect 184124 108082 184130 108084
rect 193630 108082 193690 108868
rect 226609 108628 226675 108629
rect 226558 108626 226564 108628
rect 224940 108566 226564 108626
rect 226628 108624 226675 108628
rect 226670 108568 226675 108624
rect 226558 108564 226564 108566
rect 226628 108564 226675 108568
rect 226609 108563 226675 108564
rect 184124 108022 193690 108082
rect 184124 108020 184130 108022
rect 65885 107810 65951 107813
rect 226374 107810 226380 107812
rect 65885 107808 68908 107810
rect 65885 107752 65890 107808
rect 65946 107752 68908 107808
rect 65885 107750 68908 107752
rect 65885 107747 65951 107750
rect 193630 107674 193690 107780
rect 224940 107750 226380 107810
rect 226374 107748 226380 107750
rect 226444 107748 226450 107812
rect 190410 107614 193690 107674
rect 187550 107476 187556 107540
rect 187620 107538 187626 107540
rect 190410 107538 190470 107614
rect 187620 107478 190470 107538
rect 187620 107476 187626 107478
rect 97901 107266 97967 107269
rect 94668 107264 97967 107266
rect 94668 107208 97906 107264
rect 97962 107208 97967 107264
rect 94668 107206 97967 107208
rect 97901 107203 97967 107206
rect 66662 106932 66668 106996
rect 66732 106994 66738 106996
rect 66805 106994 66871 106997
rect 190637 106994 190703 106997
rect 226701 106994 226767 106997
rect 66732 106992 68908 106994
rect 66732 106936 66810 106992
rect 66866 106936 68908 106992
rect 66732 106934 68908 106936
rect 190637 106992 193660 106994
rect 190637 106936 190642 106992
rect 190698 106936 193660 106992
rect 190637 106934 193660 106936
rect 224940 106992 226767 106994
rect 224940 106936 226706 106992
rect 226762 106936 226767 106992
rect 224940 106934 226767 106936
rect 66732 106932 66738 106934
rect 66805 106931 66871 106934
rect 190637 106931 190703 106934
rect 226701 106931 226767 106934
rect 61878 106252 61884 106316
rect 61948 106314 61954 106316
rect 68878 106314 68938 106420
rect 61948 106254 68938 106314
rect 94638 106314 94698 106692
rect 162209 106314 162275 106317
rect 94638 106312 162275 106314
rect 94638 106256 162214 106312
rect 162270 106256 162275 106312
rect 94638 106254 162275 106256
rect 61948 106252 61954 106254
rect 162209 106251 162275 106254
rect 191005 106178 191071 106181
rect 191005 106176 193660 106178
rect 191005 106120 191010 106176
rect 191066 106120 193660 106176
rect 191005 106118 193660 106120
rect 191005 106115 191071 106118
rect 100702 105906 100708 105908
rect 94668 105846 100708 105906
rect 100702 105844 100708 105846
rect 100772 105844 100778 105908
rect 226701 105906 226767 105909
rect 224940 105904 226767 105906
rect 224940 105848 226706 105904
rect 226762 105848 226767 105904
rect 224940 105846 226767 105848
rect 226701 105843 226767 105846
rect 66621 105634 66687 105637
rect 66621 105632 68908 105634
rect 66621 105576 66626 105632
rect 66682 105576 68908 105632
rect 66621 105574 68908 105576
rect 66621 105571 66687 105574
rect 96797 105090 96863 105093
rect 94668 105088 96863 105090
rect 94668 105032 96802 105088
rect 96858 105032 96863 105088
rect 94668 105030 96863 105032
rect 96797 105027 96863 105030
rect 191557 105090 191623 105093
rect 191557 105088 193660 105090
rect 191557 105032 191562 105088
rect 191618 105032 193660 105088
rect 191557 105030 193660 105032
rect 191557 105027 191623 105030
rect 224910 104954 224970 105060
rect 225045 104954 225111 104957
rect 224910 104952 225111 104954
rect 224910 104896 225050 104952
rect 225106 104896 225111 104952
rect 224910 104894 225111 104896
rect 225045 104891 225111 104894
rect 66805 104818 66871 104821
rect 66805 104816 68908 104818
rect 66805 104760 66810 104816
rect 66866 104760 68908 104816
rect 66805 104758 68908 104760
rect 66805 104755 66871 104758
rect 97901 104274 97967 104277
rect 94668 104272 97967 104274
rect 94668 104216 97906 104272
rect 97962 104216 97967 104272
rect 94668 104214 97967 104216
rect 97901 104211 97967 104214
rect 193213 104274 193279 104277
rect 226517 104274 226583 104277
rect 193213 104272 193660 104274
rect 193213 104216 193218 104272
rect 193274 104216 193660 104272
rect 193213 104214 193660 104216
rect 224940 104272 226583 104274
rect 224940 104216 226522 104272
rect 226578 104216 226583 104272
rect 224940 104214 226583 104216
rect 193213 104211 193279 104214
rect 226517 104211 226583 104214
rect 94814 104076 94820 104140
rect 94884 104138 94890 104140
rect 121545 104138 121611 104141
rect 94884 104136 121611 104138
rect 94884 104080 121550 104136
rect 121606 104080 121611 104136
rect 94884 104078 121611 104080
rect 94884 104076 94890 104078
rect 121545 104075 121611 104078
rect 67265 104002 67331 104005
rect 67265 104000 68908 104002
rect 67265 103944 67270 104000
rect 67326 103944 68908 104000
rect 67265 103942 68908 103944
rect 67265 103939 67331 103942
rect 97809 103458 97875 103461
rect 94668 103456 97875 103458
rect 94668 103400 97814 103456
rect 97870 103400 97875 103456
rect 94668 103398 97875 103400
rect 97809 103395 97875 103398
rect 191557 103458 191623 103461
rect 226609 103458 226675 103461
rect 191557 103456 193660 103458
rect 191557 103400 191562 103456
rect 191618 103400 193660 103456
rect 191557 103398 193660 103400
rect 224940 103456 226675 103458
rect 224940 103400 226614 103456
rect 226670 103400 226675 103456
rect 224940 103398 226675 103400
rect 191557 103395 191623 103398
rect 226609 103395 226675 103398
rect 67817 103186 67883 103189
rect 67817 103184 68908 103186
rect 67817 103128 67822 103184
rect 67878 103128 68908 103184
rect 67817 103126 68908 103128
rect 67817 103123 67883 103126
rect 97901 102914 97967 102917
rect 94668 102912 97967 102914
rect 94668 102856 97906 102912
rect 97962 102856 97967 102912
rect 94668 102854 97967 102856
rect 97901 102851 97967 102854
rect 66805 102642 66871 102645
rect 191465 102642 191531 102645
rect 66805 102640 68908 102642
rect 66805 102584 66810 102640
rect 66866 102584 68908 102640
rect 66805 102582 68908 102584
rect 191465 102640 193660 102642
rect 191465 102584 191470 102640
rect 191526 102584 193660 102640
rect 191465 102582 193660 102584
rect 66805 102579 66871 102582
rect 191465 102579 191531 102582
rect 227897 102370 227963 102373
rect 224940 102368 227963 102370
rect 224940 102312 227902 102368
rect 227958 102312 227963 102368
rect 224940 102310 227963 102312
rect 227897 102307 227963 102310
rect 96705 102098 96771 102101
rect 94668 102096 96771 102098
rect 94668 102040 96710 102096
rect 96766 102040 96771 102096
rect 94668 102038 96771 102040
rect 96705 102035 96771 102038
rect 66529 101826 66595 101829
rect 66529 101824 68908 101826
rect 66529 101768 66534 101824
rect 66590 101768 68908 101824
rect 66529 101766 68908 101768
rect 66529 101763 66595 101766
rect 190637 101554 190703 101557
rect 227437 101554 227503 101557
rect 190637 101552 193660 101554
rect 190637 101496 190642 101552
rect 190698 101496 193660 101552
rect 190637 101494 193660 101496
rect 224940 101552 227503 101554
rect 224940 101496 227442 101552
rect 227498 101496 227503 101552
rect 224940 101494 227503 101496
rect 190637 101491 190703 101494
rect 227437 101491 227503 101494
rect 96705 101282 96771 101285
rect 94668 101280 96771 101282
rect 94668 101224 96710 101280
rect 96766 101224 96771 101280
rect 94668 101222 96771 101224
rect 96705 101219 96771 101222
rect 66805 101010 66871 101013
rect 66805 101008 68908 101010
rect 66805 100952 66810 101008
rect 66866 100952 68908 101008
rect 66805 100950 68908 100952
rect 66805 100947 66871 100950
rect 191741 100874 191807 100877
rect 191741 100872 191850 100874
rect 191741 100816 191746 100872
rect 191802 100816 191850 100872
rect 191741 100811 191850 100816
rect 191557 100738 191623 100741
rect 191790 100738 191850 100811
rect 225137 100738 225203 100741
rect 191557 100736 193660 100738
rect 191557 100680 191562 100736
rect 191618 100680 193660 100736
rect 191557 100678 193660 100680
rect 224940 100736 225203 100738
rect 224940 100680 225142 100736
rect 225198 100680 225203 100736
rect 224940 100678 225203 100680
rect 191557 100675 191623 100678
rect 225137 100675 225203 100678
rect 97441 100466 97507 100469
rect 94668 100464 97507 100466
rect 94668 100408 97446 100464
rect 97502 100408 97507 100464
rect 94668 100406 97507 100408
rect 97441 100403 97507 100406
rect 66713 100194 66779 100197
rect 66713 100192 68908 100194
rect 66713 100136 66718 100192
rect 66774 100136 68908 100192
rect 66713 100134 68908 100136
rect 66713 100131 66779 100134
rect 191741 99922 191807 99925
rect 191741 99920 193660 99922
rect 191741 99864 191746 99920
rect 191802 99864 193660 99920
rect 191741 99862 193660 99864
rect 191741 99859 191807 99862
rect 66253 99650 66319 99653
rect 97901 99650 97967 99653
rect 226425 99650 226491 99653
rect 66253 99648 68908 99650
rect 66253 99592 66258 99648
rect 66314 99592 68908 99648
rect 66253 99590 68908 99592
rect 94668 99648 97967 99650
rect 94668 99592 97906 99648
rect 97962 99592 97967 99648
rect 94668 99590 97967 99592
rect 224940 99648 226491 99650
rect 224940 99592 226430 99648
rect 226486 99592 226491 99648
rect 224940 99590 226491 99592
rect 66253 99587 66319 99590
rect 97901 99587 97967 99590
rect 226425 99587 226491 99590
rect 582649 99514 582715 99517
rect 583520 99514 584960 99604
rect 582649 99512 584960 99514
rect 582649 99456 582654 99512
rect 582710 99456 584960 99512
rect 582649 99454 584960 99456
rect 582649 99451 582715 99454
rect 583520 99364 584960 99454
rect 97901 99106 97967 99109
rect 94668 99104 97967 99106
rect 94668 99048 97906 99104
rect 97962 99048 97967 99104
rect 94668 99046 97967 99048
rect 97901 99043 97967 99046
rect 226425 98834 226491 98837
rect 224940 98832 226491 98834
rect 68878 98290 68938 98804
rect 100753 98698 100819 98701
rect 107745 98698 107811 98701
rect 108297 98698 108363 98701
rect 100753 98696 108363 98698
rect 100753 98640 100758 98696
rect 100814 98640 107750 98696
rect 107806 98640 108302 98696
rect 108358 98640 108363 98696
rect 100753 98638 108363 98640
rect 100753 98635 100819 98638
rect 107745 98635 107811 98638
rect 108297 98635 108363 98638
rect 96521 98290 96587 98293
rect 97901 98290 97967 98293
rect 64830 98230 68938 98290
rect 94668 98288 97967 98290
rect 94668 98232 96526 98288
rect 96582 98232 97906 98288
rect 97962 98232 97967 98288
rect 94668 98230 97967 98232
rect 57830 98092 57836 98156
rect 57900 98154 57906 98156
rect 64830 98154 64890 98230
rect 96521 98227 96587 98230
rect 97901 98227 97967 98230
rect 189901 98290 189967 98293
rect 193630 98290 193690 98804
rect 224940 98776 226430 98832
rect 226486 98776 226491 98832
rect 224940 98774 226491 98776
rect 226425 98771 226491 98774
rect 189901 98288 193690 98290
rect 189901 98232 189906 98288
rect 189962 98232 193690 98288
rect 189901 98230 193690 98232
rect 189901 98227 189967 98230
rect 57900 98094 64890 98154
rect 57900 98092 57906 98094
rect 67449 98018 67515 98021
rect 191741 98018 191807 98021
rect 226701 98018 226767 98021
rect 67449 98016 68908 98018
rect 67449 97960 67454 98016
rect 67510 97960 68908 98016
rect 67449 97958 68908 97960
rect 191741 98016 193660 98018
rect 191741 97960 191746 98016
rect 191802 97960 193660 98016
rect 191741 97958 193660 97960
rect 224940 98016 226767 98018
rect 224940 97960 226706 98016
rect 226762 97960 226767 98016
rect 224940 97958 226767 97960
rect 67449 97955 67515 97958
rect 191741 97955 191807 97958
rect 226701 97955 226767 97958
rect -960 97610 480 97700
rect 3417 97610 3483 97613
rect -960 97608 3483 97610
rect -960 97552 3422 97608
rect 3478 97552 3483 97608
rect -960 97550 3483 97552
rect -960 97460 480 97550
rect 3417 97547 3483 97550
rect 67357 97202 67423 97205
rect 67357 97200 68908 97202
rect 67357 97144 67362 97200
rect 67418 97144 68908 97200
rect 67357 97142 68908 97144
rect 67357 97139 67423 97142
rect 94638 96930 94698 97444
rect 224718 97412 224724 97476
rect 224788 97474 224794 97476
rect 270585 97474 270651 97477
rect 224788 97472 270651 97474
rect 224788 97416 270590 97472
rect 270646 97416 270651 97472
rect 224788 97414 270651 97416
rect 224788 97412 224794 97414
rect 270585 97411 270651 97414
rect 190637 97202 190703 97205
rect 226517 97202 226583 97205
rect 190637 97200 193660 97202
rect 190637 97144 190642 97200
rect 190698 97144 193660 97200
rect 190637 97142 193660 97144
rect 224940 97200 226583 97202
rect 224940 97144 226522 97200
rect 226578 97144 226583 97200
rect 224940 97142 226583 97144
rect 190637 97139 190703 97142
rect 226517 97139 226583 97142
rect 191046 96930 191052 96932
rect 94638 96870 191052 96930
rect 191046 96868 191052 96870
rect 191116 96868 191122 96932
rect 96705 96658 96771 96661
rect 94668 96656 96771 96658
rect 94668 96600 96710 96656
rect 96766 96600 96771 96656
rect 94668 96598 96771 96600
rect 96705 96595 96771 96598
rect 193029 96386 193095 96389
rect 193029 96384 193660 96386
rect 68878 96114 68938 96356
rect 193029 96328 193034 96384
rect 193090 96328 193660 96384
rect 193029 96326 193660 96328
rect 193029 96323 193095 96326
rect 97809 96114 97875 96117
rect 226977 96114 227043 96117
rect 64830 96054 68938 96114
rect 94668 96112 97875 96114
rect 94668 96056 97814 96112
rect 97870 96056 97875 96112
rect 94668 96054 97875 96056
rect 224940 96112 227043 96114
rect 224940 96056 226982 96112
rect 227038 96056 227043 96112
rect 224940 96054 227043 96056
rect 64638 95372 64644 95436
rect 64708 95434 64714 95436
rect 64830 95434 64890 96054
rect 97809 96051 97875 96054
rect 226977 96051 227043 96054
rect 66897 95842 66963 95845
rect 66897 95840 68908 95842
rect 66897 95784 66902 95840
rect 66958 95784 68908 95840
rect 66897 95782 68908 95784
rect 66897 95779 66963 95782
rect 64708 95374 64890 95434
rect 64708 95372 64714 95374
rect 97901 95298 97967 95301
rect 94668 95296 97967 95298
rect 94668 95240 97906 95296
rect 97962 95240 97967 95296
rect 94668 95238 97967 95240
rect 97901 95235 97967 95238
rect 173249 95298 173315 95301
rect 226333 95298 226399 95301
rect 173249 95296 193660 95298
rect 173249 95240 173254 95296
rect 173310 95240 193660 95296
rect 224940 95296 226399 95298
rect 224940 95268 226338 95296
rect 173249 95238 193660 95240
rect 224910 95240 226338 95268
rect 226394 95240 226399 95296
rect 224910 95238 226399 95240
rect 173249 95235 173315 95238
rect 224910 95164 224970 95238
rect 226333 95235 226399 95238
rect 224902 95100 224908 95164
rect 224972 95100 224978 95164
rect 66805 95026 66871 95029
rect 97257 95026 97323 95029
rect 66805 95024 68908 95026
rect 66805 94968 66810 95024
rect 66866 94968 68908 95024
rect 66805 94966 68908 94968
rect 94638 95024 97323 95026
rect 94638 94968 97262 95024
rect 97318 94968 97323 95024
rect 94638 94966 97323 94968
rect 66805 94963 66871 94966
rect 94638 94452 94698 94966
rect 97257 94963 97323 94966
rect 153101 94754 153167 94757
rect 193438 94754 193444 94756
rect 142110 94752 193444 94754
rect 142110 94696 153106 94752
rect 153162 94696 193444 94752
rect 142110 94694 193444 94696
rect 96981 94482 97047 94485
rect 142110 94482 142170 94694
rect 153101 94691 153167 94694
rect 193438 94692 193444 94694
rect 193508 94692 193514 94756
rect 224350 94692 224356 94756
rect 224420 94754 224426 94756
rect 262213 94754 262279 94757
rect 224420 94752 262279 94754
rect 224420 94696 262218 94752
rect 262274 94696 262279 94752
rect 224420 94694 262279 94696
rect 224420 94692 224426 94694
rect 262213 94691 262279 94694
rect 226793 94482 226859 94485
rect 96981 94480 142170 94482
rect 96981 94424 96986 94480
rect 97042 94424 142170 94480
rect 224940 94480 226859 94482
rect 96981 94422 142170 94424
rect 96981 94419 97047 94422
rect 67265 94210 67331 94213
rect 193814 94212 193874 94452
rect 224940 94424 226798 94480
rect 226854 94424 226859 94480
rect 224940 94422 226859 94424
rect 226793 94419 226859 94422
rect 67265 94208 68908 94210
rect 67265 94152 67270 94208
rect 67326 94152 68908 94208
rect 67265 94150 68908 94152
rect 67265 94147 67331 94150
rect 193806 94148 193812 94212
rect 193876 94148 193882 94212
rect 97901 93666 97967 93669
rect 226885 93666 226951 93669
rect 94668 93664 97967 93666
rect 94668 93608 97906 93664
rect 97962 93608 97967 93664
rect 224940 93664 226951 93666
rect 94668 93606 97967 93608
rect 97901 93603 97967 93606
rect 68878 92850 68938 93364
rect 94773 93122 94839 93125
rect 155309 93122 155375 93125
rect 94773 93120 155375 93122
rect 94773 93064 94778 93120
rect 94834 93064 155314 93120
rect 155370 93064 155375 93120
rect 94773 93062 155375 93064
rect 94773 93059 94839 93062
rect 155309 93059 155375 93062
rect 155493 93122 155559 93125
rect 188521 93122 188587 93125
rect 155493 93120 188587 93122
rect 155493 93064 155498 93120
rect 155554 93064 188526 93120
rect 188582 93064 188587 93120
rect 155493 93062 188587 93064
rect 155493 93059 155559 93062
rect 188521 93059 188587 93062
rect 194182 92986 194242 93636
rect 224940 93608 226890 93664
rect 226946 93608 226951 93664
rect 224940 93606 226951 93608
rect 226885 93603 226951 93606
rect 211705 93396 211771 93397
rect 224769 93396 224835 93397
rect 211654 93332 211660 93396
rect 211724 93394 211771 93396
rect 211724 93392 211816 93394
rect 211766 93336 211816 93392
rect 211724 93334 211816 93336
rect 211724 93332 211771 93334
rect 224718 93332 224724 93396
rect 224788 93394 224835 93396
rect 224788 93392 224880 93394
rect 224830 93336 224880 93392
rect 224788 93334 224880 93336
rect 224788 93332 224835 93334
rect 211705 93331 211771 93332
rect 224769 93331 224835 93332
rect 222653 92986 222719 92989
rect 223430 92986 223436 92988
rect 194182 92926 194426 92986
rect 97206 92850 97212 92852
rect 68694 92790 68938 92850
rect 94668 92790 97212 92850
rect 67541 92578 67607 92581
rect 68694 92578 68754 92790
rect 97206 92788 97212 92790
rect 97276 92788 97282 92852
rect 68870 92652 68876 92716
rect 68940 92714 68946 92716
rect 69703 92714 69769 92717
rect 68940 92712 69769 92714
rect 68940 92656 69708 92712
rect 69764 92656 69769 92712
rect 68940 92654 69769 92656
rect 68940 92652 68946 92654
rect 69703 92651 69769 92654
rect 70894 92652 70900 92716
rect 70964 92714 70970 92716
rect 71175 92714 71241 92717
rect 70964 92712 71241 92714
rect 70964 92656 71180 92712
rect 71236 92656 71241 92712
rect 70964 92654 71241 92656
rect 70964 92652 70970 92654
rect 71175 92651 71241 92654
rect 72366 92652 72372 92716
rect 72436 92714 72442 92716
rect 72831 92714 72897 92717
rect 72436 92712 72897 92714
rect 72436 92656 72836 92712
rect 72892 92656 72897 92712
rect 72436 92654 72897 92656
rect 72436 92652 72442 92654
rect 72831 92651 72897 92654
rect 91783 92714 91849 92717
rect 92238 92714 92244 92716
rect 91783 92712 92244 92714
rect 91783 92656 91788 92712
rect 91844 92656 92244 92712
rect 91783 92654 92244 92656
rect 91783 92651 91849 92654
rect 92238 92652 92244 92654
rect 92308 92652 92314 92716
rect 93255 92714 93321 92717
rect 93710 92714 93716 92716
rect 93255 92712 93716 92714
rect 93255 92656 93260 92712
rect 93316 92656 93716 92712
rect 93255 92654 93716 92656
rect 93255 92651 93321 92654
rect 93710 92652 93716 92654
rect 93780 92652 93786 92716
rect 194366 92714 194426 92926
rect 222653 92984 223436 92986
rect 222653 92928 222658 92984
rect 222714 92928 223436 92984
rect 222653 92926 223436 92928
rect 222653 92923 222719 92926
rect 223430 92924 223436 92926
rect 223500 92924 223506 92988
rect 201585 92852 201651 92853
rect 205449 92852 205515 92853
rect 208393 92852 208459 92853
rect 210049 92852 210115 92853
rect 201534 92850 201540 92852
rect 201494 92790 201540 92850
rect 201604 92848 201651 92852
rect 205398 92850 205404 92852
rect 201646 92792 201651 92848
rect 201534 92788 201540 92790
rect 201604 92788 201651 92792
rect 205358 92790 205404 92850
rect 205468 92848 205515 92852
rect 208342 92850 208348 92852
rect 205510 92792 205515 92848
rect 205398 92788 205404 92790
rect 205468 92788 205515 92792
rect 208302 92790 208348 92850
rect 208412 92848 208459 92852
rect 208454 92792 208459 92848
rect 208342 92788 208348 92790
rect 208412 92788 208459 92792
rect 209998 92788 210004 92852
rect 210068 92850 210115 92852
rect 220261 92850 220327 92853
rect 220670 92850 220676 92852
rect 210068 92848 210160 92850
rect 210110 92792 210160 92848
rect 210068 92790 210160 92792
rect 220261 92848 220676 92850
rect 220261 92792 220266 92848
rect 220322 92792 220676 92848
rect 220261 92790 220676 92792
rect 210068 92788 210115 92790
rect 201585 92787 201651 92788
rect 205449 92787 205515 92788
rect 208393 92787 208459 92788
rect 210049 92787 210115 92788
rect 220261 92787 220327 92790
rect 220670 92788 220676 92790
rect 220740 92788 220746 92852
rect 223941 92850 224007 92853
rect 224350 92850 224356 92852
rect 223941 92848 224356 92850
rect 223941 92792 223946 92848
rect 224002 92792 224356 92848
rect 223941 92790 224356 92792
rect 223941 92787 224007 92790
rect 224350 92788 224356 92790
rect 224420 92788 224426 92852
rect 196157 92714 196223 92717
rect 194366 92712 196223 92714
rect 194366 92656 196162 92712
rect 196218 92656 196223 92712
rect 194366 92654 196223 92656
rect 196157 92651 196223 92654
rect 215334 92652 215340 92716
rect 215404 92714 215410 92716
rect 216029 92714 216095 92717
rect 215404 92712 216095 92714
rect 215404 92656 216034 92712
rect 216090 92656 216095 92712
rect 215404 92654 216095 92656
rect 215404 92652 215410 92654
rect 216029 92651 216095 92654
rect 69841 92578 69907 92581
rect 67541 92576 69907 92578
rect 67541 92520 67546 92576
rect 67602 92520 69846 92576
rect 69902 92520 69907 92576
rect 67541 92518 69907 92520
rect 67541 92515 67607 92518
rect 69841 92515 69907 92518
rect 193438 92516 193444 92580
rect 193508 92578 193514 92580
rect 197353 92578 197419 92581
rect 193508 92576 197419 92578
rect 193508 92520 197358 92576
rect 197414 92520 197419 92576
rect 193508 92518 197419 92520
rect 193508 92516 193514 92518
rect 197353 92515 197419 92518
rect 198733 92578 198799 92581
rect 199469 92578 199535 92581
rect 269205 92578 269271 92581
rect 198733 92576 269271 92578
rect 198733 92520 198738 92576
rect 198794 92520 199474 92576
rect 199530 92520 269210 92576
rect 269266 92520 269271 92576
rect 198733 92518 269271 92520
rect 198733 92515 198799 92518
rect 199469 92515 199535 92518
rect 269205 92515 269271 92518
rect 71630 92380 71636 92444
rect 71700 92442 71706 92444
rect 81433 92442 81499 92445
rect 71700 92440 81499 92442
rect 71700 92384 81438 92440
rect 81494 92384 81499 92440
rect 71700 92382 81499 92384
rect 71700 92380 71706 92382
rect 81433 92379 81499 92382
rect 177941 92442 178007 92445
rect 196525 92442 196591 92445
rect 177941 92440 196591 92442
rect 177941 92384 177946 92440
rect 178002 92384 196530 92440
rect 196586 92384 196591 92440
rect 177941 92382 196591 92384
rect 177941 92379 178007 92382
rect 196525 92379 196591 92382
rect 199285 92442 199351 92445
rect 203006 92442 203012 92444
rect 199285 92440 203012 92442
rect 199285 92384 199290 92440
rect 199346 92384 203012 92440
rect 199285 92382 203012 92384
rect 199285 92379 199351 92382
rect 203006 92380 203012 92382
rect 203076 92380 203082 92444
rect 212574 92380 212580 92444
rect 212644 92442 212650 92444
rect 226517 92442 226583 92445
rect 212644 92440 226583 92442
rect 212644 92384 226522 92440
rect 226578 92384 226583 92440
rect 212644 92382 226583 92384
rect 212644 92380 212650 92382
rect 226517 92379 226583 92382
rect 83549 92306 83615 92309
rect 179413 92306 179479 92309
rect 83549 92304 179479 92306
rect 83549 92248 83554 92304
rect 83610 92248 179418 92304
rect 179474 92248 179479 92304
rect 83549 92246 179479 92248
rect 83549 92243 83615 92246
rect 179413 92243 179479 92246
rect 189809 92306 189875 92309
rect 202597 92306 202663 92309
rect 189809 92304 202663 92306
rect 189809 92248 189814 92304
rect 189870 92248 202602 92304
rect 202658 92248 202663 92304
rect 189809 92246 202663 92248
rect 189809 92243 189875 92246
rect 202597 92243 202663 92246
rect 92381 92170 92447 92173
rect 94814 92170 94820 92172
rect 92381 92168 94820 92170
rect 92381 92112 92386 92168
rect 92442 92112 94820 92168
rect 92381 92110 94820 92112
rect 92381 92107 92447 92110
rect 94814 92108 94820 92110
rect 94884 92108 94890 92172
rect 204846 91972 204852 92036
rect 204916 92034 204922 92036
rect 212574 92034 212580 92036
rect 204916 91974 212580 92034
rect 204916 91972 204922 91974
rect 212574 91972 212580 91974
rect 212644 91972 212650 92036
rect 212165 91898 212231 91901
rect 251265 91898 251331 91901
rect 212165 91896 251331 91898
rect 212165 91840 212170 91896
rect 212226 91840 251270 91896
rect 251326 91840 251331 91896
rect 212165 91838 251331 91840
rect 212165 91835 212231 91838
rect 251265 91835 251331 91838
rect 93117 91762 93183 91765
rect 96613 91762 96679 91765
rect 93117 91760 96679 91762
rect 93117 91704 93122 91760
rect 93178 91704 96618 91760
rect 96674 91704 96679 91760
rect 93117 91702 96679 91704
rect 93117 91699 93183 91702
rect 96613 91699 96679 91702
rect 108297 91762 108363 91765
rect 214557 91762 214623 91765
rect 108297 91760 214623 91762
rect 108297 91704 108302 91760
rect 108358 91704 214562 91760
rect 214618 91704 214623 91760
rect 108297 91702 214623 91704
rect 108297 91699 108363 91702
rect 214557 91699 214623 91702
rect 251265 91218 251331 91221
rect 251817 91218 251883 91221
rect 251265 91216 251883 91218
rect 251265 91160 251270 91216
rect 251326 91160 251822 91216
rect 251878 91160 251883 91216
rect 251265 91158 251883 91160
rect 251265 91155 251331 91158
rect 251817 91155 251883 91158
rect 71773 91082 71839 91085
rect 72734 91082 72740 91084
rect 71773 91080 72740 91082
rect 71773 91024 71778 91080
rect 71834 91024 72740 91080
rect 71773 91022 72740 91024
rect 71773 91019 71839 91022
rect 72734 91020 72740 91022
rect 72804 91020 72810 91084
rect 215845 90946 215911 90949
rect 219709 90946 219775 90949
rect 220721 90946 220787 90949
rect 215845 90944 220787 90946
rect 215845 90888 215850 90944
rect 215906 90888 219714 90944
rect 219770 90888 220726 90944
rect 220782 90888 220787 90944
rect 215845 90886 220787 90888
rect 215845 90883 215911 90886
rect 219709 90883 219775 90886
rect 220721 90883 220787 90886
rect 224309 90946 224375 90949
rect 255313 90946 255379 90949
rect 224309 90944 255379 90946
rect 224309 90888 224314 90944
rect 224370 90888 255318 90944
rect 255374 90888 255379 90944
rect 224309 90886 255379 90888
rect 224309 90883 224375 90886
rect 255313 90883 255379 90886
rect 105537 90674 105603 90677
rect 204437 90674 204503 90677
rect 105537 90672 204503 90674
rect 105537 90616 105542 90672
rect 105598 90616 204442 90672
rect 204498 90616 204503 90672
rect 105537 90614 204503 90616
rect 105537 90611 105603 90614
rect 204437 90611 204503 90614
rect 104157 90538 104223 90541
rect 203517 90538 203583 90541
rect 104157 90536 203583 90538
rect 104157 90480 104162 90536
rect 104218 90480 203522 90536
rect 203578 90480 203583 90536
rect 104157 90478 203583 90480
rect 104157 90475 104223 90478
rect 203517 90475 203583 90478
rect 50889 90402 50955 90405
rect 73061 90402 73127 90405
rect 50889 90400 73127 90402
rect 50889 90344 50894 90400
rect 50950 90344 73066 90400
rect 73122 90344 73127 90400
rect 50889 90342 73127 90344
rect 50889 90339 50955 90342
rect 73061 90339 73127 90342
rect 104341 90402 104407 90405
rect 203701 90402 203767 90405
rect 104341 90400 203767 90402
rect 104341 90344 104346 90400
rect 104402 90344 203706 90400
rect 203762 90344 203767 90400
rect 104341 90342 203767 90344
rect 104341 90339 104407 90342
rect 203701 90339 203767 90342
rect 201861 90266 201927 90269
rect 202781 90266 202847 90269
rect 201861 90264 202847 90266
rect 201861 90208 201866 90264
rect 201922 90208 202786 90264
rect 202842 90208 202847 90264
rect 201861 90206 202847 90208
rect 201861 90203 201927 90206
rect 202781 90203 202847 90206
rect 204345 90266 204411 90269
rect 205541 90266 205607 90269
rect 204345 90264 205607 90266
rect 204345 90208 204350 90264
rect 204406 90208 205546 90264
rect 205602 90208 205607 90264
rect 204345 90206 205607 90208
rect 204345 90203 204411 90206
rect 205541 90203 205607 90206
rect 208669 90266 208735 90269
rect 209681 90266 209747 90269
rect 208669 90264 209747 90266
rect 208669 90208 208674 90264
rect 208730 90208 209686 90264
rect 209742 90208 209747 90264
rect 208669 90206 209747 90208
rect 208669 90203 208735 90206
rect 209681 90203 209747 90206
rect 219525 89994 219591 89997
rect 220077 89994 220143 89997
rect 227713 89994 227779 89997
rect 219525 89992 227779 89994
rect 219525 89936 219530 89992
rect 219586 89936 220082 89992
rect 220138 89936 227718 89992
rect 227774 89936 227779 89992
rect 219525 89934 227779 89936
rect 219525 89931 219591 89934
rect 220077 89931 220143 89934
rect 227713 89931 227779 89934
rect 78397 89722 78463 89725
rect 113817 89722 113883 89725
rect 114369 89722 114435 89725
rect 78397 89720 114435 89722
rect 78397 89664 78402 89720
rect 78458 89664 113822 89720
rect 113878 89664 114374 89720
rect 114430 89664 114435 89720
rect 78397 89662 114435 89664
rect 78397 89659 78463 89662
rect 113817 89659 113883 89662
rect 114369 89659 114435 89662
rect 115289 89722 115355 89725
rect 209221 89722 209287 89725
rect 115289 89720 209287 89722
rect 115289 89664 115294 89720
rect 115350 89664 209226 89720
rect 209282 89664 209287 89720
rect 115289 89662 209287 89664
rect 115289 89659 115355 89662
rect 209221 89659 209287 89662
rect 214833 89722 214899 89725
rect 256693 89722 256759 89725
rect 214833 89720 256759 89722
rect 214833 89664 214838 89720
rect 214894 89664 256698 89720
rect 256754 89664 256759 89720
rect 214833 89662 256759 89664
rect 214833 89659 214899 89662
rect 256693 89659 256759 89662
rect 64597 89586 64663 89589
rect 98821 89586 98887 89589
rect 64597 89584 98887 89586
rect 64597 89528 64602 89584
rect 64658 89528 98826 89584
rect 98882 89528 98887 89584
rect 64597 89526 98887 89528
rect 64597 89523 64663 89526
rect 98821 89523 98887 89526
rect 185577 89586 185643 89589
rect 206093 89586 206159 89589
rect 185577 89584 206159 89586
rect 185577 89528 185582 89584
rect 185638 89528 206098 89584
rect 206154 89528 206159 89584
rect 185577 89526 206159 89528
rect 185577 89523 185643 89526
rect 206093 89523 206159 89526
rect 220629 89586 220695 89589
rect 243537 89586 243603 89589
rect 220629 89584 243603 89586
rect 220629 89528 220634 89584
rect 220690 89528 243542 89584
rect 243598 89528 243603 89584
rect 220629 89526 243603 89528
rect 220629 89523 220695 89526
rect 243537 89523 243603 89526
rect 84101 89450 84167 89453
rect 98494 89450 98500 89452
rect 84101 89448 98500 89450
rect 84101 89392 84106 89448
rect 84162 89392 98500 89448
rect 84101 89390 98500 89392
rect 84101 89387 84167 89390
rect 98494 89388 98500 89390
rect 98564 89388 98570 89452
rect 214557 89450 214623 89453
rect 226425 89450 226491 89453
rect 214557 89448 226491 89450
rect 214557 89392 214562 89448
rect 214618 89392 226430 89448
rect 226486 89392 226491 89448
rect 214557 89390 226491 89392
rect 214557 89387 214623 89390
rect 226425 89387 226491 89390
rect 227713 89042 227779 89045
rect 580257 89042 580323 89045
rect 227713 89040 580323 89042
rect 227713 88984 227718 89040
rect 227774 88984 580262 89040
rect 580318 88984 580323 89040
rect 227713 88982 580323 88984
rect 227713 88979 227779 88982
rect 580257 88979 580323 88982
rect 92749 88226 92815 88229
rect 119337 88226 119403 88229
rect 221917 88226 221983 88229
rect 92749 88224 221983 88226
rect 92749 88168 92754 88224
rect 92810 88168 119342 88224
rect 119398 88168 221922 88224
rect 221978 88168 221983 88224
rect 92749 88166 221983 88168
rect 92749 88163 92815 88166
rect 119337 88163 119403 88166
rect 221917 88163 221983 88166
rect 86677 88090 86743 88093
rect 100109 88090 100175 88093
rect 86677 88088 100175 88090
rect 86677 88032 86682 88088
rect 86738 88032 100114 88088
rect 100170 88032 100175 88088
rect 86677 88030 100175 88032
rect 86677 88027 86743 88030
rect 100109 88027 100175 88030
rect 191046 88028 191052 88092
rect 191116 88090 191122 88092
rect 204846 88090 204852 88092
rect 191116 88030 204852 88090
rect 191116 88028 191122 88030
rect 204846 88028 204852 88030
rect 204916 88028 204922 88092
rect 204989 88090 205055 88093
rect 284385 88090 284451 88093
rect 204989 88088 287070 88090
rect 204989 88032 204994 88088
rect 205050 88032 284390 88088
rect 284446 88032 287070 88088
rect 204989 88030 287070 88032
rect 204989 88027 205055 88030
rect 284385 88027 284451 88030
rect 66478 87892 66484 87956
rect 66548 87954 66554 87956
rect 94773 87954 94839 87957
rect 66548 87952 94839 87954
rect 66548 87896 94778 87952
rect 94834 87896 94839 87952
rect 66548 87894 94839 87896
rect 66548 87892 66554 87894
rect 94773 87891 94839 87894
rect 187601 87954 187667 87957
rect 224902 87954 224908 87956
rect 187601 87952 224908 87954
rect 187601 87896 187606 87952
rect 187662 87896 224908 87952
rect 187601 87894 224908 87896
rect 187601 87891 187667 87894
rect 224902 87892 224908 87894
rect 224972 87892 224978 87956
rect 287010 87546 287070 88030
rect 582925 87546 582991 87549
rect 287010 87544 582991 87546
rect 287010 87488 582930 87544
rect 582986 87488 582991 87544
rect 287010 87486 582991 87488
rect 582925 87483 582991 87486
rect 86125 86866 86191 86869
rect 95141 86866 95207 86869
rect 86125 86864 95207 86866
rect 86125 86808 86130 86864
rect 86186 86808 95146 86864
rect 95202 86808 95207 86864
rect 86125 86806 95207 86808
rect 86125 86803 86191 86806
rect 95141 86803 95207 86806
rect 204437 86866 204503 86869
rect 288617 86866 288683 86869
rect 289721 86866 289787 86869
rect 204437 86864 289787 86866
rect 204437 86808 204442 86864
rect 204498 86808 288622 86864
rect 288678 86808 289726 86864
rect 289782 86808 289787 86864
rect 204437 86806 289787 86808
rect 204437 86803 204503 86806
rect 288617 86803 288683 86806
rect 289721 86803 289787 86806
rect 67357 86730 67423 86733
rect 100017 86730 100083 86733
rect 67357 86728 100083 86730
rect 67357 86672 67362 86728
rect 67418 86672 100022 86728
rect 100078 86672 100083 86728
rect 67357 86670 100083 86672
rect 67357 86667 67423 86670
rect 100017 86667 100083 86670
rect 180057 86730 180123 86733
rect 200757 86730 200823 86733
rect 180057 86728 200823 86730
rect 180057 86672 180062 86728
rect 180118 86672 200762 86728
rect 200818 86672 200823 86728
rect 180057 86670 200823 86672
rect 180057 86667 180123 86670
rect 200757 86667 200823 86670
rect 71773 86594 71839 86597
rect 197077 86594 197143 86597
rect 71773 86592 197143 86594
rect 71773 86536 71778 86592
rect 71834 86536 197082 86592
rect 197138 86536 197143 86592
rect 71773 86534 197143 86536
rect 71773 86531 71839 86534
rect 197077 86531 197143 86534
rect 192569 86186 192635 86189
rect 259545 86186 259611 86189
rect 583520 86186 584960 86276
rect 192569 86184 259611 86186
rect 192569 86128 192574 86184
rect 192630 86128 259550 86184
rect 259606 86128 259611 86184
rect 192569 86126 259611 86128
rect 192569 86123 192635 86126
rect 259545 86123 259611 86126
rect 583342 86126 584960 86186
rect 583342 86050 583402 86126
rect 583520 86050 584960 86126
rect 583342 86036 584960 86050
rect 583342 85990 583586 86036
rect 289721 85642 289787 85645
rect 583526 85642 583586 85990
rect 289721 85640 583586 85642
rect 289721 85584 289726 85640
rect 289782 85584 583586 85640
rect 289721 85582 583586 85584
rect 289721 85579 289787 85582
rect 66069 85506 66135 85509
rect 187734 85506 187740 85508
rect 66069 85504 187740 85506
rect 66069 85448 66074 85504
rect 66130 85448 187740 85504
rect 66069 85446 187740 85448
rect 66069 85443 66135 85446
rect 187734 85444 187740 85446
rect 187804 85506 187810 85508
rect 188337 85506 188403 85509
rect 187804 85504 188403 85506
rect 187804 85448 188342 85504
rect 188398 85448 188403 85504
rect 187804 85446 188403 85448
rect 187804 85444 187810 85446
rect 188337 85443 188403 85446
rect 79501 85370 79567 85373
rect 95182 85370 95188 85372
rect 79501 85368 95188 85370
rect 79501 85312 79506 85368
rect 79562 85312 95188 85368
rect 79501 85310 95188 85312
rect 79501 85307 79567 85310
rect 95182 85308 95188 85310
rect 95252 85308 95258 85372
rect 182909 85370 182975 85373
rect 200389 85370 200455 85373
rect 201309 85370 201375 85373
rect 182909 85368 201375 85370
rect 182909 85312 182914 85368
rect 182970 85312 200394 85368
rect 200450 85312 201314 85368
rect 201370 85312 201375 85368
rect 182909 85310 201375 85312
rect 182909 85307 182975 85310
rect 200389 85307 200455 85310
rect 201309 85307 201375 85310
rect -960 84690 480 84780
rect 3141 84690 3207 84693
rect -960 84688 3207 84690
rect -960 84632 3146 84688
rect 3202 84632 3207 84688
rect -960 84630 3207 84632
rect -960 84540 480 84630
rect 3141 84627 3207 84630
rect 191097 84282 191163 84285
rect 191465 84282 191531 84285
rect 309777 84282 309843 84285
rect 191097 84280 309843 84282
rect 191097 84224 191102 84280
rect 191158 84224 191470 84280
rect 191526 84224 309782 84280
rect 309838 84224 309843 84280
rect 191097 84222 309843 84224
rect 191097 84219 191163 84222
rect 191465 84219 191531 84222
rect 309777 84219 309843 84222
rect 91093 84146 91159 84149
rect 219433 84146 219499 84149
rect 91093 84144 219499 84146
rect 91093 84088 91098 84144
rect 91154 84088 219438 84144
rect 219494 84088 219499 84144
rect 91093 84086 219499 84088
rect 91093 84083 91159 84086
rect 219433 84083 219499 84086
rect 178769 84010 178835 84013
rect 230473 84010 230539 84013
rect 178769 84008 230539 84010
rect 178769 83952 178774 84008
rect 178830 83952 230478 84008
rect 230534 83952 230539 84008
rect 178769 83950 230539 83952
rect 178769 83947 178835 83950
rect 230473 83947 230539 83950
rect 3417 83466 3483 83469
rect 95325 83466 95391 83469
rect 3417 83464 95391 83466
rect 3417 83408 3422 83464
rect 3478 83408 95330 83464
rect 95386 83408 95391 83464
rect 3417 83406 95391 83408
rect 3417 83403 3483 83406
rect 95325 83403 95391 83406
rect 209773 82786 209839 82789
rect 281533 82786 281599 82789
rect 209773 82784 281599 82786
rect 209773 82728 209778 82784
rect 209834 82728 281538 82784
rect 281594 82728 281599 82784
rect 209773 82726 281599 82728
rect 209773 82723 209839 82726
rect 281533 82723 281599 82726
rect 89989 82650 90055 82653
rect 98729 82650 98795 82653
rect 89989 82648 98795 82650
rect 89989 82592 89994 82648
rect 90050 82592 98734 82648
rect 98790 82592 98795 82648
rect 89989 82590 98795 82592
rect 89989 82587 90055 82590
rect 98729 82587 98795 82590
rect 157977 82650 158043 82653
rect 226374 82650 226380 82652
rect 157977 82648 226380 82650
rect 157977 82592 157982 82648
rect 158038 82592 226380 82648
rect 157977 82590 226380 82592
rect 157977 82587 158043 82590
rect 226374 82588 226380 82590
rect 226444 82588 226450 82652
rect 82813 82514 82879 82517
rect 209998 82514 210004 82516
rect 82813 82512 210004 82514
rect 82813 82456 82818 82512
rect 82874 82456 210004 82512
rect 82813 82454 210004 82456
rect 82813 82451 82879 82454
rect 209998 82452 210004 82454
rect 210068 82452 210074 82516
rect 184289 81426 184355 81429
rect 227989 81426 228055 81429
rect 184289 81424 228055 81426
rect 184289 81368 184294 81424
rect 184350 81368 227994 81424
rect 228050 81368 228055 81424
rect 184289 81366 228055 81368
rect 184289 81363 184355 81366
rect 227989 81363 228055 81366
rect 77569 81290 77635 81293
rect 105537 81290 105603 81293
rect 77569 81288 105603 81290
rect 77569 81232 77574 81288
rect 77630 81232 105542 81288
rect 105598 81232 105603 81288
rect 77569 81230 105603 81232
rect 77569 81227 77635 81230
rect 105537 81227 105603 81230
rect 61745 81154 61811 81157
rect 187049 81154 187115 81157
rect 61745 81152 187115 81154
rect 61745 81096 61750 81152
rect 61806 81096 187054 81152
rect 187110 81096 187115 81152
rect 61745 81094 187115 81096
rect 61745 81091 61811 81094
rect 187049 81091 187115 81094
rect 192702 80684 192708 80748
rect 192772 80746 192778 80748
rect 327073 80746 327139 80749
rect 192772 80744 327139 80746
rect 192772 80688 327078 80744
rect 327134 80688 327139 80744
rect 192772 80686 327139 80688
rect 192772 80684 192778 80686
rect 327073 80683 327139 80686
rect 77293 80066 77359 80069
rect 104341 80066 104407 80069
rect 77293 80064 104407 80066
rect 77293 80008 77298 80064
rect 77354 80008 104346 80064
rect 104402 80008 104407 80064
rect 77293 80006 104407 80008
rect 77293 80003 77359 80006
rect 104341 80003 104407 80006
rect 204161 80066 204227 80069
rect 241605 80066 241671 80069
rect 204161 80064 241671 80066
rect 204161 80008 204166 80064
rect 204222 80008 241610 80064
rect 241666 80008 241671 80064
rect 204161 80006 241671 80008
rect 204161 80003 204227 80006
rect 241605 80003 241671 80006
rect 184381 79930 184447 79933
rect 213269 79930 213335 79933
rect 184381 79928 213335 79930
rect 184381 79872 184386 79928
rect 184442 79872 213274 79928
rect 213330 79872 213335 79928
rect 184381 79870 213335 79872
rect 184381 79867 184447 79870
rect 213269 79867 213335 79870
rect 111149 79794 111215 79797
rect 204345 79794 204411 79797
rect 111149 79792 204411 79794
rect 111149 79736 111154 79792
rect 111210 79736 204350 79792
rect 204406 79736 204411 79792
rect 111149 79734 204411 79736
rect 111149 79731 111215 79734
rect 204345 79731 204411 79734
rect 203517 79658 203583 79661
rect 204161 79658 204227 79661
rect 203517 79656 204227 79658
rect 203517 79600 203522 79656
rect 203578 79600 204166 79656
rect 204222 79600 204227 79656
rect 203517 79598 204227 79600
rect 203517 79595 203583 79598
rect 204161 79595 204227 79598
rect 204345 79522 204411 79525
rect 204897 79522 204963 79525
rect 204345 79520 204963 79522
rect 204345 79464 204350 79520
rect 204406 79464 204902 79520
rect 204958 79464 204963 79520
rect 204345 79462 204963 79464
rect 204345 79459 204411 79462
rect 204897 79459 204963 79462
rect 197445 78570 197511 78573
rect 273345 78570 273411 78573
rect 582649 78570 582715 78573
rect 197445 78568 582715 78570
rect 197445 78512 197450 78568
rect 197506 78512 273350 78568
rect 273406 78512 582654 78568
rect 582710 78512 582715 78568
rect 197445 78510 582715 78512
rect 197445 78507 197511 78510
rect 273345 78507 273411 78510
rect 582649 78507 582715 78510
rect 193029 78434 193095 78437
rect 238109 78434 238175 78437
rect 193029 78432 238175 78434
rect 193029 78376 193034 78432
rect 193090 78376 238114 78432
rect 238170 78376 238175 78432
rect 193029 78374 238175 78376
rect 193029 78371 193095 78374
rect 238109 78371 238175 78374
rect 73061 78026 73127 78029
rect 101397 78026 101463 78029
rect 73061 78024 101463 78026
rect 73061 77968 73066 78024
rect 73122 77968 101402 78024
rect 101458 77968 101463 78024
rect 73061 77966 101463 77968
rect 73061 77963 73127 77966
rect 101397 77963 101463 77966
rect 70301 77890 70367 77893
rect 182817 77890 182883 77893
rect 70301 77888 182883 77890
rect 70301 77832 70306 77888
rect 70362 77832 182822 77888
rect 182878 77832 182883 77888
rect 70301 77830 182883 77832
rect 70301 77827 70367 77830
rect 182817 77827 182883 77830
rect 89897 77210 89963 77213
rect 220077 77210 220143 77213
rect 89897 77208 220143 77210
rect 89897 77152 89902 77208
rect 89958 77152 220082 77208
rect 220138 77152 220143 77208
rect 89897 77150 220143 77152
rect 89897 77147 89963 77150
rect 220077 77147 220143 77150
rect 196566 76468 196572 76532
rect 196636 76530 196642 76532
rect 262213 76530 262279 76533
rect 196636 76528 262279 76530
rect 196636 76472 262218 76528
rect 262274 76472 262279 76528
rect 196636 76470 262279 76472
rect 196636 76468 196642 76470
rect 262213 76467 262279 76470
rect 193305 75850 193371 75853
rect 193857 75850 193923 75853
rect 269113 75850 269179 75853
rect 193305 75848 269179 75850
rect 193305 75792 193310 75848
rect 193366 75792 193862 75848
rect 193918 75792 269118 75848
rect 269174 75792 269179 75848
rect 193305 75790 269179 75792
rect 193305 75787 193371 75790
rect 193857 75787 193923 75790
rect 269113 75787 269179 75790
rect 75821 75170 75887 75173
rect 167637 75170 167703 75173
rect 75821 75168 167703 75170
rect 75821 75112 75826 75168
rect 75882 75112 167642 75168
rect 167698 75112 167703 75168
rect 75821 75110 167703 75112
rect 75821 75107 75887 75110
rect 167637 75107 167703 75110
rect 76557 73810 76623 73813
rect 230606 73810 230612 73812
rect 76557 73808 230612 73810
rect 76557 73752 76562 73808
rect 76618 73752 230612 73808
rect 76557 73750 230612 73752
rect 76557 73747 76623 73750
rect 230606 73748 230612 73750
rect 230676 73748 230682 73812
rect 580257 72994 580323 72997
rect 583520 72994 584960 73084
rect 580257 72992 584960 72994
rect 580257 72936 580262 72992
rect 580318 72936 584960 72992
rect 580257 72934 584960 72936
rect 580257 72931 580323 72934
rect 583520 72844 584960 72934
rect 91001 72450 91067 72453
rect 234613 72450 234679 72453
rect 91001 72448 234679 72450
rect 91001 72392 91006 72448
rect 91062 72392 234618 72448
rect 234674 72392 234679 72448
rect 91001 72390 234679 72392
rect 91001 72387 91067 72390
rect 234613 72387 234679 72390
rect 187693 71770 187759 71773
rect 188889 71770 188955 71773
rect 274582 71770 274588 71772
rect 187693 71768 274588 71770
rect -960 71634 480 71724
rect 187693 71712 187698 71768
rect 187754 71712 188894 71768
rect 188950 71712 274588 71768
rect 187693 71710 274588 71712
rect 187693 71707 187759 71710
rect 188889 71707 188955 71710
rect 274582 71708 274588 71710
rect 274652 71770 274658 71772
rect 274652 71710 277410 71770
rect 274652 71708 274658 71710
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 277350 71090 277410 71710
rect 288433 71090 288499 71093
rect 277350 71088 288499 71090
rect 277350 71032 288438 71088
rect 288494 71032 288499 71088
rect 277350 71030 288499 71032
rect 288433 71027 288499 71030
rect 98637 69594 98703 69597
rect 232078 69594 232084 69596
rect 98637 69592 232084 69594
rect 98637 69536 98642 69592
rect 98698 69536 232084 69592
rect 98637 69534 232084 69536
rect 98637 69531 98703 69534
rect 232078 69532 232084 69534
rect 232148 69532 232154 69596
rect 194593 66194 194659 66197
rect 195237 66194 195303 66197
rect 247718 66194 247724 66196
rect 194593 66192 247724 66194
rect 194593 66136 194598 66192
rect 194654 66136 195242 66192
rect 195298 66136 247724 66192
rect 194593 66134 247724 66136
rect 194593 66131 194659 66134
rect 195237 66131 195303 66134
rect 247718 66132 247724 66134
rect 247788 66132 247794 66196
rect 67265 63474 67331 63477
rect 193806 63474 193812 63476
rect 67265 63472 193812 63474
rect 67265 63416 67270 63472
rect 67326 63416 193812 63472
rect 67265 63414 193812 63416
rect 67265 63411 67331 63414
rect 193806 63412 193812 63414
rect 193876 63412 193882 63476
rect 84101 61434 84167 61437
rect 233182 61434 233188 61436
rect 84101 61432 233188 61434
rect 84101 61376 84106 61432
rect 84162 61376 233188 61432
rect 84101 61374 233188 61376
rect 84101 61371 84167 61374
rect 233182 61372 233188 61374
rect 233252 61372 233258 61436
rect 193806 60556 193812 60620
rect 193876 60618 193882 60620
rect 285673 60618 285739 60621
rect 286409 60618 286475 60621
rect 193876 60616 286475 60618
rect 193876 60560 285678 60616
rect 285734 60560 286414 60616
rect 286470 60560 286475 60616
rect 193876 60558 286475 60560
rect 193876 60556 193882 60558
rect 285673 60555 285739 60558
rect 286409 60555 286475 60558
rect 583017 59666 583083 59669
rect 583520 59666 584960 59756
rect 583017 59664 584960 59666
rect 583017 59608 583022 59664
rect 583078 59608 584960 59664
rect 583017 59606 584960 59608
rect 583017 59603 583083 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 2957 58578 3023 58581
rect -960 58576 3023 58578
rect -960 58520 2962 58576
rect 3018 58520 3023 58576
rect -960 58518 3023 58520
rect -960 58428 480 58518
rect 2957 58515 3023 58518
rect 95141 54498 95207 54501
rect 234654 54498 234660 54500
rect 95141 54496 234660 54498
rect 95141 54440 95146 54496
rect 95202 54440 234660 54496
rect 95141 54438 234660 54440
rect 95141 54435 95207 54438
rect 234654 54436 234660 54438
rect 234724 54436 234730 54500
rect 88241 48922 88307 48925
rect 233550 48922 233556 48924
rect 88241 48920 233556 48922
rect 88241 48864 88246 48920
rect 88302 48864 233556 48920
rect 88241 48862 233556 48864
rect 88241 48859 88307 48862
rect 233550 48860 233556 48862
rect 233620 48860 233626 48924
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 582833 33146 582899 33149
rect 583520 33146 584960 33236
rect 582833 33144 584960 33146
rect 582833 33088 582838 33144
rect 582894 33088 584960 33144
rect 582833 33086 584960 33088
rect 582833 33083 582899 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3509 32466 3575 32469
rect -960 32464 3575 32466
rect -960 32408 3514 32464
rect 3570 32408 3575 32464
rect -960 32406 3575 32408
rect -960 32316 480 32406
rect 3509 32403 3575 32406
rect 582557 19818 582623 19821
rect 583520 19818 584960 19908
rect 582557 19816 584960 19818
rect 582557 19760 582562 19816
rect 582618 19760 584960 19816
rect 582557 19758 584960 19760
rect 582557 19755 582623 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 81341 14514 81407 14517
rect 232262 14514 232268 14516
rect 81341 14512 232268 14514
rect 81341 14456 81346 14512
rect 81402 14456 232268 14512
rect 81341 14454 232268 14456
rect 81341 14451 81407 14454
rect 232262 14452 232268 14454
rect 232332 14452 232338 14516
rect 197854 7516 197860 7580
rect 197924 7578 197930 7580
rect 301957 7578 302023 7581
rect 197924 7576 302023 7578
rect 197924 7520 301962 7576
rect 302018 7520 302023 7576
rect 197924 7518 302023 7520
rect 197924 7516 197930 7518
rect 301957 7515 302023 7518
rect 582925 6626 582991 6629
rect 583520 6626 584960 6716
rect 582925 6624 584960 6626
rect -960 6490 480 6580
rect 582925 6568 582930 6624
rect 582986 6568 584960 6624
rect 582925 6566 584960 6568
rect 582925 6563 582991 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 73797 6218 73863 6221
rect 230422 6218 230428 6220
rect 73797 6216 230428 6218
rect 73797 6160 73802 6216
rect 73858 6160 230428 6216
rect 73797 6158 230428 6160
rect 73797 6155 73863 6158
rect 230422 6156 230428 6158
rect 230492 6156 230498 6220
rect 305637 6218 305703 6221
rect 319713 6218 319779 6221
rect 305637 6216 319779 6218
rect 305637 6160 305642 6216
rect 305698 6160 319718 6216
rect 319774 6160 319779 6216
rect 305637 6158 319779 6160
rect 305637 6155 305703 6158
rect 319713 6155 319779 6158
rect 110505 3498 110571 3501
rect 111558 3498 111564 3500
rect 110505 3496 111564 3498
rect 110505 3440 110510 3496
rect 110566 3440 111564 3496
rect 110505 3438 111564 3440
rect 110505 3435 110571 3438
rect 111558 3436 111564 3438
rect 111628 3436 111634 3500
rect 348049 3498 348115 3501
rect 353293 3498 353359 3501
rect 348049 3496 353359 3498
rect 348049 3440 348054 3496
rect 348110 3440 353298 3496
rect 353354 3440 353359 3496
rect 348049 3438 353359 3440
rect 348049 3435 348115 3438
rect 353293 3435 353359 3438
rect 63217 3362 63283 3365
rect 100293 3362 100359 3365
rect 63217 3360 100359 3362
rect 63217 3304 63222 3360
rect 63278 3304 100298 3360
rect 100354 3304 100359 3360
rect 63217 3302 100359 3304
rect 63217 3299 63283 3302
rect 100293 3299 100359 3302
<< via3 >>
rect 258580 702476 258644 702540
rect 75868 585108 75932 585172
rect 80652 581164 80716 581228
rect 75684 581028 75748 581092
rect 101260 581028 101324 581092
rect 70348 580756 70412 580820
rect 79916 580816 79980 580820
rect 79916 580760 79930 580816
rect 79930 580760 79980 580816
rect 79916 580756 79980 580760
rect 83964 580756 84028 580820
rect 88932 580816 88996 580820
rect 88932 580760 88946 580816
rect 88946 580760 88996 580816
rect 88932 580756 88996 580760
rect 92612 580816 92676 580820
rect 92612 580760 92626 580816
rect 92626 580760 92676 580816
rect 92612 580756 92676 580760
rect 104940 565796 105004 565860
rect 67772 561988 67836 562052
rect 96660 554100 96724 554164
rect 100708 549340 100772 549404
rect 96844 547028 96908 547092
rect 69060 546756 69124 546820
rect 67956 543356 68020 543420
rect 69244 541588 69308 541652
rect 75868 539548 75932 539612
rect 96844 537372 96908 537436
rect 105124 535468 105188 535532
rect 79732 534652 79796 534716
rect 72740 523636 72804 523700
rect 114508 522276 114572 522340
rect 69796 520916 69860 520980
rect 88748 520916 88812 520980
rect 67772 482156 67836 482220
rect 91324 482156 91388 482220
rect 73292 478076 73356 478140
rect 92612 478076 92676 478140
rect 69612 476716 69676 476780
rect 104204 476716 104268 476780
rect 75868 475356 75932 475420
rect 96844 473996 96908 474060
rect 111932 472500 111996 472564
rect 67956 471820 68020 471884
rect 67772 467876 67836 467940
rect 70348 467876 70412 467940
rect 269068 465156 269132 465220
rect 75684 464340 75748 464404
rect 258580 462844 258644 462908
rect 114324 460124 114388 460188
rect 101996 459580 102060 459644
rect 253060 458492 253124 458556
rect 197124 458280 197188 458284
rect 197124 458224 197138 458280
rect 197138 458224 197188 458280
rect 197124 458220 197188 458224
rect 80652 456044 80716 456108
rect 96660 456104 96724 456108
rect 96660 456048 96674 456104
rect 96674 456048 96724 456104
rect 96660 456044 96724 456048
rect 96660 455908 96724 455972
rect 267780 455636 267844 455700
rect 266492 454140 266556 454204
rect 194548 453052 194612 453116
rect 241652 452916 241716 452980
rect 247724 451556 247788 451620
rect 193812 450332 193876 450396
rect 194548 450256 194612 450260
rect 194548 450200 194598 450256
rect 194598 450200 194612 450256
rect 194548 450196 194612 450200
rect 256740 450060 256804 450124
rect 244412 449924 244476 449988
rect 249748 449924 249812 449988
rect 193444 449712 193508 449716
rect 193444 449656 193494 449712
rect 193494 449656 193508 449712
rect 193444 449652 193508 449656
rect 242940 449712 243004 449716
rect 242940 449656 242990 449712
rect 242990 449656 243004 449712
rect 242940 449652 243004 449656
rect 96476 446388 96540 446452
rect 193444 442852 193508 442916
rect 258396 442036 258460 442100
rect 107700 440812 107764 440876
rect 192708 440676 192772 440740
rect 67956 440268 68020 440332
rect 252876 440268 252940 440332
rect 69428 438908 69492 438972
rect 88932 438772 88996 438836
rect 88932 438228 88996 438292
rect 101996 438092 102060 438156
rect 112116 438092 112180 438156
rect 82124 437412 82188 437476
rect 83964 437412 84028 437476
rect 113220 436792 113284 436796
rect 113220 436736 113270 436792
rect 113270 436736 113284 436792
rect 113220 436732 113284 436736
rect 253060 436732 253124 436796
rect 95004 436460 95068 436524
rect 96292 436324 96356 436388
rect 73660 436188 73724 436252
rect 83964 436188 84028 436252
rect 102732 436052 102796 436116
rect 118740 434828 118804 434892
rect 70164 434556 70228 434620
rect 92980 434556 93044 434620
rect 71636 434420 71700 434484
rect 72556 433740 72620 433804
rect 90220 433740 90284 433804
rect 94452 433740 94516 433804
rect 99972 433740 100036 433804
rect 74580 433604 74644 433668
rect 76420 433664 76484 433668
rect 76420 433608 76434 433664
rect 76434 433608 76484 433664
rect 76420 433604 76484 433608
rect 77340 433604 77404 433668
rect 81940 433664 82004 433668
rect 81940 433608 81954 433664
rect 81954 433608 82004 433664
rect 81940 433604 82004 433608
rect 84700 433664 84764 433668
rect 84700 433608 84714 433664
rect 84714 433608 84764 433664
rect 84700 433604 84764 433608
rect 85804 433604 85868 433668
rect 87092 433604 87156 433668
rect 87460 433604 87524 433668
rect 91140 433664 91204 433668
rect 91140 433608 91190 433664
rect 91190 433608 91204 433664
rect 91140 433604 91204 433608
rect 92612 433604 92676 433668
rect 96476 433604 96540 433668
rect 98132 433664 98196 433668
rect 98132 433608 98182 433664
rect 98182 433608 98196 433664
rect 98132 433604 98196 433608
rect 98316 433604 98380 433668
rect 100156 433604 100220 433668
rect 102548 433604 102612 433668
rect 106412 433604 106476 433668
rect 108988 433664 109052 433668
rect 108988 433608 109038 433664
rect 109038 433608 109052 433664
rect 108988 433604 109052 433608
rect 110644 433664 110708 433668
rect 110644 433608 110694 433664
rect 110694 433608 110708 433664
rect 110644 433604 110708 433608
rect 111748 433664 111812 433668
rect 111748 433608 111798 433664
rect 111798 433608 111812 433664
rect 111748 433604 111812 433608
rect 112116 432788 112180 432852
rect 193444 432516 193508 432580
rect 193260 430884 193324 430948
rect 69428 426124 69492 426188
rect 262260 424220 262324 424284
rect 188844 420956 188908 421020
rect 114324 418236 114388 418300
rect 114692 417828 114756 417892
rect 188292 414020 188356 414084
rect 114508 410484 114572 410548
rect 67772 409668 67836 409732
rect 59124 405724 59188 405788
rect 252876 404772 252940 404836
rect 270540 403548 270604 403612
rect 66668 398788 66732 398852
rect 160692 396612 160756 396676
rect 67956 396340 68020 396404
rect 113220 396340 113284 396404
rect 253980 395524 254044 395588
rect 193812 392532 193876 392596
rect 69612 391988 69676 392052
rect 193260 391232 193324 391236
rect 193260 391176 193310 391232
rect 193310 391176 193324 391232
rect 193260 391172 193324 391176
rect 73476 390900 73540 390964
rect 82124 390688 82188 390692
rect 82124 390632 82138 390688
rect 82138 390632 82188 390688
rect 82124 390628 82188 390632
rect 96476 390628 96540 390692
rect 96660 390688 96724 390692
rect 96660 390632 96710 390688
rect 96710 390632 96724 390688
rect 96660 390628 96724 390632
rect 104204 390688 104268 390692
rect 104204 390632 104254 390688
rect 104254 390632 104268 390688
rect 104204 390628 104268 390632
rect 105124 390688 105188 390692
rect 105124 390632 105138 390688
rect 105138 390632 105188 390688
rect 105124 390628 105188 390632
rect 107700 390688 107764 390692
rect 107700 390632 107750 390688
rect 107750 390632 107764 390688
rect 107700 390628 107764 390632
rect 111932 390688 111996 390692
rect 111932 390632 111982 390688
rect 111982 390632 111996 390688
rect 111932 390628 111996 390632
rect 88748 390492 88812 390556
rect 100708 390492 100772 390556
rect 91324 390356 91388 390420
rect 96844 390356 96908 390420
rect 104940 390492 105004 390556
rect 253980 389132 254044 389196
rect 72740 388996 72804 389060
rect 79732 388996 79796 389060
rect 80100 389056 80164 389060
rect 80100 389000 80150 389056
rect 80150 389000 80164 389056
rect 80100 388996 80164 389000
rect 100156 388452 100220 388516
rect 102548 388452 102612 388516
rect 281580 388316 281644 388380
rect 70348 388180 70412 388244
rect 95004 388180 95068 388244
rect 93900 387908 93964 387972
rect 68876 387772 68940 387836
rect 188292 387500 188356 387564
rect 266308 387636 266372 387700
rect 86724 386956 86788 387020
rect 201540 386956 201604 387020
rect 263548 386276 263612 386340
rect 285628 386336 285692 386340
rect 285628 386280 285678 386336
rect 285678 386280 285692 386336
rect 285628 386276 285692 386280
rect 208348 385596 208412 385660
rect 285628 385596 285692 385660
rect 244412 384372 244476 384436
rect 66668 384236 66732 384300
rect 242940 384236 243004 384300
rect 216444 384024 216508 384028
rect 216444 383968 216458 384024
rect 216458 383968 216508 384024
rect 216444 383964 216508 383968
rect 74580 383692 74644 383756
rect 96292 383692 96356 383756
rect 87460 382876 87524 382940
rect 114692 382876 114756 382940
rect 69612 380836 69676 380900
rect 192708 380156 192772 380220
rect 276244 379536 276308 379540
rect 276244 379480 276258 379536
rect 276258 379480 276308 379536
rect 276244 379476 276308 379480
rect 242756 377980 242820 378044
rect 67772 376620 67836 376684
rect 197124 375940 197188 376004
rect 203012 375940 203076 376004
rect 258396 375260 258460 375324
rect 160692 372540 160756 372604
rect 236500 370636 236564 370700
rect 247724 370636 247788 370700
rect 252692 368324 252756 368388
rect 218652 366284 218716 366348
rect 249748 366284 249812 366348
rect 215156 364924 215220 364988
rect 269252 363020 269316 363084
rect 221228 360844 221292 360908
rect 193812 357988 193876 358052
rect 267964 357988 268028 358052
rect 72740 356628 72804 356692
rect 188844 355404 188908 355468
rect 68876 355268 68940 355332
rect 266492 339552 266556 339556
rect 266492 339496 266506 339552
rect 266506 339496 266556 339552
rect 266492 339492 266556 339496
rect 193812 338676 193876 338740
rect 72556 338132 72620 338196
rect 252508 338056 252572 338060
rect 252508 338000 252558 338056
rect 252558 338000 252572 338056
rect 252508 337996 252572 338000
rect 238892 337316 238956 337380
rect 252692 336636 252756 336700
rect 252508 334596 252572 334660
rect 262444 332556 262508 332620
rect 260972 331740 261036 331804
rect 252324 328340 252388 328404
rect 252324 327116 252388 327180
rect 77340 326300 77404 326364
rect 110644 323580 110708 323644
rect 199332 323036 199396 323100
rect 217180 322900 217244 322964
rect 66484 322084 66548 322148
rect 94452 320724 94516 320788
rect 85804 320180 85868 320244
rect 102732 320240 102796 320244
rect 102732 320184 102746 320240
rect 102746 320184 102796 320240
rect 102732 320180 102796 320184
rect 98132 319364 98196 319428
rect 111748 319364 111812 319428
rect 84700 318684 84764 318748
rect 106412 318004 106476 318068
rect 270724 318004 270788 318068
rect 81940 317460 82004 317524
rect 90220 316780 90284 316844
rect 118740 316644 118804 316708
rect 191604 316644 191668 316708
rect 263732 316644 263796 316708
rect 260052 316508 260116 316572
rect 259500 313924 259564 313988
rect 277164 313924 277228 313988
rect 256740 309436 256804 309500
rect 206140 307668 206204 307732
rect 224172 307668 224236 307732
rect 255268 306988 255332 307052
rect 230244 306444 230308 306508
rect 273300 305764 273364 305828
rect 108988 305628 109052 305692
rect 184060 305220 184124 305284
rect 220492 305220 220556 305284
rect 81940 304948 82004 305012
rect 91140 305084 91204 305148
rect 226196 305084 226260 305148
rect 241468 305084 241532 305148
rect 90956 304948 91020 305012
rect 241652 304132 241716 304196
rect 217548 303860 217612 303924
rect 186820 303724 186884 303788
rect 213684 303724 213748 303788
rect 211660 303588 211724 303652
rect 274588 303724 274652 303788
rect 200620 303452 200684 303516
rect 99972 302772 100036 302836
rect 192708 302288 192772 302292
rect 192708 302232 192758 302288
rect 192758 302232 192772 302288
rect 192708 302228 192772 302232
rect 194548 302228 194612 302292
rect 214420 302228 214484 302292
rect 240732 302228 240796 302292
rect 220860 301820 220924 301884
rect 191604 301548 191668 301612
rect 193260 301548 193324 301612
rect 91140 301412 91204 301476
rect 204300 301472 204364 301476
rect 204300 301416 204350 301472
rect 204350 301416 204364 301472
rect 204300 301412 204364 301416
rect 207060 301472 207124 301476
rect 207060 301416 207074 301472
rect 207074 301416 207124 301472
rect 207060 301412 207124 301416
rect 210556 301472 210620 301476
rect 210556 301416 210606 301472
rect 210606 301416 210620 301472
rect 210556 301412 210620 301416
rect 215892 301412 215956 301476
rect 219204 301412 219268 301476
rect 222332 301548 222396 301612
rect 226564 301548 226628 301612
rect 230428 301548 230492 301612
rect 234660 301548 234724 301612
rect 237604 301548 237668 301612
rect 222700 301412 222764 301476
rect 223620 301412 223684 301476
rect 224908 301412 224972 301476
rect 226748 301472 226812 301476
rect 226748 301416 226762 301472
rect 226762 301416 226812 301472
rect 226748 301412 226812 301416
rect 227668 301412 227732 301476
rect 229692 301412 229756 301476
rect 230612 301472 230676 301476
rect 230612 301416 230626 301472
rect 230626 301416 230676 301472
rect 230612 301412 230676 301416
rect 232084 301472 232148 301476
rect 232084 301416 232134 301472
rect 232134 301416 232148 301472
rect 232084 301412 232148 301416
rect 232268 301412 232332 301476
rect 233188 301412 233252 301476
rect 233556 301412 233620 301476
rect 234844 301472 234908 301476
rect 234844 301416 234858 301472
rect 234858 301416 234908 301472
rect 234844 301412 234908 301416
rect 236684 301472 236748 301476
rect 236684 301416 236698 301472
rect 236698 301416 236748 301472
rect 236684 301412 236748 301416
rect 237788 301412 237852 301476
rect 238524 301412 238588 301476
rect 242940 301412 243004 301476
rect 245516 301412 245580 301476
rect 245884 301548 245948 301612
rect 247724 301412 247788 301476
rect 258396 301412 258460 301476
rect 84700 300732 84764 300796
rect 87460 300732 87524 300796
rect 252876 300596 252940 300660
rect 193260 300052 193324 300116
rect 191972 299508 192036 299572
rect 272564 299432 272628 299436
rect 272564 299376 272578 299432
rect 272578 299376 272628 299432
rect 272564 299372 272628 299376
rect 173020 298828 173084 298892
rect 91508 298692 91572 298756
rect 265756 298692 265820 298756
rect 188292 298148 188356 298212
rect 191420 298072 191484 298076
rect 191420 298016 191470 298072
rect 191470 298016 191484 298072
rect 191420 298012 191484 298016
rect 267780 298012 267844 298076
rect 192708 297332 192772 297396
rect 255268 295836 255332 295900
rect 268332 295292 268396 295356
rect 87092 294476 87156 294540
rect 98316 294476 98380 294540
rect 75684 293932 75748 293996
rect 191972 293116 192036 293180
rect 192708 293116 192772 293180
rect 86540 292572 86604 292636
rect 192708 292572 192772 292636
rect 92980 291892 93044 291956
rect 83964 291756 84028 291820
rect 83964 291212 84028 291276
rect 191604 291272 191668 291276
rect 191604 291216 191618 291272
rect 191618 291216 191668 291272
rect 191604 291212 191668 291216
rect 92612 290396 92676 290460
rect 262444 290668 262508 290732
rect 73292 289988 73356 290052
rect 73476 289852 73540 289916
rect 252876 289444 252940 289508
rect 98500 287268 98564 287332
rect 98684 285636 98748 285700
rect 76420 284820 76484 284884
rect 70164 284276 70228 284340
rect 72924 284276 72988 284340
rect 73108 284200 73172 284204
rect 73108 284144 73158 284200
rect 73158 284144 73172 284200
rect 73108 284140 73172 284144
rect 87092 284140 87156 284204
rect 69980 283460 70044 283524
rect 71636 283460 71700 283524
rect 89484 283460 89548 283524
rect 68692 283324 68756 283388
rect 83412 283384 83476 283388
rect 83412 283328 83462 283384
rect 83462 283328 83476 283384
rect 83412 283324 83476 283328
rect 87092 283188 87156 283252
rect 69980 283052 70044 283116
rect 75684 283052 75748 283116
rect 67404 281556 67468 281620
rect 268332 280876 268396 280940
rect 260972 276796 261036 276860
rect 256740 275572 256804 275636
rect 190316 274620 190380 274684
rect 188844 273260 188908 273324
rect 67404 273124 67468 273188
rect 260052 273124 260116 273188
rect 98684 271084 98748 271148
rect 258396 270540 258460 270604
rect 259500 269316 259564 269380
rect 188292 268500 188356 268564
rect 184060 267140 184124 267204
rect 98868 267004 98932 267068
rect 266860 267064 266924 267068
rect 266860 267008 266874 267064
rect 266874 267008 266924 267064
rect 266860 267004 266924 267008
rect 276244 266732 276308 266796
rect 193444 265508 193508 265572
rect 269068 264828 269132 264892
rect 281580 264148 281644 264212
rect 262444 263604 262508 263668
rect 270724 263604 270788 263668
rect 276244 263604 276308 263668
rect 266492 262652 266556 262716
rect 263548 261700 263612 261764
rect 100892 261488 100956 261492
rect 100892 261432 100906 261488
rect 100906 261432 100956 261488
rect 100892 261428 100956 261432
rect 173020 261428 173084 261492
rect 263732 261292 263796 261356
rect 254532 261020 254596 261084
rect 255268 260612 255332 260676
rect 259500 259796 259564 259860
rect 263732 259524 263796 259588
rect 270724 259584 270788 259588
rect 270724 259528 270738 259584
rect 270738 259528 270788 259584
rect 270724 259524 270788 259528
rect 262260 259388 262324 259452
rect 270540 258844 270604 258908
rect 59124 258164 59188 258228
rect 66116 257892 66180 257956
rect 66668 256864 66732 256868
rect 66668 256808 66682 256864
rect 66682 256808 66732 256864
rect 66668 256804 66732 256808
rect 267964 256804 268028 256868
rect 61884 255852 61948 255916
rect 269252 255172 269316 255236
rect 285628 254492 285692 254556
rect 98132 254356 98196 254420
rect 258396 253676 258460 253740
rect 269068 252588 269132 252652
rect 100708 252452 100772 252516
rect 193260 251772 193324 251836
rect 177252 251228 177316 251292
rect 66484 251152 66548 251156
rect 66484 251096 66498 251152
rect 66498 251096 66548 251152
rect 66484 251092 66548 251096
rect 272564 251092 272628 251156
rect 262076 249732 262140 249796
rect 262444 249732 262508 249796
rect 267780 248372 267844 248436
rect 252876 248100 252940 248164
rect 262812 247828 262876 247892
rect 266308 247828 266372 247892
rect 57836 247148 57900 247212
rect 160692 246196 160756 246260
rect 184244 245652 184308 245716
rect 64644 244428 64708 244492
rect 193260 242796 193324 242860
rect 273300 242796 273364 242860
rect 259684 242252 259748 242316
rect 277164 242252 277228 242316
rect 66300 242116 66364 242180
rect 68692 241708 68756 241772
rect 72740 241768 72804 241772
rect 72740 241712 72754 241768
rect 72754 241712 72804 241768
rect 72740 241708 72804 241712
rect 73292 241768 73356 241772
rect 73292 241712 73306 241768
rect 73306 241712 73356 241768
rect 73292 241708 73356 241712
rect 84700 241708 84764 241772
rect 86724 241708 86788 241772
rect 87092 241768 87156 241772
rect 87092 241712 87142 241768
rect 87142 241712 87156 241768
rect 87092 241708 87156 241712
rect 90956 241708 91020 241772
rect 91508 241768 91572 241772
rect 91508 241712 91558 241768
rect 91558 241712 91572 241768
rect 91508 241708 91572 241712
rect 93900 241708 93964 241772
rect 87460 241572 87524 241636
rect 188292 241572 188356 241636
rect 70348 241496 70412 241500
rect 70348 241440 70362 241496
rect 70362 241440 70412 241496
rect 70348 241436 70412 241440
rect 86540 241496 86604 241500
rect 86540 241440 86590 241496
rect 86590 241440 86604 241496
rect 86540 241436 86604 241440
rect 68876 241300 68940 241364
rect 201540 241496 201604 241500
rect 201540 241440 201590 241496
rect 201590 241440 201604 241496
rect 201540 241436 201604 241440
rect 208348 241496 208412 241500
rect 208348 241440 208398 241496
rect 208398 241440 208412 241496
rect 208348 241436 208412 241440
rect 215156 241496 215220 241500
rect 215156 241440 215206 241496
rect 215206 241440 215220 241496
rect 215156 241436 215220 241440
rect 218652 241496 218716 241500
rect 218652 241440 218666 241496
rect 218666 241440 218716 241496
rect 218652 241436 218716 241440
rect 221228 241436 221292 241500
rect 226196 241436 226260 241500
rect 236500 241436 236564 241500
rect 238892 241436 238956 241500
rect 242756 241436 242820 241500
rect 245516 241436 245580 241500
rect 210372 240892 210436 240956
rect 262076 240756 262140 240820
rect 66300 240212 66364 240276
rect 93900 240212 93964 240276
rect 70900 240076 70964 240140
rect 72740 240076 72804 240140
rect 97764 240076 97828 240140
rect 188844 240076 188908 240140
rect 203012 240076 203076 240140
rect 210556 240076 210620 240140
rect 229692 240076 229756 240140
rect 234844 240076 234908 240140
rect 238892 240076 238956 240140
rect 263732 240076 263796 240140
rect 216444 239940 216508 240004
rect 224172 239804 224236 239868
rect 84700 238716 84764 238780
rect 230244 238716 230308 238780
rect 254532 238580 254596 238644
rect 216444 238036 216508 238100
rect 111564 237900 111628 237964
rect 201540 237900 201604 237964
rect 205404 237900 205468 237964
rect 245700 237900 245764 237964
rect 265756 237900 265820 237964
rect 73108 237492 73172 237556
rect 93716 237492 93780 237556
rect 258396 236676 258460 236740
rect 200620 235724 200684 235788
rect 263548 235724 263612 235788
rect 229876 235588 229940 235652
rect 208348 232460 208412 232524
rect 259500 231780 259564 231844
rect 236684 231100 236748 231164
rect 222700 230284 222764 230348
rect 223436 229876 223500 229940
rect 226564 229740 226628 229804
rect 211660 229060 211724 229124
rect 61884 228924 61948 228988
rect 206140 228380 206204 228444
rect 262260 228380 262324 228444
rect 266492 228244 266556 228308
rect 184060 227700 184124 227764
rect 220676 227700 220740 227764
rect 237604 226884 237668 226948
rect 240732 226884 240796 226948
rect 66116 226340 66180 226404
rect 238524 225660 238588 225724
rect 207060 225524 207124 225588
rect 253060 224708 253124 224772
rect 220860 224164 220924 224228
rect 259684 222940 259748 223004
rect 262812 222804 262876 222868
rect 237788 222668 237852 222732
rect 186820 220084 186884 220148
rect 270724 219268 270788 219332
rect 253060 219132 253124 219196
rect 212580 218044 212644 218108
rect 267780 217908 267844 217972
rect 192708 217228 192772 217292
rect 57836 215868 57900 215932
rect 190316 215868 190380 215932
rect 203012 214644 203076 214708
rect 255268 214508 255332 214572
rect 276244 214508 276308 214572
rect 72740 212468 72804 212532
rect 254532 211924 254596 211988
rect 215892 211788 215956 211852
rect 64644 210292 64708 210356
rect 215340 210292 215404 210356
rect 253060 206212 253124 206276
rect 97212 204988 97276 205052
rect 226748 204852 226812 204916
rect 222332 203492 222396 203556
rect 204300 202132 204364 202196
rect 188844 201376 188908 201380
rect 188844 201320 188894 201376
rect 188894 201320 188908 201376
rect 188844 201316 188908 201320
rect 223620 200636 223684 200700
rect 224908 197916 224972 197980
rect 227668 189620 227732 189684
rect 228220 189620 228284 189684
rect 258396 184180 258460 184244
rect 187556 182820 187620 182884
rect 86724 181324 86788 181388
rect 269068 181324 269132 181388
rect 214420 179964 214484 180028
rect 97948 179420 98012 179484
rect 242940 178604 243004 178668
rect 220492 177380 220556 177444
rect 89484 175884 89548 175948
rect 88932 172484 88996 172548
rect 213684 167588 213748 167652
rect 190316 161604 190380 161668
rect 199332 161664 199396 161668
rect 199332 161608 199382 161664
rect 199382 161608 199396 161664
rect 199332 161604 199396 161608
rect 72924 156496 72988 156500
rect 72924 156440 72938 156496
rect 72938 156440 72988 156496
rect 72924 156436 72988 156440
rect 224908 156164 224972 156228
rect 195836 155212 195900 155276
rect 217548 155212 217612 155276
rect 226380 154532 226444 154596
rect 193812 153036 193876 153100
rect 193812 152628 193876 152692
rect 184244 152356 184308 152420
rect 177252 150996 177316 151060
rect 66668 149092 66732 149156
rect 83412 149092 83476 149156
rect 227668 149228 227732 149292
rect 223620 147732 223684 147796
rect 219204 147052 219268 147116
rect 188292 146916 188356 146980
rect 226932 146236 226996 146300
rect 91508 144740 91572 144804
rect 211660 143788 211724 143852
rect 67772 143516 67836 143580
rect 197860 143108 197924 143172
rect 66116 142700 66180 142764
rect 224724 142156 224788 142220
rect 83412 141476 83476 141540
rect 69980 140116 70044 140180
rect 197860 140524 197924 140588
rect 196572 140388 196636 140452
rect 94820 139572 94884 139636
rect 69980 139436 70044 139500
rect 71636 138756 71700 138820
rect 69428 138348 69492 138412
rect 70164 138212 70228 138276
rect 96292 138076 96356 138140
rect 194180 137668 194244 137732
rect 83412 136716 83476 136780
rect 88932 136716 88996 136780
rect 226932 136308 226996 136372
rect 224724 135900 224788 135964
rect 90956 135492 91020 135556
rect 227668 135492 227732 135556
rect 95188 135356 95252 135420
rect 69244 135220 69308 135284
rect 188844 135084 188908 135148
rect 72372 134676 72436 134740
rect 69428 133452 69492 133516
rect 94820 132092 94884 132156
rect 190316 131140 190380 131204
rect 224908 130596 224972 130660
rect 191420 129236 191484 129300
rect 69244 128420 69308 128484
rect 192708 128420 192772 128484
rect 67772 124340 67836 124404
rect 224356 124068 224420 124132
rect 96292 119988 96356 120052
rect 191604 117948 191668 118012
rect 66116 116996 66180 117060
rect 100892 116588 100956 116652
rect 66484 108564 66548 108628
rect 98500 108292 98564 108356
rect 97948 108020 98012 108084
rect 184060 108020 184124 108084
rect 226564 108624 226628 108628
rect 226564 108568 226614 108624
rect 226614 108568 226628 108624
rect 226564 108564 226628 108568
rect 226380 107748 226444 107812
rect 187556 107476 187620 107540
rect 66668 106932 66732 106996
rect 61884 106252 61948 106316
rect 100708 105844 100772 105908
rect 94820 104076 94884 104140
rect 57836 98092 57900 98156
rect 224724 97412 224788 97476
rect 191052 96868 191116 96932
rect 64644 95372 64708 95436
rect 224908 95100 224972 95164
rect 193444 94692 193508 94756
rect 224356 94692 224420 94756
rect 193812 94148 193876 94212
rect 211660 93392 211724 93396
rect 211660 93336 211710 93392
rect 211710 93336 211724 93392
rect 211660 93332 211724 93336
rect 224724 93392 224788 93396
rect 224724 93336 224774 93392
rect 224774 93336 224788 93392
rect 224724 93332 224788 93336
rect 97212 92788 97276 92852
rect 68876 92652 68940 92716
rect 70900 92652 70964 92716
rect 72372 92652 72436 92716
rect 92244 92652 92308 92716
rect 93716 92652 93780 92716
rect 223436 92924 223500 92988
rect 201540 92848 201604 92852
rect 201540 92792 201590 92848
rect 201590 92792 201604 92848
rect 201540 92788 201604 92792
rect 205404 92848 205468 92852
rect 205404 92792 205454 92848
rect 205454 92792 205468 92848
rect 205404 92788 205468 92792
rect 208348 92848 208412 92852
rect 208348 92792 208398 92848
rect 208398 92792 208412 92848
rect 208348 92788 208412 92792
rect 210004 92848 210068 92852
rect 210004 92792 210054 92848
rect 210054 92792 210068 92848
rect 210004 92788 210068 92792
rect 220676 92788 220740 92852
rect 224356 92788 224420 92852
rect 215340 92652 215404 92716
rect 193444 92516 193508 92580
rect 71636 92380 71700 92444
rect 203012 92380 203076 92444
rect 212580 92380 212644 92444
rect 94820 92108 94884 92172
rect 204852 91972 204916 92036
rect 212580 91972 212644 92036
rect 72740 91020 72804 91084
rect 98500 89388 98564 89452
rect 191052 88028 191116 88092
rect 204852 88028 204916 88092
rect 66484 87892 66548 87956
rect 224908 87892 224972 87956
rect 187740 85444 187804 85508
rect 95188 85308 95252 85372
rect 226380 82588 226444 82652
rect 210004 82452 210068 82516
rect 192708 80684 192772 80748
rect 196572 76468 196636 76532
rect 230612 73748 230676 73812
rect 274588 71708 274652 71772
rect 232084 69532 232148 69596
rect 247724 66132 247788 66196
rect 193812 63412 193876 63476
rect 233188 61372 233252 61436
rect 193812 60556 193876 60620
rect 234660 54436 234724 54500
rect 233556 48860 233620 48924
rect 232268 14452 232332 14516
rect 197860 7516 197924 7580
rect 230428 6156 230492 6220
rect 111564 3436 111628 3500
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 529174 60134 564618
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 59514 493174 60134 528618
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59514 457174 60134 492618
rect 59514 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 60134 457174
rect 59514 456854 60134 456938
rect 59514 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 60134 456854
rect 59514 421174 60134 456618
rect 59514 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 60134 421174
rect 59514 420854 60134 420938
rect 59514 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 60134 420854
rect 59123 405788 59189 405789
rect 59123 405724 59124 405788
rect 59188 405724 59189 405788
rect 59123 405723 59189 405724
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 59126 258229 59186 405723
rect 59514 385174 60134 420618
rect 59514 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 60134 385174
rect 59514 384854 60134 384938
rect 59514 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 60134 384854
rect 59514 349174 60134 384618
rect 59514 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 60134 349174
rect 59514 348854 60134 348938
rect 59514 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 60134 348854
rect 59514 313174 60134 348618
rect 59514 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 60134 313174
rect 59514 312854 60134 312938
rect 59514 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 60134 312854
rect 59514 277174 60134 312618
rect 59514 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 60134 277174
rect 59514 276854 60134 276938
rect 59514 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 60134 276854
rect 59123 258228 59189 258229
rect 59123 258164 59124 258228
rect 59188 258164 59189 258228
rect 59123 258163 59189 258164
rect 57835 247212 57901 247213
rect 57835 247148 57836 247212
rect 57900 247148 57901 247212
rect 57835 247147 57901 247148
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 57838 215933 57898 247147
rect 59514 241174 60134 276618
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 583166 67574 608058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 583166 74414 614898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 75867 585172 75933 585173
rect 75867 585108 75868 585172
rect 75932 585108 75933 585172
rect 75867 585107 75933 585108
rect 75683 581092 75749 581093
rect 75683 581028 75684 581092
rect 75748 581028 75749 581092
rect 75683 581027 75749 581028
rect 70347 580820 70413 580821
rect 70347 580756 70348 580820
rect 70412 580756 70413 580820
rect 70347 580755 70413 580756
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 532894 63854 568338
rect 67771 562052 67837 562053
rect 67771 561988 67772 562052
rect 67836 561988 67837 562052
rect 67771 561987 67837 561988
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 63234 460894 63854 496338
rect 63234 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 63854 460894
rect 63234 460574 63854 460658
rect 63234 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 63854 460574
rect 63234 424894 63854 460338
rect 66954 536614 67574 537166
rect 66954 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 67574 536614
rect 66954 536294 67574 536378
rect 66954 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 67574 536294
rect 66954 500614 67574 536058
rect 66954 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 67574 500614
rect 66954 500294 67574 500378
rect 66954 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 67574 500294
rect 66954 464614 67574 500058
rect 67774 482221 67834 561987
rect 69059 546820 69125 546821
rect 69059 546756 69060 546820
rect 69124 546756 69125 546820
rect 69059 546755 69125 546756
rect 67955 543420 68021 543421
rect 67955 543356 67956 543420
rect 68020 543356 68021 543420
rect 67955 543355 68021 543356
rect 67771 482220 67837 482221
rect 67771 482156 67772 482220
rect 67836 482156 67837 482220
rect 67771 482155 67837 482156
rect 67958 471885 68018 543355
rect 69062 538230 69122 546755
rect 69243 541652 69309 541653
rect 69243 541588 69244 541652
rect 69308 541650 69309 541652
rect 69308 541590 69858 541650
rect 69308 541588 69309 541590
rect 69243 541587 69309 541588
rect 69062 538170 69674 538230
rect 69614 476781 69674 538170
rect 69798 520981 69858 541590
rect 69795 520980 69861 520981
rect 69795 520916 69796 520980
rect 69860 520916 69861 520980
rect 69795 520915 69861 520916
rect 69611 476780 69677 476781
rect 69611 476716 69612 476780
rect 69676 476716 69677 476780
rect 69611 476715 69677 476716
rect 67955 471884 68021 471885
rect 67955 471820 67956 471884
rect 68020 471820 68021 471884
rect 67955 471819 68021 471820
rect 70350 467941 70410 580755
rect 73679 543454 73999 543486
rect 73679 543218 73721 543454
rect 73957 543218 73999 543454
rect 73679 543134 73999 543218
rect 73679 542898 73721 543134
rect 73957 542898 73999 543134
rect 73679 542866 73999 542898
rect 72739 523700 72805 523701
rect 72739 523636 72740 523700
rect 72804 523636 72805 523700
rect 72739 523635 72805 523636
rect 67771 467940 67837 467941
rect 67771 467876 67772 467940
rect 67836 467876 67837 467940
rect 67771 467875 67837 467876
rect 70347 467940 70413 467941
rect 70347 467876 70348 467940
rect 70412 467876 70413 467940
rect 70347 467875 70413 467876
rect 66954 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 67574 464614
rect 66954 464294 67574 464378
rect 66954 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 67574 464294
rect 66954 436356 67574 464058
rect 63234 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 63854 424894
rect 63234 424574 63854 424658
rect 63234 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 63854 424574
rect 63234 388894 63854 424338
rect 67774 409733 67834 467875
rect 67955 440332 68021 440333
rect 67955 440268 67956 440332
rect 68020 440268 68021 440332
rect 67955 440267 68021 440268
rect 67771 409732 67837 409733
rect 67771 409668 67772 409732
rect 67836 409668 67837 409732
rect 67771 409667 67837 409668
rect 66667 398852 66733 398853
rect 66667 398788 66668 398852
rect 66732 398788 66733 398852
rect 66667 398787 66733 398788
rect 63234 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 63854 388894
rect 63234 388574 63854 388658
rect 63234 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 63854 388574
rect 63234 352894 63854 388338
rect 66670 384301 66730 398787
rect 66667 384300 66733 384301
rect 66667 384236 66668 384300
rect 66732 384236 66733 384300
rect 66667 384235 66733 384236
rect 63234 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 63854 352894
rect 63234 352574 63854 352658
rect 63234 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 63854 352574
rect 63234 316894 63854 352338
rect 66954 356614 67574 388356
rect 67774 376685 67834 409667
rect 67958 396405 68018 440267
rect 69427 438972 69493 438973
rect 69427 438908 69428 438972
rect 69492 438908 69493 438972
rect 69427 438907 69493 438908
rect 69430 426189 69490 438907
rect 70163 434620 70229 434621
rect 70163 434556 70164 434620
rect 70228 434556 70229 434620
rect 70163 434555 70229 434556
rect 69427 426188 69493 426189
rect 69427 426124 69428 426188
rect 69492 426124 69493 426188
rect 69427 426123 69493 426124
rect 67955 396404 68021 396405
rect 67955 396340 67956 396404
rect 68020 396340 68021 396404
rect 67955 396339 68021 396340
rect 69611 392052 69677 392053
rect 69611 391988 69612 392052
rect 69676 391988 69677 392052
rect 69611 391987 69677 391988
rect 68875 387836 68941 387837
rect 68875 387772 68876 387836
rect 68940 387772 68941 387836
rect 68875 387771 68941 387772
rect 67771 376684 67837 376685
rect 67771 376620 67772 376684
rect 67836 376620 67837 376684
rect 67771 376619 67837 376620
rect 66954 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 67574 356614
rect 66954 356294 67574 356378
rect 66954 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 67574 356294
rect 66483 322148 66549 322149
rect 66483 322084 66484 322148
rect 66548 322084 66549 322148
rect 66483 322083 66549 322084
rect 63234 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 63854 316894
rect 63234 316574 63854 316658
rect 63234 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 63854 316574
rect 63234 280894 63854 316338
rect 63234 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 63854 280894
rect 63234 280574 63854 280658
rect 63234 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 63854 280574
rect 61883 255916 61949 255917
rect 61883 255852 61884 255916
rect 61948 255852 61949 255916
rect 61883 255851 61949 255852
rect 59514 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 60134 241174
rect 59514 240854 60134 240938
rect 59514 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 60134 240854
rect 57835 215932 57901 215933
rect 57835 215868 57836 215932
rect 57900 215868 57901 215932
rect 57835 215867 57901 215868
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 57838 98157 57898 215867
rect 59514 205174 60134 240618
rect 61886 228989 61946 255851
rect 63234 244894 63854 280338
rect 66115 257956 66181 257957
rect 66115 257892 66116 257956
rect 66180 257892 66181 257956
rect 66115 257891 66181 257892
rect 63234 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 63854 244894
rect 63234 244574 63854 244658
rect 63234 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 63854 244574
rect 64643 244492 64709 244493
rect 64643 244428 64644 244492
rect 64708 244428 64709 244492
rect 64643 244427 64709 244428
rect 61883 228988 61949 228989
rect 61883 228924 61884 228988
rect 61948 228924 61949 228988
rect 61883 228923 61949 228924
rect 59514 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 60134 205174
rect 59514 204854 60134 204938
rect 59514 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 60134 204854
rect 59514 169174 60134 204618
rect 59514 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 60134 169174
rect 59514 168854 60134 168938
rect 59514 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 60134 168854
rect 59514 133174 60134 168618
rect 59514 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 60134 133174
rect 59514 132854 60134 132938
rect 59514 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 60134 132854
rect 57835 98156 57901 98157
rect 57835 98092 57836 98156
rect 57900 98092 57901 98156
rect 57835 98091 57901 98092
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 97174 60134 132618
rect 61886 106317 61946 228923
rect 63234 208894 63854 244338
rect 64646 210357 64706 244427
rect 66118 226405 66178 257891
rect 66486 251157 66546 322083
rect 66954 320614 67574 356058
rect 68878 355333 68938 387771
rect 69614 380901 69674 391987
rect 69611 380900 69677 380901
rect 69611 380836 69612 380900
rect 69676 380836 69677 380900
rect 69611 380835 69677 380836
rect 68875 355332 68941 355333
rect 68875 355268 68876 355332
rect 68940 355268 68941 355332
rect 68875 355267 68941 355268
rect 66954 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 67574 320614
rect 66954 320294 67574 320378
rect 66954 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 67574 320294
rect 66954 285592 67574 320058
rect 68691 283388 68757 283389
rect 68691 283324 68692 283388
rect 68756 283324 68757 283388
rect 68691 283323 68757 283324
rect 67403 281620 67469 281621
rect 67403 281556 67404 281620
rect 67468 281556 67469 281620
rect 67403 281555 67469 281556
rect 67406 273189 67466 281555
rect 67403 273188 67469 273189
rect 67403 273124 67404 273188
rect 67468 273124 67469 273188
rect 67403 273123 67469 273124
rect 66667 256868 66733 256869
rect 66667 256804 66668 256868
rect 66732 256804 66733 256868
rect 66667 256803 66733 256804
rect 66483 251156 66549 251157
rect 66483 251092 66484 251156
rect 66548 251092 66549 251156
rect 66483 251091 66549 251092
rect 66299 242180 66365 242181
rect 66299 242116 66300 242180
rect 66364 242116 66365 242180
rect 66299 242115 66365 242116
rect 66302 240277 66362 242115
rect 66299 240276 66365 240277
rect 66299 240212 66300 240276
rect 66364 240212 66365 240276
rect 66299 240211 66365 240212
rect 66115 226404 66181 226405
rect 66115 226340 66116 226404
rect 66180 226340 66181 226404
rect 66115 226339 66181 226340
rect 64643 210356 64709 210357
rect 64643 210292 64644 210356
rect 64708 210292 64709 210356
rect 64643 210291 64709 210292
rect 63234 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 63854 208894
rect 63234 208574 63854 208658
rect 63234 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 63854 208574
rect 63234 172894 63854 208338
rect 63234 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 63854 172894
rect 63234 172574 63854 172658
rect 63234 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 63854 172574
rect 63234 136894 63854 172338
rect 63234 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 63854 136894
rect 63234 136574 63854 136658
rect 63234 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 63854 136574
rect 61883 106316 61949 106317
rect 61883 106252 61884 106316
rect 61948 106252 61949 106316
rect 61883 106251 61949 106252
rect 59514 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 60134 97174
rect 59514 96854 60134 96938
rect 59514 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 60134 96854
rect 59514 61174 60134 96618
rect 59514 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 60134 61174
rect 59514 60854 60134 60938
rect 59514 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 60134 60854
rect 59514 25174 60134 60618
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 100894 63854 136338
rect 63234 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 63854 100894
rect 63234 100574 63854 100658
rect 63234 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 63854 100574
rect 63234 64894 63854 100338
rect 64646 95437 64706 210291
rect 66670 149157 66730 256803
rect 68694 241773 68754 283323
rect 68691 241772 68757 241773
rect 68691 241708 68692 241772
rect 68756 241708 68757 241772
rect 68691 241707 68757 241708
rect 66954 212614 67574 239592
rect 68694 238770 68754 241707
rect 68878 241365 68938 355267
rect 70166 287070 70226 434555
rect 71635 434484 71701 434485
rect 71635 434420 71636 434484
rect 71700 434420 71701 434484
rect 71635 434419 71701 434420
rect 70347 388244 70413 388245
rect 70347 388180 70348 388244
rect 70412 388180 70413 388244
rect 70347 388179 70413 388180
rect 70350 292590 70410 388179
rect 70350 292530 70594 292590
rect 69982 287010 70226 287070
rect 69982 283525 70042 287010
rect 70163 284340 70229 284341
rect 70163 284276 70164 284340
rect 70228 284276 70229 284340
rect 70163 284275 70229 284276
rect 69979 283524 70045 283525
rect 69979 283460 69980 283524
rect 70044 283460 70045 283524
rect 69979 283459 70045 283460
rect 69979 283116 70045 283117
rect 69979 283052 69980 283116
rect 70044 283052 70045 283116
rect 69979 283051 70045 283052
rect 68875 241364 68941 241365
rect 68875 241300 68876 241364
rect 68940 241300 68941 241364
rect 68875 241299 68941 241300
rect 68694 238710 68938 238770
rect 66954 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 67574 212614
rect 66954 212294 67574 212378
rect 66954 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 67574 212294
rect 66954 176614 67574 212058
rect 66954 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 67574 176614
rect 66954 176294 67574 176378
rect 66954 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 67574 176294
rect 66667 149156 66733 149157
rect 66667 149092 66668 149156
rect 66732 149092 66733 149156
rect 66667 149091 66733 149092
rect 66115 142764 66181 142765
rect 66115 142700 66116 142764
rect 66180 142700 66181 142764
rect 66115 142699 66181 142700
rect 66118 117061 66178 142699
rect 66115 117060 66181 117061
rect 66115 116996 66116 117060
rect 66180 116996 66181 117060
rect 66115 116995 66181 116996
rect 66483 108628 66549 108629
rect 66483 108564 66484 108628
rect 66548 108564 66549 108628
rect 66483 108563 66549 108564
rect 64643 95436 64709 95437
rect 64643 95372 64644 95436
rect 64708 95372 64709 95436
rect 64643 95371 64709 95372
rect 66486 87957 66546 108563
rect 66670 106997 66730 149091
rect 66954 140614 67574 176058
rect 67771 143580 67837 143581
rect 67771 143516 67772 143580
rect 67836 143516 67837 143580
rect 67771 143515 67837 143516
rect 66954 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 67574 140614
rect 66954 140294 67574 140378
rect 66954 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 67574 140294
rect 66954 136782 67574 140058
rect 67774 124405 67834 143515
rect 67771 124404 67837 124405
rect 67771 124340 67772 124404
rect 67836 124340 67837 124404
rect 67771 124339 67837 124340
rect 66667 106996 66733 106997
rect 66667 106932 66668 106996
rect 66732 106932 66733 106996
rect 66667 106931 66733 106932
rect 68878 92717 68938 238710
rect 69982 140181 70042 283051
rect 69979 140180 70045 140181
rect 69979 140116 69980 140180
rect 70044 140116 70045 140180
rect 69979 140115 70045 140116
rect 69982 139501 70042 140115
rect 69979 139500 70045 139501
rect 69979 139436 69980 139500
rect 70044 139436 70045 139500
rect 69979 139435 70045 139436
rect 69427 138412 69493 138413
rect 69427 138348 69428 138412
rect 69492 138348 69493 138412
rect 69427 138347 69493 138348
rect 69243 135284 69309 135285
rect 69243 135220 69244 135284
rect 69308 135220 69309 135284
rect 69243 135219 69309 135220
rect 69246 128485 69306 135219
rect 69430 133517 69490 138347
rect 70166 138277 70226 284275
rect 70534 282930 70594 292530
rect 71638 283525 71698 434419
rect 72555 433804 72621 433805
rect 72555 433740 72556 433804
rect 72620 433740 72621 433804
rect 72555 433739 72621 433740
rect 72558 338197 72618 433739
rect 72742 389061 72802 523635
rect 73794 507454 74414 537166
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73291 478140 73357 478141
rect 73291 478076 73292 478140
rect 73356 478076 73357 478140
rect 73291 478075 73357 478076
rect 73294 441630 73354 478075
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73294 441570 73538 441630
rect 72978 399454 73298 399486
rect 72978 399218 73020 399454
rect 73256 399218 73298 399454
rect 72978 399134 73298 399218
rect 72978 398898 73020 399134
rect 73256 398898 73298 399134
rect 72978 398866 73298 398898
rect 73478 390965 73538 441570
rect 73794 436356 74414 470898
rect 75686 464405 75746 581027
rect 75870 539613 75930 585107
rect 77514 583166 78134 618618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 586894 81854 622338
rect 81234 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 81854 586894
rect 81234 586574 81854 586658
rect 81234 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 81854 586574
rect 81234 583166 81854 586338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 590614 85574 626058
rect 84954 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 85574 590614
rect 84954 590294 85574 590378
rect 84954 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 85574 590294
rect 84954 583166 85574 590058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 583166 92414 596898
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 95514 583166 96134 600618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 80651 581228 80717 581229
rect 80651 581164 80652 581228
rect 80716 581164 80717 581228
rect 80651 581163 80717 581164
rect 79915 580820 79981 580821
rect 79915 580756 79916 580820
rect 79980 580756 79981 580820
rect 79915 580755 79981 580756
rect 77644 561454 77964 561486
rect 77644 561218 77686 561454
rect 77922 561218 77964 561454
rect 77644 561134 77964 561218
rect 77644 560898 77686 561134
rect 77922 560898 77964 561134
rect 77644 560866 77964 560898
rect 75867 539612 75933 539613
rect 75867 539548 75868 539612
rect 75932 539548 75933 539612
rect 75867 539547 75933 539548
rect 75870 475421 75930 539547
rect 77514 511174 78134 537166
rect 79731 534716 79797 534717
rect 79731 534652 79732 534716
rect 79796 534652 79797 534716
rect 79731 534651 79797 534652
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 75867 475420 75933 475421
rect 75867 475356 75868 475420
rect 75932 475356 75933 475420
rect 75867 475355 75933 475356
rect 77514 475174 78134 510618
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 75683 464404 75749 464405
rect 75683 464340 75684 464404
rect 75748 464340 75749 464404
rect 75683 464339 75749 464340
rect 77514 439174 78134 474618
rect 77514 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 78134 439174
rect 77514 438854 78134 438938
rect 77514 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 78134 438854
rect 77514 436356 78134 438618
rect 73659 436252 73725 436253
rect 73659 436188 73660 436252
rect 73724 436188 73725 436252
rect 73659 436187 73725 436188
rect 73662 402990 73722 436187
rect 74579 433668 74645 433669
rect 74579 433604 74580 433668
rect 74644 433604 74645 433668
rect 74579 433603 74645 433604
rect 76419 433668 76485 433669
rect 76419 433604 76420 433668
rect 76484 433604 76485 433668
rect 76419 433603 76485 433604
rect 77339 433668 77405 433669
rect 77339 433604 77340 433668
rect 77404 433604 77405 433668
rect 77339 433603 77405 433604
rect 73662 402930 73906 402990
rect 73475 390964 73541 390965
rect 73475 390900 73476 390964
rect 73540 390900 73541 390964
rect 73475 390899 73541 390900
rect 73846 389190 73906 402930
rect 73478 389130 73906 389190
rect 72739 389060 72805 389061
rect 72739 388996 72740 389060
rect 72804 388996 72805 389060
rect 72739 388995 72805 388996
rect 72739 356692 72805 356693
rect 72739 356628 72740 356692
rect 72804 356628 72805 356692
rect 72739 356627 72805 356628
rect 72555 338196 72621 338197
rect 72555 338132 72556 338196
rect 72620 338132 72621 338196
rect 72555 338131 72621 338132
rect 71635 283524 71701 283525
rect 71635 283460 71636 283524
rect 71700 283460 71701 283524
rect 71635 283459 71701 283460
rect 70350 282870 70594 282930
rect 70350 241501 70410 282870
rect 72742 241773 72802 356627
rect 73291 290052 73357 290053
rect 73291 289988 73292 290052
rect 73356 289988 73357 290052
rect 73291 289987 73357 289988
rect 72923 284340 72989 284341
rect 72923 284276 72924 284340
rect 72988 284276 72989 284340
rect 72923 284275 72989 284276
rect 72739 241772 72805 241773
rect 72739 241708 72740 241772
rect 72804 241708 72805 241772
rect 72739 241707 72805 241708
rect 70347 241500 70413 241501
rect 70347 241436 70348 241500
rect 70412 241436 70413 241500
rect 70347 241435 70413 241436
rect 70899 240140 70965 240141
rect 70899 240076 70900 240140
rect 70964 240076 70965 240140
rect 70899 240075 70965 240076
rect 72739 240140 72805 240141
rect 72739 240076 72740 240140
rect 72804 240076 72805 240140
rect 72739 240075 72805 240076
rect 70163 138276 70229 138277
rect 70163 138212 70164 138276
rect 70228 138212 70229 138276
rect 70163 138211 70229 138212
rect 69427 133516 69493 133517
rect 69427 133452 69428 133516
rect 69492 133452 69493 133516
rect 69427 133451 69493 133452
rect 69243 128484 69309 128485
rect 69243 128420 69244 128484
rect 69308 128420 69309 128484
rect 69243 128419 69309 128420
rect 70902 92717 70962 240075
rect 72742 212533 72802 240075
rect 72739 212532 72805 212533
rect 72739 212468 72740 212532
rect 72804 212468 72805 212532
rect 72739 212467 72805 212468
rect 71635 138820 71701 138821
rect 71635 138756 71636 138820
rect 71700 138756 71701 138820
rect 71635 138755 71701 138756
rect 68875 92716 68941 92717
rect 68875 92652 68876 92716
rect 68940 92652 68941 92716
rect 68875 92651 68941 92652
rect 70899 92716 70965 92717
rect 70899 92652 70900 92716
rect 70964 92652 70965 92716
rect 70899 92651 70965 92652
rect 71638 92445 71698 138755
rect 72371 134740 72437 134741
rect 72371 134676 72372 134740
rect 72436 134676 72437 134740
rect 72371 134675 72437 134676
rect 72374 92717 72434 134675
rect 72371 92716 72437 92717
rect 72371 92652 72372 92716
rect 72436 92652 72437 92716
rect 72371 92651 72437 92652
rect 71635 92444 71701 92445
rect 71635 92380 71636 92444
rect 71700 92380 71701 92444
rect 71635 92379 71701 92380
rect 72742 91085 72802 212467
rect 72926 156501 72986 284275
rect 73107 284204 73173 284205
rect 73107 284140 73108 284204
rect 73172 284140 73173 284204
rect 73107 284139 73173 284140
rect 73110 237557 73170 284139
rect 73294 241773 73354 289987
rect 73478 289917 73538 389130
rect 73794 363454 74414 388356
rect 74582 383757 74642 433603
rect 74579 383756 74645 383757
rect 74579 383692 74580 383756
rect 74644 383692 74645 383756
rect 74579 383691 74645 383692
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 75683 293996 75749 293997
rect 75683 293932 75684 293996
rect 75748 293932 75749 293996
rect 75683 293931 75749 293932
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73475 289916 73541 289917
rect 73475 289852 73476 289916
rect 73540 289852 73541 289916
rect 73475 289851 73541 289852
rect 73794 285592 74414 290898
rect 75686 283117 75746 293931
rect 76422 284885 76482 433603
rect 77342 326365 77402 433603
rect 79734 389061 79794 534651
rect 79918 435570 79978 580755
rect 80654 456109 80714 581163
rect 83963 580820 84029 580821
rect 83963 580756 83964 580820
rect 84028 580756 84029 580820
rect 83963 580755 84029 580756
rect 88931 580820 88997 580821
rect 88931 580756 88932 580820
rect 88996 580756 88997 580820
rect 88931 580755 88997 580756
rect 92611 580820 92677 580821
rect 92611 580756 92612 580820
rect 92676 580756 92677 580820
rect 92611 580755 92677 580756
rect 81609 543454 81929 543486
rect 81609 543218 81651 543454
rect 81887 543218 81929 543454
rect 81609 543134 81929 543218
rect 81609 542898 81651 543134
rect 81887 542898 81929 543134
rect 81609 542866 81929 542898
rect 81234 514894 81854 537166
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 81234 478894 81854 514338
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 80651 456108 80717 456109
rect 80651 456044 80652 456108
rect 80716 456044 80717 456108
rect 80651 456043 80717 456044
rect 81234 442894 81854 478338
rect 81234 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 81854 442894
rect 81234 442574 81854 442658
rect 81234 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 81854 442574
rect 81234 436356 81854 442338
rect 83966 437477 84026 580755
rect 85575 561454 85895 561486
rect 85575 561218 85617 561454
rect 85853 561218 85895 561454
rect 85575 561134 85895 561218
rect 85575 560898 85617 561134
rect 85853 560898 85895 561134
rect 85575 560866 85895 560898
rect 84954 518614 85574 537166
rect 88747 520980 88813 520981
rect 88747 520916 88748 520980
rect 88812 520916 88813 520980
rect 88747 520915 88813 520916
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 84954 482614 85574 518058
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 84954 446614 85574 482058
rect 84954 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 85574 446614
rect 84954 446294 85574 446378
rect 84954 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 85574 446294
rect 82123 437476 82189 437477
rect 82123 437412 82124 437476
rect 82188 437412 82189 437476
rect 82123 437411 82189 437412
rect 83963 437476 84029 437477
rect 83963 437412 83964 437476
rect 84028 437412 84029 437476
rect 83963 437411 84029 437412
rect 79918 435510 80162 435570
rect 80102 389061 80162 435510
rect 81939 433668 82005 433669
rect 81939 433604 81940 433668
rect 82004 433604 82005 433668
rect 81939 433603 82005 433604
rect 79731 389060 79797 389061
rect 79731 388996 79732 389060
rect 79796 388996 79797 389060
rect 79731 388995 79797 388996
rect 80099 389060 80165 389061
rect 80099 388996 80100 389060
rect 80164 388996 80165 389060
rect 80099 388995 80165 388996
rect 77514 367174 78134 388356
rect 77514 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 78134 367174
rect 77514 366854 78134 366938
rect 77514 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 78134 366854
rect 77514 331174 78134 366618
rect 77514 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 78134 331174
rect 77514 330854 78134 330938
rect 77514 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 78134 330854
rect 77339 326364 77405 326365
rect 77339 326300 77340 326364
rect 77404 326300 77405 326364
rect 77339 326299 77405 326300
rect 77514 295174 78134 330618
rect 77514 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 78134 295174
rect 77514 294854 78134 294938
rect 77514 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 78134 294854
rect 77514 285592 78134 294618
rect 81234 370894 81854 388356
rect 81234 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 81854 370894
rect 81234 370574 81854 370658
rect 81234 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 81854 370574
rect 81234 334894 81854 370338
rect 81234 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 81854 334894
rect 81234 334574 81854 334658
rect 81234 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 81854 334574
rect 81234 298894 81854 334338
rect 81942 317525 82002 433603
rect 82126 390693 82186 437411
rect 84954 436356 85574 446058
rect 83963 436252 84029 436253
rect 83963 436188 83964 436252
rect 84028 436188 84029 436252
rect 83963 436187 84029 436188
rect 82123 390692 82189 390693
rect 82123 390628 82124 390692
rect 82188 390628 82189 390692
rect 82123 390627 82189 390628
rect 81939 317524 82005 317525
rect 81939 317460 81940 317524
rect 82004 317460 82005 317524
rect 81939 317459 82005 317460
rect 81942 305013 82002 317459
rect 81939 305012 82005 305013
rect 81939 304948 81940 305012
rect 82004 304948 82005 305012
rect 81939 304947 82005 304948
rect 81234 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 81854 298894
rect 81234 298574 81854 298658
rect 81234 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 81854 298574
rect 81234 285592 81854 298338
rect 83966 291821 84026 436187
rect 84699 433668 84765 433669
rect 84699 433604 84700 433668
rect 84764 433604 84765 433668
rect 84699 433603 84765 433604
rect 85803 433668 85869 433669
rect 85803 433604 85804 433668
rect 85868 433604 85869 433668
rect 85803 433603 85869 433604
rect 87091 433668 87157 433669
rect 87091 433604 87092 433668
rect 87156 433604 87157 433668
rect 87091 433603 87157 433604
rect 87459 433668 87525 433669
rect 87459 433604 87460 433668
rect 87524 433604 87525 433668
rect 87459 433603 87525 433604
rect 84702 318749 84762 433603
rect 84954 374614 85574 388356
rect 84954 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 85574 374614
rect 84954 374294 85574 374378
rect 84954 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 85574 374294
rect 84954 338614 85574 374058
rect 84954 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 85574 338614
rect 84954 338294 85574 338378
rect 84954 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 85574 338294
rect 84699 318748 84765 318749
rect 84699 318684 84700 318748
rect 84764 318684 84765 318748
rect 84699 318683 84765 318684
rect 84954 302614 85574 338058
rect 85806 320245 85866 433603
rect 86723 387020 86789 387021
rect 86723 386956 86724 387020
rect 86788 386956 86789 387020
rect 86723 386955 86789 386956
rect 85803 320244 85869 320245
rect 85803 320180 85804 320244
rect 85868 320180 85869 320244
rect 85803 320179 85869 320180
rect 84954 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 85574 302614
rect 84954 302294 85574 302378
rect 84954 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 85574 302294
rect 84699 300796 84765 300797
rect 84699 300732 84700 300796
rect 84764 300732 84765 300796
rect 84699 300731 84765 300732
rect 83963 291820 84029 291821
rect 83963 291756 83964 291820
rect 84028 291756 84029 291820
rect 83963 291755 84029 291756
rect 83966 291277 84026 291755
rect 83963 291276 84029 291277
rect 83963 291212 83964 291276
rect 84028 291212 84029 291276
rect 83963 291211 84029 291212
rect 76419 284884 76485 284885
rect 76419 284820 76420 284884
rect 76484 284820 76485 284884
rect 76419 284819 76485 284820
rect 83411 283388 83477 283389
rect 83411 283324 83412 283388
rect 83476 283324 83477 283388
rect 83411 283323 83477 283324
rect 75683 283116 75749 283117
rect 75683 283052 75684 283116
rect 75748 283052 75749 283116
rect 75683 283051 75749 283052
rect 78977 273454 79297 273486
rect 78977 273218 79019 273454
rect 79255 273218 79297 273454
rect 78977 273134 79297 273218
rect 78977 272898 79019 273134
rect 79255 272898 79297 273134
rect 78977 272866 79297 272898
rect 74345 255454 74665 255486
rect 74345 255218 74387 255454
rect 74623 255218 74665 255454
rect 74345 255134 74665 255218
rect 74345 254898 74387 255134
rect 74623 254898 74665 255134
rect 74345 254866 74665 254898
rect 73291 241772 73357 241773
rect 73291 241708 73292 241772
rect 73356 241708 73357 241772
rect 73291 241707 73357 241708
rect 73107 237556 73173 237557
rect 73107 237492 73108 237556
rect 73172 237492 73173 237556
rect 73107 237491 73173 237492
rect 73794 219454 74414 239592
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 72923 156500 72989 156501
rect 72923 156436 72924 156500
rect 72988 156436 72989 156500
rect 72923 156435 72989 156436
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 136782 74414 146898
rect 77514 223174 78134 239592
rect 77514 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 78134 223174
rect 77514 222854 78134 222938
rect 77514 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 78134 222854
rect 77514 187174 78134 222618
rect 77514 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 78134 187174
rect 77514 186854 78134 186938
rect 77514 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 78134 186854
rect 77514 151174 78134 186618
rect 77514 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 78134 151174
rect 77514 150854 78134 150938
rect 77514 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 78134 150854
rect 77514 136782 78134 150618
rect 81234 226894 81854 239592
rect 81234 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 81854 226894
rect 81234 226574 81854 226658
rect 81234 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 81854 226574
rect 81234 190894 81854 226338
rect 81234 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 81854 190894
rect 81234 190574 81854 190658
rect 81234 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 81854 190574
rect 81234 154894 81854 190338
rect 81234 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 81854 154894
rect 81234 154574 81854 154658
rect 81234 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 81854 154574
rect 81234 136782 81854 154338
rect 83414 149157 83474 283323
rect 83609 255454 83929 255486
rect 83609 255218 83651 255454
rect 83887 255218 83929 255454
rect 83609 255134 83929 255218
rect 83609 254898 83651 255134
rect 83887 254898 83929 255134
rect 83609 254866 83929 254898
rect 84702 241773 84762 300731
rect 84954 285592 85574 302058
rect 86539 292636 86605 292637
rect 86539 292572 86540 292636
rect 86604 292572 86605 292636
rect 86539 292571 86605 292572
rect 84699 241772 84765 241773
rect 84699 241708 84700 241772
rect 84764 241708 84765 241772
rect 84699 241707 84765 241708
rect 84702 238781 84762 241707
rect 86542 241501 86602 292571
rect 86726 241773 86786 386955
rect 87094 294541 87154 433603
rect 87462 382941 87522 433603
rect 88338 417454 88658 417486
rect 88338 417218 88380 417454
rect 88616 417218 88658 417454
rect 88338 417134 88658 417218
rect 88338 416898 88380 417134
rect 88616 416898 88658 417134
rect 88338 416866 88658 416898
rect 88750 390557 88810 520915
rect 88934 438837 88994 580755
rect 89540 543454 89860 543486
rect 89540 543218 89582 543454
rect 89818 543218 89860 543454
rect 89540 543134 89860 543218
rect 89540 542898 89582 543134
rect 89818 542898 89860 543134
rect 89540 542866 89860 542898
rect 91794 525454 92414 537166
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91323 482220 91389 482221
rect 91323 482156 91324 482220
rect 91388 482156 91389 482220
rect 91323 482155 91389 482156
rect 88931 438836 88997 438837
rect 88931 438772 88932 438836
rect 88996 438772 88997 438836
rect 88931 438771 88997 438772
rect 88934 438293 88994 438771
rect 88931 438292 88997 438293
rect 88931 438228 88932 438292
rect 88996 438228 88997 438292
rect 88931 438227 88997 438228
rect 90219 433804 90285 433805
rect 90219 433740 90220 433804
rect 90284 433740 90285 433804
rect 90219 433739 90285 433740
rect 88747 390556 88813 390557
rect 88747 390492 88748 390556
rect 88812 390492 88813 390556
rect 88747 390491 88813 390492
rect 87459 382940 87525 382941
rect 87459 382876 87460 382940
rect 87524 382876 87525 382940
rect 87459 382875 87525 382876
rect 90222 316845 90282 433739
rect 91139 433668 91205 433669
rect 91139 433604 91140 433668
rect 91204 433604 91205 433668
rect 91139 433603 91205 433604
rect 90219 316844 90285 316845
rect 90219 316780 90220 316844
rect 90284 316780 90285 316844
rect 90219 316779 90285 316780
rect 91142 305149 91202 433603
rect 91326 390421 91386 482155
rect 91794 453454 92414 488898
rect 92614 478141 92674 580755
rect 99234 568894 99854 604338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 101259 581092 101325 581093
rect 101259 581028 101260 581092
rect 101324 581028 101325 581092
rect 101259 581027 101325 581028
rect 99234 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 99854 568894
rect 99234 568574 99854 568658
rect 99234 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 99854 568574
rect 96659 554164 96725 554165
rect 96659 554100 96660 554164
rect 96724 554100 96725 554164
rect 96659 554099 96725 554100
rect 95514 529174 96134 537166
rect 95514 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 96134 529174
rect 95514 528854 96134 528938
rect 95514 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 96134 528854
rect 95514 493174 96134 528618
rect 95514 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 96134 493174
rect 95514 492854 96134 492938
rect 95514 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 96134 492854
rect 92611 478140 92677 478141
rect 92611 478076 92612 478140
rect 92676 478076 92677 478140
rect 92611 478075 92677 478076
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 436356 92414 452898
rect 95514 457174 96134 492618
rect 95514 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 96134 457174
rect 95514 456854 96134 456938
rect 95514 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 96134 456854
rect 95003 436524 95069 436525
rect 95003 436460 95004 436524
rect 95068 436460 95069 436524
rect 95003 436459 95069 436460
rect 92979 434620 93045 434621
rect 92979 434556 92980 434620
rect 93044 434556 93045 434620
rect 92979 434555 93045 434556
rect 92611 433668 92677 433669
rect 92611 433604 92612 433668
rect 92676 433604 92677 433668
rect 92611 433603 92677 433604
rect 91323 390420 91389 390421
rect 91323 390356 91324 390420
rect 91388 390356 91389 390420
rect 91323 390355 91389 390356
rect 91794 381454 92414 388356
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91139 305148 91205 305149
rect 91139 305084 91140 305148
rect 91204 305084 91205 305148
rect 91139 305083 91205 305084
rect 90955 305012 91021 305013
rect 90955 304948 90956 305012
rect 91020 304948 91021 305012
rect 90955 304947 91021 304948
rect 87459 300796 87525 300797
rect 87459 300732 87460 300796
rect 87524 300732 87525 300796
rect 87459 300731 87525 300732
rect 87091 294540 87157 294541
rect 87091 294476 87092 294540
rect 87156 294476 87157 294540
rect 87091 294475 87157 294476
rect 87091 284204 87157 284205
rect 87091 284140 87092 284204
rect 87156 284140 87157 284204
rect 87091 284139 87157 284140
rect 87094 283253 87154 284139
rect 87091 283252 87157 283253
rect 87091 283188 87092 283252
rect 87156 283188 87157 283252
rect 87091 283187 87157 283188
rect 87094 241773 87154 283187
rect 86723 241772 86789 241773
rect 86723 241708 86724 241772
rect 86788 241708 86789 241772
rect 86723 241707 86789 241708
rect 87091 241772 87157 241773
rect 87091 241708 87092 241772
rect 87156 241708 87157 241772
rect 87091 241707 87157 241708
rect 86539 241500 86605 241501
rect 86539 241436 86540 241500
rect 86604 241436 86605 241500
rect 86539 241435 86605 241436
rect 84699 238780 84765 238781
rect 84699 238716 84700 238780
rect 84764 238716 84765 238780
rect 84699 238715 84765 238716
rect 84954 230614 85574 239592
rect 84954 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 85574 230614
rect 84954 230294 85574 230378
rect 84954 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 85574 230294
rect 84954 194614 85574 230058
rect 84954 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 85574 194614
rect 84954 194294 85574 194378
rect 84954 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 85574 194294
rect 84954 158614 85574 194058
rect 86726 181389 86786 241707
rect 87462 241637 87522 300731
rect 89483 283524 89549 283525
rect 89483 283460 89484 283524
rect 89548 283460 89549 283524
rect 89483 283459 89549 283460
rect 88241 273454 88561 273486
rect 88241 273218 88283 273454
rect 88519 273218 88561 273454
rect 88241 273134 88561 273218
rect 88241 272898 88283 273134
rect 88519 272898 88561 273134
rect 88241 272866 88561 272898
rect 87459 241636 87525 241637
rect 87459 241572 87460 241636
rect 87524 241572 87525 241636
rect 87459 241571 87525 241572
rect 86723 181388 86789 181389
rect 86723 181324 86724 181388
rect 86788 181324 86789 181388
rect 86723 181323 86789 181324
rect 89486 175949 89546 283459
rect 90958 241773 91018 304947
rect 91142 301477 91202 305083
rect 91139 301476 91205 301477
rect 91139 301412 91140 301476
rect 91204 301412 91205 301476
rect 91139 301411 91205 301412
rect 91507 298756 91573 298757
rect 91507 298692 91508 298756
rect 91572 298692 91573 298756
rect 91507 298691 91573 298692
rect 91510 241773 91570 298691
rect 91794 285592 92414 308898
rect 92614 290461 92674 433603
rect 92982 291957 93042 434555
rect 94451 433804 94517 433805
rect 94451 433740 94452 433804
rect 94516 433740 94517 433804
rect 94451 433739 94517 433740
rect 93899 387972 93965 387973
rect 93899 387908 93900 387972
rect 93964 387908 93965 387972
rect 93899 387907 93965 387908
rect 92979 291956 93045 291957
rect 92979 291892 92980 291956
rect 93044 291892 93045 291956
rect 92979 291891 93045 291892
rect 92611 290460 92677 290461
rect 92611 290396 92612 290460
rect 92676 290396 92677 290460
rect 92611 290395 92677 290396
rect 92873 255454 93193 255486
rect 92873 255218 92915 255454
rect 93151 255218 93193 255454
rect 92873 255134 93193 255218
rect 92873 254898 92915 255134
rect 93151 254898 93193 255134
rect 92873 254866 93193 254898
rect 93902 241773 93962 387907
rect 94454 320789 94514 433739
rect 95006 388245 95066 436459
rect 95514 436356 96134 456618
rect 96662 456109 96722 554099
rect 96843 547092 96909 547093
rect 96843 547028 96844 547092
rect 96908 547028 96909 547092
rect 96843 547027 96909 547028
rect 96846 537437 96906 547027
rect 96843 537436 96909 537437
rect 96843 537372 96844 537436
rect 96908 537372 96909 537436
rect 96843 537371 96909 537372
rect 99234 532894 99854 568338
rect 100707 549404 100773 549405
rect 100707 549340 100708 549404
rect 100772 549340 100773 549404
rect 100707 549339 100773 549340
rect 99234 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 99854 532894
rect 99234 532574 99854 532658
rect 99234 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 99854 532574
rect 99234 496894 99854 532338
rect 99234 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 99854 496894
rect 99234 496574 99854 496658
rect 99234 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 99854 496574
rect 96843 474060 96909 474061
rect 96843 473996 96844 474060
rect 96908 473996 96909 474060
rect 96843 473995 96909 473996
rect 96659 456108 96725 456109
rect 96659 456044 96660 456108
rect 96724 456044 96725 456108
rect 96659 456043 96725 456044
rect 96659 455972 96725 455973
rect 96659 455908 96660 455972
rect 96724 455908 96725 455972
rect 96659 455907 96725 455908
rect 96475 446452 96541 446453
rect 96475 446388 96476 446452
rect 96540 446388 96541 446452
rect 96475 446387 96541 446388
rect 96291 436388 96357 436389
rect 96291 436324 96292 436388
rect 96356 436324 96357 436388
rect 96291 436323 96357 436324
rect 95003 388244 95069 388245
rect 95003 388180 95004 388244
rect 95068 388180 95069 388244
rect 95003 388179 95069 388180
rect 95514 385174 96134 388356
rect 95514 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 96134 385174
rect 95514 384854 96134 384938
rect 95514 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 96134 384854
rect 95514 349174 96134 384618
rect 96294 383757 96354 436323
rect 96478 433669 96538 446387
rect 96475 433668 96541 433669
rect 96475 433604 96476 433668
rect 96540 433604 96541 433668
rect 96475 433603 96541 433604
rect 96478 390693 96538 433603
rect 96662 390693 96722 455907
rect 96475 390692 96541 390693
rect 96475 390628 96476 390692
rect 96540 390628 96541 390692
rect 96475 390627 96541 390628
rect 96659 390692 96725 390693
rect 96659 390628 96660 390692
rect 96724 390628 96725 390692
rect 96659 390627 96725 390628
rect 96846 390421 96906 473995
rect 99234 460894 99854 496338
rect 99234 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 99854 460894
rect 99234 460574 99854 460658
rect 99234 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 99854 460574
rect 99234 436356 99854 460338
rect 99971 433804 100037 433805
rect 99971 433740 99972 433804
rect 100036 433740 100037 433804
rect 99971 433739 100037 433740
rect 98131 433668 98197 433669
rect 98131 433604 98132 433668
rect 98196 433604 98197 433668
rect 98131 433603 98197 433604
rect 98315 433668 98381 433669
rect 98315 433604 98316 433668
rect 98380 433604 98381 433668
rect 98315 433603 98381 433604
rect 96843 390420 96909 390421
rect 96843 390356 96844 390420
rect 96908 390356 96909 390420
rect 96843 390355 96909 390356
rect 96291 383756 96357 383757
rect 96291 383692 96292 383756
rect 96356 383692 96357 383756
rect 96291 383691 96357 383692
rect 95514 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 96134 349174
rect 95514 348854 96134 348938
rect 95514 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 96134 348854
rect 94451 320788 94517 320789
rect 94451 320724 94452 320788
rect 94516 320724 94517 320788
rect 94451 320723 94517 320724
rect 95514 313174 96134 348618
rect 98134 319429 98194 433603
rect 98131 319428 98197 319429
rect 98131 319364 98132 319428
rect 98196 319364 98197 319428
rect 98131 319363 98197 319364
rect 95514 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 96134 313174
rect 95514 312854 96134 312938
rect 95514 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 96134 312854
rect 95514 285592 96134 312618
rect 98318 294541 98378 433603
rect 99234 352894 99854 388356
rect 99234 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 99854 352894
rect 99234 352574 99854 352658
rect 99234 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 99854 352574
rect 99234 316894 99854 352338
rect 99234 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 99854 316894
rect 99234 316574 99854 316658
rect 99234 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 99854 316574
rect 98315 294540 98381 294541
rect 98315 294476 98316 294540
rect 98380 294476 98381 294540
rect 98315 294475 98381 294476
rect 98499 287332 98565 287333
rect 98499 287268 98500 287332
rect 98564 287268 98565 287332
rect 98499 287267 98565 287268
rect 98502 267750 98562 287267
rect 98683 285700 98749 285701
rect 98683 285636 98684 285700
rect 98748 285636 98749 285700
rect 98683 285635 98749 285636
rect 98686 271149 98746 285635
rect 99234 285592 99854 316338
rect 99974 302837 100034 433739
rect 100155 433668 100221 433669
rect 100155 433604 100156 433668
rect 100220 433604 100221 433668
rect 100155 433603 100221 433604
rect 100158 388517 100218 433603
rect 100710 390557 100770 549339
rect 101262 460950 101322 581027
rect 102954 572614 103574 608058
rect 102954 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 103574 572614
rect 102954 572294 103574 572378
rect 102954 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 103574 572294
rect 102954 536614 103574 572058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 104939 565860 105005 565861
rect 104939 565796 104940 565860
rect 105004 565796 105005 565860
rect 104939 565795 105005 565796
rect 102954 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 103574 536614
rect 102954 536294 103574 536378
rect 102954 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 103574 536294
rect 102954 500614 103574 536058
rect 102954 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 103574 500614
rect 102954 500294 103574 500378
rect 102954 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 103574 500294
rect 102954 464614 103574 500058
rect 104203 476780 104269 476781
rect 104203 476716 104204 476780
rect 104268 476716 104269 476780
rect 104203 476715 104269 476716
rect 102954 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 103574 464614
rect 102954 464294 103574 464378
rect 102954 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 103574 464294
rect 101262 460890 102058 460950
rect 101998 459645 102058 460890
rect 101995 459644 102061 459645
rect 101995 459580 101996 459644
rect 102060 459580 102061 459644
rect 101995 459579 102061 459580
rect 101998 438157 102058 459579
rect 101995 438156 102061 438157
rect 101995 438092 101996 438156
rect 102060 438092 102061 438156
rect 101995 438091 102061 438092
rect 102954 436356 103574 464058
rect 102731 436116 102797 436117
rect 102731 436052 102732 436116
rect 102796 436052 102797 436116
rect 102731 436051 102797 436052
rect 102547 433668 102613 433669
rect 102547 433604 102548 433668
rect 102612 433604 102613 433668
rect 102547 433603 102613 433604
rect 100707 390556 100773 390557
rect 100707 390492 100708 390556
rect 100772 390492 100773 390556
rect 100707 390491 100773 390492
rect 102550 388517 102610 433603
rect 100155 388516 100221 388517
rect 100155 388452 100156 388516
rect 100220 388452 100221 388516
rect 100155 388451 100221 388452
rect 102547 388516 102613 388517
rect 102547 388452 102548 388516
rect 102612 388452 102613 388516
rect 102547 388451 102613 388452
rect 102734 320245 102794 436051
rect 103698 399454 104018 399486
rect 103698 399218 103740 399454
rect 103976 399218 104018 399454
rect 103698 399134 104018 399218
rect 103698 398898 103740 399134
rect 103976 398898 104018 399134
rect 103698 398866 104018 398898
rect 104206 390693 104266 476715
rect 104203 390692 104269 390693
rect 104203 390628 104204 390692
rect 104268 390628 104269 390692
rect 104203 390627 104269 390628
rect 104942 390557 105002 565795
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 105123 535532 105189 535533
rect 105123 535468 105124 535532
rect 105188 535468 105189 535532
rect 105123 535467 105189 535468
rect 105126 390693 105186 535467
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 113514 547174 114134 582618
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 113514 511174 114134 546618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117234 550894 117854 586338
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 114507 522340 114573 522341
rect 114507 522276 114508 522340
rect 114572 522276 114573 522340
rect 114507 522275 114573 522276
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 113514 475174 114134 510618
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 111931 472564 111997 472565
rect 111931 472500 111932 472564
rect 111996 472500 111997 472564
rect 111931 472499 111997 472500
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 107699 440876 107765 440877
rect 107699 440812 107700 440876
rect 107764 440812 107765 440876
rect 107699 440811 107765 440812
rect 106411 433668 106477 433669
rect 106411 433604 106412 433668
rect 106476 433604 106477 433668
rect 106411 433603 106477 433604
rect 105123 390692 105189 390693
rect 105123 390628 105124 390692
rect 105188 390628 105189 390692
rect 105123 390627 105189 390628
rect 104939 390556 105005 390557
rect 104939 390492 104940 390556
rect 105004 390492 105005 390556
rect 104939 390491 105005 390492
rect 102954 356614 103574 388356
rect 102954 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 103574 356614
rect 102954 356294 103574 356378
rect 102954 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 103574 356294
rect 102954 320614 103574 356058
rect 102954 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 103574 320614
rect 102954 320294 103574 320378
rect 102731 320244 102797 320245
rect 102731 320180 102732 320244
rect 102796 320180 102797 320244
rect 102731 320179 102797 320180
rect 102954 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 103574 320294
rect 99971 302836 100037 302837
rect 99971 302772 99972 302836
rect 100036 302772 100037 302836
rect 99971 302771 100037 302772
rect 102954 284614 103574 320058
rect 106414 318069 106474 433603
rect 107702 390693 107762 440811
rect 109794 436356 110414 470898
rect 108987 433668 109053 433669
rect 108987 433604 108988 433668
rect 109052 433604 109053 433668
rect 108987 433603 109053 433604
rect 110643 433668 110709 433669
rect 110643 433604 110644 433668
rect 110708 433604 110709 433668
rect 110643 433603 110709 433604
rect 111747 433668 111813 433669
rect 111747 433604 111748 433668
rect 111812 433604 111813 433668
rect 111747 433603 111813 433604
rect 108990 433530 109050 433603
rect 108806 433470 109050 433530
rect 108806 427830 108866 433470
rect 108806 427770 109050 427830
rect 108990 398850 109050 427770
rect 108806 398790 109050 398850
rect 107699 390692 107765 390693
rect 107699 390628 107700 390692
rect 107764 390628 107765 390692
rect 107699 390627 107765 390628
rect 108806 389190 108866 398790
rect 108806 389130 109050 389190
rect 106411 318068 106477 318069
rect 106411 318004 106412 318068
rect 106476 318004 106477 318068
rect 106411 318003 106477 318004
rect 108990 305693 109050 389130
rect 109794 363454 110414 388356
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 108987 305692 109053 305693
rect 108987 305628 108988 305692
rect 109052 305628 109053 305692
rect 108987 305627 109053 305628
rect 102954 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 103574 284614
rect 102954 284294 103574 284378
rect 102954 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 103574 284294
rect 98683 271148 98749 271149
rect 98683 271084 98684 271148
rect 98748 271084 98749 271148
rect 98683 271083 98749 271084
rect 98502 267690 98930 267750
rect 98870 267069 98930 267690
rect 98867 267068 98933 267069
rect 98867 267004 98868 267068
rect 98932 267004 98933 267068
rect 98867 267003 98933 267004
rect 100891 261492 100957 261493
rect 100891 261428 100892 261492
rect 100956 261428 100957 261492
rect 100891 261427 100957 261428
rect 98131 254420 98197 254421
rect 98131 254356 98132 254420
rect 98196 254356 98197 254420
rect 98131 254355 98197 254356
rect 90955 241772 91021 241773
rect 90955 241708 90956 241772
rect 91020 241708 91021 241772
rect 90955 241707 91021 241708
rect 91507 241772 91573 241773
rect 91507 241708 91508 241772
rect 91572 241708 91573 241772
rect 91507 241707 91573 241708
rect 93899 241772 93965 241773
rect 93899 241708 93900 241772
rect 93964 241708 93965 241772
rect 93899 241707 93965 241708
rect 89483 175948 89549 175949
rect 89483 175884 89484 175948
rect 89548 175884 89549 175948
rect 89483 175883 89549 175884
rect 88931 172548 88997 172549
rect 88931 172484 88932 172548
rect 88996 172484 88997 172548
rect 88931 172483 88997 172484
rect 84954 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 85574 158614
rect 84954 158294 85574 158378
rect 84954 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 85574 158294
rect 83411 149156 83477 149157
rect 83411 149092 83412 149156
rect 83476 149092 83477 149156
rect 83411 149091 83477 149092
rect 83411 141540 83477 141541
rect 83411 141476 83412 141540
rect 83476 141476 83477 141540
rect 83411 141475 83477 141476
rect 83414 136781 83474 141475
rect 84954 136782 85574 158058
rect 88934 136781 88994 172483
rect 83411 136780 83477 136781
rect 83411 136716 83412 136780
rect 83476 136716 83477 136780
rect 83411 136715 83477 136716
rect 88931 136780 88997 136781
rect 88931 136716 88932 136780
rect 88996 136716 88997 136780
rect 88931 136715 88997 136716
rect 90958 135557 91018 241707
rect 93902 240277 93962 241707
rect 93899 240276 93965 240277
rect 93899 240212 93900 240276
rect 93964 240212 93965 240276
rect 93899 240211 93965 240212
rect 97763 240140 97829 240141
rect 97763 240076 97764 240140
rect 97828 240076 97829 240140
rect 97763 240075 97829 240076
rect 91794 237454 92414 239592
rect 93715 237556 93781 237557
rect 93715 237492 93716 237556
rect 93780 237492 93781 237556
rect 93715 237491 93781 237492
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91507 144804 91573 144805
rect 91507 144740 91508 144804
rect 91572 144740 91573 144804
rect 91507 144739 91573 144740
rect 90955 135556 91021 135557
rect 90955 135492 90956 135556
rect 91020 135492 91021 135556
rect 90955 135491 91021 135492
rect 91510 132970 91570 144739
rect 91794 136782 92414 164898
rect 91510 132910 91754 132970
rect 77644 129454 77964 129486
rect 77644 129218 77686 129454
rect 77922 129218 77964 129454
rect 77644 129134 77964 129218
rect 77644 128898 77686 129134
rect 77922 128898 77964 129134
rect 77644 128866 77964 128898
rect 85575 129454 85895 129486
rect 85575 129218 85617 129454
rect 85853 129218 85895 129454
rect 85575 129134 85895 129218
rect 85575 128898 85617 129134
rect 85853 128898 85895 129134
rect 85575 128866 85895 128898
rect 91694 128370 91754 132910
rect 91694 128310 92306 128370
rect 73679 111454 73999 111486
rect 73679 111218 73721 111454
rect 73957 111218 73999 111454
rect 73679 111134 73999 111218
rect 73679 110898 73721 111134
rect 73957 110898 73999 111134
rect 73679 110866 73999 110898
rect 81609 111454 81929 111486
rect 81609 111218 81651 111454
rect 81887 111218 81929 111454
rect 81609 111134 81929 111218
rect 81609 110898 81651 111134
rect 81887 110898 81929 111134
rect 81609 110866 81929 110898
rect 89540 111454 89860 111486
rect 89540 111218 89582 111454
rect 89818 111218 89860 111454
rect 89540 111134 89860 111218
rect 89540 110898 89582 111134
rect 89818 110898 89860 111134
rect 89540 110866 89860 110898
rect 92246 92717 92306 128310
rect 93718 92717 93778 237491
rect 95514 205174 96134 239592
rect 97766 209790 97826 240075
rect 98134 238770 98194 254355
rect 100707 252516 100773 252517
rect 100707 252452 100708 252516
rect 100772 252452 100773 252516
rect 100707 252451 100773 252452
rect 95514 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 96134 205174
rect 97214 209730 97826 209790
rect 97950 238710 98194 238770
rect 97214 205053 97274 209730
rect 97211 205052 97277 205053
rect 97211 204988 97212 205052
rect 97276 204988 97277 205052
rect 97211 204987 97277 204988
rect 95514 204854 96134 204938
rect 95514 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 96134 204854
rect 95514 169174 96134 204618
rect 95514 168938 95546 169174
rect 95782 168938 95866 169174
rect 96102 168938 96134 169174
rect 95514 168854 96134 168938
rect 95514 168618 95546 168854
rect 95782 168618 95866 168854
rect 96102 168618 96134 168854
rect 94819 139636 94885 139637
rect 94819 139572 94820 139636
rect 94884 139572 94885 139636
rect 94819 139571 94885 139572
rect 94822 132157 94882 139571
rect 95514 136782 96134 168618
rect 96291 138140 96357 138141
rect 96291 138076 96292 138140
rect 96356 138076 96357 138140
rect 96291 138075 96357 138076
rect 95187 135420 95253 135421
rect 95187 135356 95188 135420
rect 95252 135356 95253 135420
rect 95187 135355 95253 135356
rect 94819 132156 94885 132157
rect 94819 132092 94820 132156
rect 94884 132092 94885 132156
rect 94819 132091 94885 132092
rect 94819 104140 94885 104141
rect 94819 104076 94820 104140
rect 94884 104076 94885 104140
rect 94819 104075 94885 104076
rect 92243 92716 92309 92717
rect 92243 92652 92244 92716
rect 92308 92652 92309 92716
rect 92243 92651 92309 92652
rect 93715 92716 93781 92717
rect 93715 92652 93716 92716
rect 93780 92652 93781 92716
rect 93715 92651 93781 92652
rect 94822 92173 94882 104075
rect 94819 92172 94885 92173
rect 94819 92108 94820 92172
rect 94884 92108 94885 92172
rect 94819 92107 94885 92108
rect 72739 91084 72805 91085
rect 72739 91020 72740 91084
rect 72804 91020 72805 91084
rect 72739 91019 72805 91020
rect 66483 87956 66549 87957
rect 66483 87892 66484 87956
rect 66548 87892 66549 87956
rect 66483 87891 66549 87892
rect 63234 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 63854 64894
rect 63234 64574 63854 64658
rect 63234 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 63854 64574
rect 63234 28894 63854 64338
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 68614 67574 90782
rect 66954 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 67574 68614
rect 66954 68294 67574 68378
rect 66954 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 67574 68294
rect 66954 32614 67574 68058
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 75454 74414 90782
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 79174 78134 90782
rect 77514 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 78134 79174
rect 77514 78854 78134 78938
rect 77514 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 78134 78854
rect 77514 43174 78134 78618
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 82894 81854 90782
rect 81234 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 81854 82894
rect 81234 82574 81854 82658
rect 81234 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 81854 82574
rect 81234 46894 81854 82338
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 86614 85574 90782
rect 84954 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 85574 86614
rect 84954 86294 85574 86378
rect 84954 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 85574 86294
rect 84954 50614 85574 86058
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 57454 92414 90782
rect 95190 85373 95250 135355
rect 96294 120053 96354 138075
rect 96291 120052 96357 120053
rect 96291 119988 96292 120052
rect 96356 119988 96357 120052
rect 96291 119987 96357 119988
rect 97214 92853 97274 204987
rect 97950 179485 98010 238710
rect 99234 208894 99854 239592
rect 99234 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 99854 208894
rect 99234 208574 99854 208658
rect 99234 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 99854 208574
rect 97947 179484 98013 179485
rect 97947 179420 97948 179484
rect 98012 179420 98013 179484
rect 97947 179419 98013 179420
rect 97950 108085 98010 179419
rect 99234 172894 99854 208338
rect 99234 172658 99266 172894
rect 99502 172658 99586 172894
rect 99822 172658 99854 172894
rect 99234 172574 99854 172658
rect 99234 172338 99266 172574
rect 99502 172338 99586 172574
rect 99822 172338 99854 172574
rect 99234 136894 99854 172338
rect 99234 136658 99266 136894
rect 99502 136658 99586 136894
rect 99822 136658 99854 136894
rect 99234 136574 99854 136658
rect 99234 136338 99266 136574
rect 99502 136338 99586 136574
rect 99822 136338 99854 136574
rect 98499 108356 98565 108357
rect 98499 108292 98500 108356
rect 98564 108292 98565 108356
rect 98499 108291 98565 108292
rect 97947 108084 98013 108085
rect 97947 108020 97948 108084
rect 98012 108020 98013 108084
rect 97947 108019 98013 108020
rect 97211 92852 97277 92853
rect 97211 92788 97212 92852
rect 97276 92788 97277 92852
rect 97211 92787 97277 92788
rect 95187 85372 95253 85373
rect 95187 85308 95188 85372
rect 95252 85308 95253 85372
rect 95187 85307 95253 85308
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 61174 96134 90782
rect 98502 89453 98562 108291
rect 99234 100894 99854 136338
rect 100710 105909 100770 252451
rect 100894 116653 100954 261427
rect 102954 248614 103574 284058
rect 102954 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 103574 248614
rect 102954 248294 103574 248378
rect 102954 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 103574 248294
rect 102954 212614 103574 248058
rect 102954 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 103574 212614
rect 102954 212294 103574 212378
rect 102954 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 103574 212294
rect 102954 176614 103574 212058
rect 102954 176378 102986 176614
rect 103222 176378 103306 176614
rect 103542 176378 103574 176614
rect 102954 176294 103574 176378
rect 102954 176058 102986 176294
rect 103222 176058 103306 176294
rect 103542 176058 103574 176294
rect 102954 140614 103574 176058
rect 102954 140378 102986 140614
rect 103222 140378 103306 140614
rect 103542 140378 103574 140614
rect 102954 140294 103574 140378
rect 102954 140058 102986 140294
rect 103222 140058 103306 140294
rect 103542 140058 103574 140294
rect 100891 116652 100957 116653
rect 100891 116588 100892 116652
rect 100956 116588 100957 116652
rect 100891 116587 100957 116588
rect 100707 105908 100773 105909
rect 100707 105844 100708 105908
rect 100772 105844 100773 105908
rect 100707 105843 100773 105844
rect 99234 100658 99266 100894
rect 99502 100658 99586 100894
rect 99822 100658 99854 100894
rect 99234 100574 99854 100658
rect 99234 100338 99266 100574
rect 99502 100338 99586 100574
rect 99822 100338 99854 100574
rect 98499 89452 98565 89453
rect 98499 89388 98500 89452
rect 98564 89388 98565 89452
rect 98499 89387 98565 89388
rect 95514 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 96134 61174
rect 95514 60854 96134 60938
rect 95514 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 96134 60854
rect 95514 25174 96134 60618
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 64894 99854 100338
rect 99234 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 99854 64894
rect 99234 64574 99854 64658
rect 99234 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 99854 64574
rect 99234 28894 99854 64338
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 104614 103574 140058
rect 102954 104378 102986 104614
rect 103222 104378 103306 104614
rect 103542 104378 103574 104614
rect 102954 104294 103574 104378
rect 102954 104058 102986 104294
rect 103222 104058 103306 104294
rect 103542 104058 103574 104294
rect 102954 68614 103574 104058
rect 102954 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 103574 68614
rect 102954 68294 103574 68378
rect 102954 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 103574 68294
rect 102954 32614 103574 68058
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 291454 110414 326898
rect 110646 323645 110706 433603
rect 110643 323644 110709 323645
rect 110643 323580 110644 323644
rect 110708 323580 110709 323644
rect 110643 323579 110709 323580
rect 111750 319429 111810 433603
rect 111934 390693 111994 472499
rect 113514 439174 114134 474618
rect 114323 460188 114389 460189
rect 114323 460124 114324 460188
rect 114388 460124 114389 460188
rect 114323 460123 114389 460124
rect 113514 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 114134 439174
rect 113514 438854 114134 438938
rect 113514 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 114134 438854
rect 112115 438156 112181 438157
rect 112115 438092 112116 438156
rect 112180 438092 112181 438156
rect 112115 438091 112181 438092
rect 112118 432853 112178 438091
rect 113219 436796 113285 436797
rect 113219 436732 113220 436796
rect 113284 436732 113285 436796
rect 113219 436731 113285 436732
rect 112115 432852 112181 432853
rect 112115 432788 112116 432852
rect 112180 432788 112181 432852
rect 112115 432787 112181 432788
rect 113222 396405 113282 436731
rect 113514 436356 114134 438618
rect 114326 418301 114386 460123
rect 114323 418300 114389 418301
rect 114323 418236 114324 418300
rect 114388 418236 114389 418300
rect 114323 418235 114389 418236
rect 114510 410549 114570 522275
rect 117234 514894 117854 550338
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 117234 478894 117854 514338
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 117234 442894 117854 478338
rect 117234 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 117854 442894
rect 117234 442574 117854 442658
rect 117234 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 117854 442574
rect 114691 417892 114757 417893
rect 114691 417828 114692 417892
rect 114756 417828 114757 417892
rect 114691 417827 114757 417828
rect 114507 410548 114573 410549
rect 114507 410484 114508 410548
rect 114572 410484 114573 410548
rect 114507 410483 114573 410484
rect 113219 396404 113285 396405
rect 113219 396340 113220 396404
rect 113284 396340 113285 396404
rect 113219 396339 113285 396340
rect 111931 390692 111997 390693
rect 111931 390628 111932 390692
rect 111996 390628 111997 390692
rect 111931 390627 111997 390628
rect 113514 367174 114134 388356
rect 114694 382941 114754 417827
rect 117234 406894 117854 442338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 120954 554614 121574 590058
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 518614 121574 554058
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 120954 482614 121574 518058
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120954 446614 121574 482058
rect 120954 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 121574 446614
rect 120954 446294 121574 446378
rect 120954 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 121574 446294
rect 118739 434892 118805 434893
rect 118739 434828 118740 434892
rect 118804 434828 118805 434892
rect 118739 434827 118805 434828
rect 117234 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 117854 406894
rect 117234 406574 117854 406658
rect 117234 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 117854 406574
rect 114691 382940 114757 382941
rect 114691 382876 114692 382940
rect 114756 382876 114757 382940
rect 114691 382875 114757 382876
rect 113514 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 114134 367174
rect 113514 366854 114134 366938
rect 113514 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 114134 366854
rect 113514 331174 114134 366618
rect 113514 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 114134 331174
rect 113514 330854 114134 330938
rect 113514 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 114134 330854
rect 111747 319428 111813 319429
rect 111747 319364 111748 319428
rect 111812 319364 111813 319428
rect 111747 319363 111813 319364
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 219454 110414 254898
rect 113514 295174 114134 330618
rect 113514 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 114134 295174
rect 113514 294854 114134 294938
rect 113514 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 114134 294854
rect 113514 259174 114134 294618
rect 113514 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 114134 259174
rect 113514 258854 114134 258938
rect 113514 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 114134 258854
rect 111563 237964 111629 237965
rect 111563 237900 111564 237964
rect 111628 237900 111629 237964
rect 111563 237899 111629 237900
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 111566 3501 111626 237899
rect 113514 223174 114134 258618
rect 113514 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 114134 223174
rect 113514 222854 114134 222938
rect 113514 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 114134 222854
rect 113514 187174 114134 222618
rect 113514 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 114134 187174
rect 113514 186854 114134 186938
rect 113514 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 114134 186854
rect 113514 151174 114134 186618
rect 113514 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 114134 151174
rect 113514 150854 114134 150938
rect 113514 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 114134 150854
rect 113514 115174 114134 150618
rect 113514 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 114134 115174
rect 113514 114854 114134 114938
rect 113514 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 114134 114854
rect 113514 79174 114134 114618
rect 113514 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 114134 79174
rect 113514 78854 114134 78938
rect 113514 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 114134 78854
rect 113514 43174 114134 78618
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 111563 3500 111629 3501
rect 111563 3436 111564 3500
rect 111628 3436 111629 3500
rect 111563 3435 111629 3436
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 370894 117854 406338
rect 117234 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 117854 370894
rect 117234 370574 117854 370658
rect 117234 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 117854 370574
rect 117234 334894 117854 370338
rect 117234 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 117854 334894
rect 117234 334574 117854 334658
rect 117234 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 117854 334574
rect 117234 298894 117854 334338
rect 118742 316709 118802 434827
rect 120954 410614 121574 446058
rect 120954 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 121574 410614
rect 120954 410294 121574 410378
rect 120954 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 121574 410294
rect 120954 374614 121574 410058
rect 120954 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 121574 374614
rect 120954 374294 121574 374378
rect 120954 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 121574 374294
rect 120954 338614 121574 374058
rect 120954 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 121574 338614
rect 120954 338294 121574 338378
rect 120954 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 121574 338294
rect 118739 316708 118805 316709
rect 118739 316644 118740 316708
rect 118804 316644 118805 316708
rect 118739 316643 118805 316644
rect 117234 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 117854 298894
rect 117234 298574 117854 298658
rect 117234 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 117854 298574
rect 117234 262894 117854 298338
rect 117234 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 117854 262894
rect 117234 262574 117854 262658
rect 117234 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 117854 262574
rect 117234 226894 117854 262338
rect 117234 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 117854 226894
rect 117234 226574 117854 226658
rect 117234 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 117854 226574
rect 117234 190894 117854 226338
rect 117234 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 117854 190894
rect 117234 190574 117854 190658
rect 117234 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 117854 190574
rect 117234 154894 117854 190338
rect 117234 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 117854 154894
rect 117234 154574 117854 154658
rect 117234 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 117854 154574
rect 117234 118894 117854 154338
rect 117234 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 117854 118894
rect 117234 118574 117854 118658
rect 117234 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 117854 118574
rect 117234 82894 117854 118338
rect 117234 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 117854 82894
rect 117234 82574 117854 82658
rect 117234 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 117854 82574
rect 117234 46894 117854 82338
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 302614 121574 338058
rect 120954 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 121574 302614
rect 120954 302294 121574 302378
rect 120954 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 121574 302294
rect 120954 266614 121574 302058
rect 120954 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 121574 266614
rect 120954 266294 121574 266378
rect 120954 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 121574 266294
rect 120954 230614 121574 266058
rect 120954 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 121574 230614
rect 120954 230294 121574 230378
rect 120954 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 121574 230294
rect 120954 194614 121574 230058
rect 120954 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 121574 194614
rect 120954 194294 121574 194378
rect 120954 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 121574 194294
rect 120954 158614 121574 194058
rect 120954 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 121574 158614
rect 120954 158294 121574 158378
rect 120954 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 121574 158294
rect 120954 122614 121574 158058
rect 120954 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 121574 122614
rect 120954 122294 121574 122378
rect 120954 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 121574 122294
rect 120954 86614 121574 122058
rect 120954 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 121574 86614
rect 120954 86294 121574 86378
rect 120954 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 121574 86294
rect 120954 50614 121574 86058
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 127794 165454 128414 200898
rect 127794 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 128414 165454
rect 127794 165134 128414 165218
rect 127794 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 128414 165134
rect 127794 129454 128414 164898
rect 127794 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 128414 129454
rect 127794 129134 128414 129218
rect 127794 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 128414 129134
rect 127794 93454 128414 128898
rect 127794 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 128414 93454
rect 127794 93134 128414 93218
rect 127794 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 128414 93134
rect 127794 57454 128414 92898
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 529174 132134 564618
rect 131514 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 132134 529174
rect 131514 528854 132134 528938
rect 131514 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 132134 528854
rect 131514 493174 132134 528618
rect 131514 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 132134 493174
rect 131514 492854 132134 492938
rect 131514 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 132134 492854
rect 131514 457174 132134 492618
rect 131514 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 132134 457174
rect 131514 456854 132134 456938
rect 131514 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 132134 456854
rect 131514 421174 132134 456618
rect 131514 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 132134 421174
rect 131514 420854 132134 420938
rect 131514 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 132134 420854
rect 131514 385174 132134 420618
rect 131514 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 132134 385174
rect 131514 384854 132134 384938
rect 131514 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 132134 384854
rect 131514 349174 132134 384618
rect 131514 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 132134 349174
rect 131514 348854 132134 348938
rect 131514 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 132134 348854
rect 131514 313174 132134 348618
rect 131514 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 132134 313174
rect 131514 312854 132134 312938
rect 131514 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 132134 312854
rect 131514 277174 132134 312618
rect 131514 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 132134 277174
rect 131514 276854 132134 276938
rect 131514 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 132134 276854
rect 131514 241174 132134 276618
rect 131514 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 132134 241174
rect 131514 240854 132134 240938
rect 131514 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 132134 240854
rect 131514 205174 132134 240618
rect 131514 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 132134 205174
rect 131514 204854 132134 204938
rect 131514 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 132134 204854
rect 131514 169174 132134 204618
rect 131514 168938 131546 169174
rect 131782 168938 131866 169174
rect 132102 168938 132134 169174
rect 131514 168854 132134 168938
rect 131514 168618 131546 168854
rect 131782 168618 131866 168854
rect 132102 168618 132134 168854
rect 131514 133174 132134 168618
rect 131514 132938 131546 133174
rect 131782 132938 131866 133174
rect 132102 132938 132134 133174
rect 131514 132854 132134 132938
rect 131514 132618 131546 132854
rect 131782 132618 131866 132854
rect 132102 132618 132134 132854
rect 131514 97174 132134 132618
rect 131514 96938 131546 97174
rect 131782 96938 131866 97174
rect 132102 96938 132134 97174
rect 131514 96854 132134 96938
rect 131514 96618 131546 96854
rect 131782 96618 131866 96854
rect 132102 96618 132134 96854
rect 131514 61174 132134 96618
rect 131514 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 132134 61174
rect 131514 60854 132134 60938
rect 131514 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 132134 60854
rect 131514 25174 132134 60618
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 532894 135854 568338
rect 135234 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 135854 532894
rect 135234 532574 135854 532658
rect 135234 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 135854 532574
rect 135234 496894 135854 532338
rect 135234 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 135854 496894
rect 135234 496574 135854 496658
rect 135234 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 135854 496574
rect 135234 460894 135854 496338
rect 135234 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 135854 460894
rect 135234 460574 135854 460658
rect 135234 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 135854 460574
rect 135234 424894 135854 460338
rect 135234 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 135854 424894
rect 135234 424574 135854 424658
rect 135234 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 135854 424574
rect 135234 388894 135854 424338
rect 135234 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 135854 388894
rect 135234 388574 135854 388658
rect 135234 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 135854 388574
rect 135234 352894 135854 388338
rect 135234 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 135854 352894
rect 135234 352574 135854 352658
rect 135234 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 135854 352574
rect 135234 316894 135854 352338
rect 135234 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 135854 316894
rect 135234 316574 135854 316658
rect 135234 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 135854 316574
rect 135234 280894 135854 316338
rect 135234 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 135854 280894
rect 135234 280574 135854 280658
rect 135234 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 135854 280574
rect 135234 244894 135854 280338
rect 135234 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 135854 244894
rect 135234 244574 135854 244658
rect 135234 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 135854 244574
rect 135234 208894 135854 244338
rect 135234 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 135854 208894
rect 135234 208574 135854 208658
rect 135234 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 135854 208574
rect 135234 172894 135854 208338
rect 135234 172658 135266 172894
rect 135502 172658 135586 172894
rect 135822 172658 135854 172894
rect 135234 172574 135854 172658
rect 135234 172338 135266 172574
rect 135502 172338 135586 172574
rect 135822 172338 135854 172574
rect 135234 136894 135854 172338
rect 135234 136658 135266 136894
rect 135502 136658 135586 136894
rect 135822 136658 135854 136894
rect 135234 136574 135854 136658
rect 135234 136338 135266 136574
rect 135502 136338 135586 136574
rect 135822 136338 135854 136574
rect 135234 100894 135854 136338
rect 135234 100658 135266 100894
rect 135502 100658 135586 100894
rect 135822 100658 135854 100894
rect 135234 100574 135854 100658
rect 135234 100338 135266 100574
rect 135502 100338 135586 100574
rect 135822 100338 135854 100574
rect 135234 64894 135854 100338
rect 135234 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 135854 64894
rect 135234 64574 135854 64658
rect 135234 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 135854 64574
rect 135234 28894 135854 64338
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 536614 139574 572058
rect 138954 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 139574 536614
rect 138954 536294 139574 536378
rect 138954 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 139574 536294
rect 138954 500614 139574 536058
rect 138954 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 139574 500614
rect 138954 500294 139574 500378
rect 138954 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 139574 500294
rect 138954 464614 139574 500058
rect 138954 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 139574 464614
rect 138954 464294 139574 464378
rect 138954 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 139574 464294
rect 138954 428614 139574 464058
rect 138954 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 139574 428614
rect 138954 428294 139574 428378
rect 138954 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 139574 428294
rect 138954 392614 139574 428058
rect 138954 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 139574 392614
rect 138954 392294 139574 392378
rect 138954 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 139574 392294
rect 138954 356614 139574 392058
rect 138954 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 139574 356614
rect 138954 356294 139574 356378
rect 138954 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 139574 356294
rect 138954 320614 139574 356058
rect 138954 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 139574 320614
rect 138954 320294 139574 320378
rect 138954 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 139574 320294
rect 138954 284614 139574 320058
rect 138954 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 139574 284614
rect 138954 284294 139574 284378
rect 138954 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 139574 284294
rect 138954 248614 139574 284058
rect 138954 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 139574 248614
rect 138954 248294 139574 248378
rect 138954 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 139574 248294
rect 138954 212614 139574 248058
rect 138954 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 139574 212614
rect 138954 212294 139574 212378
rect 138954 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 139574 212294
rect 138954 176614 139574 212058
rect 138954 176378 138986 176614
rect 139222 176378 139306 176614
rect 139542 176378 139574 176614
rect 138954 176294 139574 176378
rect 138954 176058 138986 176294
rect 139222 176058 139306 176294
rect 139542 176058 139574 176294
rect 138954 140614 139574 176058
rect 138954 140378 138986 140614
rect 139222 140378 139306 140614
rect 139542 140378 139574 140614
rect 138954 140294 139574 140378
rect 138954 140058 138986 140294
rect 139222 140058 139306 140294
rect 139542 140058 139574 140294
rect 138954 104614 139574 140058
rect 138954 104378 138986 104614
rect 139222 104378 139306 104614
rect 139542 104378 139574 104614
rect 138954 104294 139574 104378
rect 138954 104058 138986 104294
rect 139222 104058 139306 104294
rect 139542 104058 139574 104294
rect 138954 68614 139574 104058
rect 138954 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 139574 68614
rect 138954 68294 139574 68378
rect 138954 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 139574 68294
rect 138954 32614 139574 68058
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 147454 146414 182898
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 111454 146414 146898
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 145794 75454 146414 110898
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 149514 475174 150134 510618
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 439174 150134 474618
rect 149514 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 150134 439174
rect 149514 438854 150134 438938
rect 149514 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 150134 438854
rect 149514 403174 150134 438618
rect 149514 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 150134 403174
rect 149514 402854 150134 402938
rect 149514 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 150134 402854
rect 149514 367174 150134 402618
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 149514 331174 150134 366618
rect 149514 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 150134 331174
rect 149514 330854 150134 330938
rect 149514 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 150134 330854
rect 149514 295174 150134 330618
rect 149514 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 150134 295174
rect 149514 294854 150134 294938
rect 149514 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 150134 294854
rect 149514 259174 150134 294618
rect 149514 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 150134 259174
rect 149514 258854 150134 258938
rect 149514 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 150134 258854
rect 149514 223174 150134 258618
rect 149514 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 150134 223174
rect 149514 222854 150134 222938
rect 149514 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 150134 222854
rect 149514 187174 150134 222618
rect 149514 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 150134 187174
rect 149514 186854 150134 186938
rect 149514 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 150134 186854
rect 149514 151174 150134 186618
rect 149514 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 150134 151174
rect 149514 150854 150134 150938
rect 149514 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 150134 150854
rect 149514 115174 150134 150618
rect 149514 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 150134 115174
rect 149514 114854 150134 114938
rect 149514 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 150134 114854
rect 149514 79174 150134 114618
rect 149514 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 150134 79174
rect 149514 78854 150134 78938
rect 149514 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 150134 78854
rect 149514 43174 150134 78618
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 514894 153854 550338
rect 153234 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 153854 514894
rect 153234 514574 153854 514658
rect 153234 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 153854 514574
rect 153234 478894 153854 514338
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 442894 153854 478338
rect 153234 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 153854 442894
rect 153234 442574 153854 442658
rect 153234 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 153854 442574
rect 153234 406894 153854 442338
rect 153234 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 153854 406894
rect 153234 406574 153854 406658
rect 153234 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 153854 406574
rect 153234 370894 153854 406338
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 153234 334894 153854 370338
rect 153234 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 153854 334894
rect 153234 334574 153854 334658
rect 153234 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 153854 334574
rect 153234 298894 153854 334338
rect 153234 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 153854 298894
rect 153234 298574 153854 298658
rect 153234 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 153854 298574
rect 153234 262894 153854 298338
rect 153234 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 153854 262894
rect 153234 262574 153854 262658
rect 153234 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 153854 262574
rect 153234 226894 153854 262338
rect 153234 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 153854 226894
rect 153234 226574 153854 226658
rect 153234 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 153854 226574
rect 153234 190894 153854 226338
rect 153234 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 153854 190894
rect 153234 190574 153854 190658
rect 153234 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 153854 190574
rect 153234 154894 153854 190338
rect 153234 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 153854 154894
rect 153234 154574 153854 154658
rect 153234 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 153854 154574
rect 153234 118894 153854 154338
rect 153234 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 153854 118894
rect 153234 118574 153854 118658
rect 153234 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 153854 118574
rect 153234 82894 153854 118338
rect 153234 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 153854 82894
rect 153234 82574 153854 82658
rect 153234 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 153854 82574
rect 153234 46894 153854 82338
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 518614 157574 554058
rect 156954 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 157574 518614
rect 156954 518294 157574 518378
rect 156954 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 157574 518294
rect 156954 482614 157574 518058
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156954 446614 157574 482058
rect 156954 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 157574 446614
rect 156954 446294 157574 446378
rect 156954 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 157574 446294
rect 156954 410614 157574 446058
rect 156954 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 157574 410614
rect 156954 410294 157574 410378
rect 156954 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 157574 410294
rect 156954 374614 157574 410058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 160691 396676 160757 396677
rect 160691 396612 160692 396676
rect 160756 396612 160757 396676
rect 160691 396611 160757 396612
rect 156954 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 157574 374614
rect 156954 374294 157574 374378
rect 156954 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 157574 374294
rect 156954 338614 157574 374058
rect 160694 372605 160754 396611
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 160691 372604 160757 372605
rect 160691 372540 160692 372604
rect 160756 372540 160757 372604
rect 160691 372539 160757 372540
rect 156954 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 157574 338614
rect 156954 338294 157574 338378
rect 156954 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 157574 338294
rect 156954 302614 157574 338058
rect 156954 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 157574 302614
rect 156954 302294 157574 302378
rect 156954 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 157574 302294
rect 156954 266614 157574 302058
rect 156954 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 157574 266614
rect 156954 266294 157574 266378
rect 156954 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 157574 266294
rect 156954 230614 157574 266058
rect 160694 246261 160754 372539
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 160691 246260 160757 246261
rect 160691 246196 160692 246260
rect 160756 246196 160757 246260
rect 160691 246195 160757 246196
rect 156954 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 157574 230614
rect 156954 230294 157574 230378
rect 156954 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 157574 230294
rect 156954 194614 157574 230058
rect 156954 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 157574 194614
rect 156954 194294 157574 194378
rect 156954 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 157574 194294
rect 156954 158614 157574 194058
rect 156954 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 157574 158614
rect 156954 158294 157574 158378
rect 156954 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 157574 158294
rect 156954 122614 157574 158058
rect 156954 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 157574 122614
rect 156954 122294 157574 122378
rect 156954 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 157574 122294
rect 156954 86614 157574 122058
rect 156954 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 157574 86614
rect 156954 86294 157574 86378
rect 156954 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 157574 86294
rect 156954 50614 157574 86058
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 163794 165454 164414 200898
rect 163794 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 164414 165454
rect 163794 165134 164414 165218
rect 163794 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 164414 165134
rect 163794 129454 164414 164898
rect 163794 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 164414 129454
rect 163794 129134 164414 129218
rect 163794 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 164414 129134
rect 163794 93454 164414 128898
rect 163794 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 164414 93454
rect 163794 93134 164414 93218
rect 163794 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 164414 93134
rect 163794 57454 164414 92898
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 565174 168134 600618
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 529174 168134 564618
rect 167514 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 168134 529174
rect 167514 528854 168134 528938
rect 167514 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 168134 528854
rect 167514 493174 168134 528618
rect 167514 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 168134 493174
rect 167514 492854 168134 492938
rect 167514 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 168134 492854
rect 167514 457174 168134 492618
rect 167514 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 168134 457174
rect 167514 456854 168134 456938
rect 167514 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 168134 456854
rect 167514 421174 168134 456618
rect 167514 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 168134 421174
rect 167514 420854 168134 420938
rect 167514 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 168134 420854
rect 167514 385174 168134 420618
rect 167514 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 168134 385174
rect 167514 384854 168134 384938
rect 167514 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 168134 384854
rect 167514 349174 168134 384618
rect 167514 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 168134 349174
rect 167514 348854 168134 348938
rect 167514 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 168134 348854
rect 167514 313174 168134 348618
rect 167514 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 168134 313174
rect 167514 312854 168134 312938
rect 167514 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 168134 312854
rect 167514 277174 168134 312618
rect 167514 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 168134 277174
rect 167514 276854 168134 276938
rect 167514 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 168134 276854
rect 167514 241174 168134 276618
rect 167514 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 168134 241174
rect 167514 240854 168134 240938
rect 167514 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 168134 240854
rect 167514 205174 168134 240618
rect 167514 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 168134 205174
rect 167514 204854 168134 204938
rect 167514 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 168134 204854
rect 167514 169174 168134 204618
rect 167514 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 168134 169174
rect 167514 168854 168134 168938
rect 167514 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 168134 168854
rect 167514 133174 168134 168618
rect 167514 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 168134 133174
rect 167514 132854 168134 132938
rect 167514 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 168134 132854
rect 167514 97174 168134 132618
rect 167514 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 168134 97174
rect 167514 96854 168134 96938
rect 167514 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 168134 96854
rect 167514 61174 168134 96618
rect 167514 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 168134 61174
rect 167514 60854 168134 60938
rect 167514 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 168134 60854
rect 167514 25174 168134 60618
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 171234 568894 171854 604338
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 171234 532894 171854 568338
rect 171234 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 171854 532894
rect 171234 532574 171854 532658
rect 171234 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 171854 532574
rect 171234 496894 171854 532338
rect 171234 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 171854 496894
rect 171234 496574 171854 496658
rect 171234 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 171854 496574
rect 171234 460894 171854 496338
rect 171234 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 171854 460894
rect 171234 460574 171854 460658
rect 171234 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 171854 460574
rect 171234 424894 171854 460338
rect 171234 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 171854 424894
rect 171234 424574 171854 424658
rect 171234 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 171854 424574
rect 171234 388894 171854 424338
rect 171234 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 171854 388894
rect 171234 388574 171854 388658
rect 171234 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 171854 388574
rect 171234 352894 171854 388338
rect 171234 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 171854 352894
rect 171234 352574 171854 352658
rect 171234 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 171854 352574
rect 171234 316894 171854 352338
rect 171234 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 171854 316894
rect 171234 316574 171854 316658
rect 171234 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 171854 316574
rect 171234 280894 171854 316338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 572614 175574 608058
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 536614 175574 572058
rect 174954 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 175574 536614
rect 174954 536294 175574 536378
rect 174954 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 175574 536294
rect 174954 500614 175574 536058
rect 174954 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 175574 500614
rect 174954 500294 175574 500378
rect 174954 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 175574 500294
rect 174954 464614 175574 500058
rect 174954 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 175574 464614
rect 174954 464294 175574 464378
rect 174954 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 175574 464294
rect 174954 428614 175574 464058
rect 174954 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 175574 428614
rect 174954 428294 175574 428378
rect 174954 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 175574 428294
rect 174954 392614 175574 428058
rect 174954 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 175574 392614
rect 174954 392294 175574 392378
rect 174954 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 175574 392294
rect 174954 356614 175574 392058
rect 174954 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 175574 356614
rect 174954 356294 175574 356378
rect 174954 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 175574 356294
rect 174954 320614 175574 356058
rect 174954 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 175574 320614
rect 174954 320294 175574 320378
rect 174954 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 175574 320294
rect 173019 298892 173085 298893
rect 173019 298828 173020 298892
rect 173084 298828 173085 298892
rect 173019 298827 173085 298828
rect 171234 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 171854 280894
rect 171234 280574 171854 280658
rect 171234 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 171854 280574
rect 171234 244894 171854 280338
rect 173022 261493 173082 298827
rect 174954 284614 175574 320058
rect 174954 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 175574 284614
rect 174954 284294 175574 284378
rect 174954 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 175574 284294
rect 173019 261492 173085 261493
rect 173019 261428 173020 261492
rect 173084 261428 173085 261492
rect 173019 261427 173085 261428
rect 171234 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 171854 244894
rect 171234 244574 171854 244658
rect 171234 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 171854 244574
rect 171234 208894 171854 244338
rect 171234 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 171854 208894
rect 171234 208574 171854 208658
rect 171234 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 171854 208574
rect 171234 172894 171854 208338
rect 171234 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 171854 172894
rect 171234 172574 171854 172658
rect 171234 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 171854 172574
rect 171234 136894 171854 172338
rect 171234 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 171854 136894
rect 171234 136574 171854 136658
rect 171234 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 171854 136574
rect 171234 100894 171854 136338
rect 171234 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 171854 100894
rect 171234 100574 171854 100658
rect 171234 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 171854 100574
rect 171234 64894 171854 100338
rect 171234 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 171854 64894
rect 171234 64574 171854 64658
rect 171234 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 171854 64574
rect 171234 28894 171854 64338
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 248614 175574 284058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 547174 186134 582618
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 475174 186134 510618
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 439174 186134 474618
rect 185514 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 186134 439174
rect 185514 438854 186134 438938
rect 185514 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 186134 438854
rect 185514 403174 186134 438618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 550894 189854 586338
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 514894 189854 550338
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 189234 478894 189854 514338
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 189234 442894 189854 478338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 554614 193574 590058
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 518614 193574 554058
rect 192954 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 193574 518614
rect 192954 518294 193574 518378
rect 192954 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 193574 518294
rect 192954 482614 193574 518058
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 192954 452356 193574 482058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 197123 458284 197189 458285
rect 197123 458220 197124 458284
rect 197188 458220 197189 458284
rect 197123 458219 197189 458220
rect 194547 453116 194613 453117
rect 194547 453052 194548 453116
rect 194612 453052 194613 453116
rect 194547 453051 194613 453052
rect 193811 450396 193877 450397
rect 193811 450332 193812 450396
rect 193876 450332 193877 450396
rect 193811 450331 193877 450332
rect 193443 449716 193509 449717
rect 193443 449652 193444 449716
rect 193508 449652 193509 449716
rect 193443 449651 193509 449652
rect 193446 442917 193506 449651
rect 189234 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 189854 442894
rect 193443 442916 193509 442917
rect 193443 442852 193444 442916
rect 193508 442852 193509 442916
rect 193443 442851 193509 442852
rect 189234 442574 189854 442658
rect 189234 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 189854 442574
rect 188843 421020 188909 421021
rect 188843 420956 188844 421020
rect 188908 420956 188909 421020
rect 188843 420955 188909 420956
rect 188291 414084 188357 414085
rect 188291 414020 188292 414084
rect 188356 414020 188357 414084
rect 188291 414019 188357 414020
rect 185514 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 186134 403174
rect 185514 402854 186134 402938
rect 185514 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 186134 402854
rect 185514 367174 186134 402618
rect 188294 387565 188354 414019
rect 188291 387564 188357 387565
rect 188291 387500 188292 387564
rect 188356 387500 188357 387564
rect 188291 387499 188357 387500
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 185514 331174 186134 366618
rect 188846 355469 188906 420955
rect 189234 406894 189854 442338
rect 193814 441630 193874 450331
rect 194550 450261 194610 453051
rect 194547 450260 194613 450261
rect 194547 450196 194548 450260
rect 194612 450196 194613 450260
rect 194547 450195 194613 450196
rect 193446 441570 193874 441630
rect 192707 440740 192773 440741
rect 192707 440676 192708 440740
rect 192772 440676 192773 440740
rect 192707 440675 192773 440676
rect 189234 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 189854 406894
rect 189234 406574 189854 406658
rect 189234 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 189854 406574
rect 189234 370894 189854 406338
rect 192710 380221 192770 440675
rect 193446 432581 193506 441570
rect 193443 432580 193509 432581
rect 193443 432516 193444 432580
rect 193508 432516 193509 432580
rect 193443 432515 193509 432516
rect 193259 430948 193325 430949
rect 193259 430884 193260 430948
rect 193324 430884 193325 430948
rect 193259 430883 193325 430884
rect 193262 391237 193322 430883
rect 193811 392596 193877 392597
rect 193811 392532 193812 392596
rect 193876 392532 193877 392596
rect 193811 392531 193877 392532
rect 193259 391236 193325 391237
rect 193259 391172 193260 391236
rect 193324 391172 193325 391236
rect 193259 391171 193325 391172
rect 192707 380220 192773 380221
rect 192707 380156 192708 380220
rect 192772 380156 192773 380220
rect 192707 380155 192773 380156
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 188843 355468 188909 355469
rect 188843 355404 188844 355468
rect 188908 355404 188909 355468
rect 188843 355403 188909 355404
rect 185514 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 186134 331174
rect 185514 330854 186134 330938
rect 185514 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 186134 330854
rect 184059 305284 184125 305285
rect 184059 305220 184060 305284
rect 184124 305220 184125 305284
rect 184059 305219 184125 305220
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 184062 267205 184122 305219
rect 185514 295174 186134 330618
rect 189234 334894 189854 370338
rect 189234 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 189854 334894
rect 189234 334574 189854 334658
rect 189234 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 189854 334574
rect 186819 303788 186885 303789
rect 186819 303724 186820 303788
rect 186884 303724 186885 303788
rect 186819 303723 186885 303724
rect 185514 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 186134 295174
rect 185514 294854 186134 294938
rect 185514 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 186134 294854
rect 184059 267204 184125 267205
rect 184059 267140 184060 267204
rect 184124 267140 184125 267204
rect 184059 267139 184125 267140
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 177251 251292 177317 251293
rect 177251 251228 177252 251292
rect 177316 251228 177317 251292
rect 177251 251227 177317 251228
rect 174954 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 175574 248614
rect 174954 248294 175574 248378
rect 174954 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 175574 248294
rect 174954 212614 175574 248058
rect 174954 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 175574 212614
rect 174954 212294 175574 212378
rect 174954 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 175574 212294
rect 174954 176614 175574 212058
rect 174954 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 175574 176614
rect 174954 176294 175574 176378
rect 174954 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 175574 176294
rect 174954 140614 175574 176058
rect 177254 151061 177314 251227
rect 181794 219454 182414 254898
rect 185514 259174 186134 294618
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 184243 245716 184309 245717
rect 184243 245652 184244 245716
rect 184308 245652 184309 245716
rect 184243 245651 184309 245652
rect 184059 227764 184125 227765
rect 184059 227700 184060 227764
rect 184124 227700 184125 227764
rect 184059 227699 184125 227700
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 177251 151060 177317 151061
rect 177251 150996 177252 151060
rect 177316 150996 177317 151060
rect 177251 150995 177317 150996
rect 174954 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 175574 140614
rect 174954 140294 175574 140378
rect 174954 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 175574 140294
rect 174954 104614 175574 140058
rect 174954 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 175574 104614
rect 174954 104294 175574 104378
rect 174954 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 175574 104294
rect 174954 68614 175574 104058
rect 174954 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 175574 68614
rect 174954 68294 175574 68378
rect 174954 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 175574 68294
rect 174954 32614 175574 68058
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 184062 108085 184122 227699
rect 184246 152421 184306 245651
rect 185514 223174 186134 258618
rect 185514 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 186134 223174
rect 185514 222854 186134 222938
rect 185514 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 186134 222854
rect 185514 187174 186134 222618
rect 186822 220149 186882 303723
rect 189234 298894 189854 334338
rect 192954 374614 193574 388356
rect 192954 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 193574 374614
rect 192954 374294 193574 374378
rect 192954 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 193574 374294
rect 192954 338614 193574 374058
rect 193814 358053 193874 392531
rect 193811 358052 193877 358053
rect 193811 357988 193812 358052
rect 193876 357988 193877 358052
rect 193811 357987 193877 357988
rect 193814 338741 193874 357987
rect 193811 338740 193877 338741
rect 193811 338676 193812 338740
rect 193876 338676 193877 338740
rect 193811 338675 193877 338676
rect 192954 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 193574 338614
rect 192954 338294 193574 338378
rect 192954 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 193574 338294
rect 191603 316708 191669 316709
rect 191603 316644 191604 316708
rect 191668 316644 191669 316708
rect 191603 316643 191669 316644
rect 191606 301613 191666 316643
rect 192954 303592 193574 338058
rect 194550 302293 194610 450195
rect 197126 376005 197186 458219
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 452356 200414 452898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 203514 565174 204134 600618
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 203514 529174 204134 564618
rect 203514 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 204134 529174
rect 203514 528854 204134 528938
rect 203514 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 204134 528854
rect 203514 493174 204134 528618
rect 203514 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 204134 493174
rect 203514 492854 204134 492938
rect 203514 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 204134 492854
rect 203514 457174 204134 492618
rect 203514 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 204134 457174
rect 203514 456854 204134 456938
rect 203514 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 204134 456854
rect 203514 452356 204134 456618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 532894 207854 568338
rect 207234 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 207854 532894
rect 207234 532574 207854 532658
rect 207234 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 207854 532574
rect 207234 496894 207854 532338
rect 207234 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 207854 496894
rect 207234 496574 207854 496658
rect 207234 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 207854 496574
rect 207234 460894 207854 496338
rect 207234 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 207854 460894
rect 207234 460574 207854 460658
rect 207234 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 207854 460574
rect 207234 452356 207854 460338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 536614 211574 572058
rect 210954 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 211574 536614
rect 210954 536294 211574 536378
rect 210954 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 211574 536294
rect 210954 500614 211574 536058
rect 210954 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 211574 500614
rect 210954 500294 211574 500378
rect 210954 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 211574 500294
rect 210954 464614 211574 500058
rect 210954 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 211574 464614
rect 210954 464294 211574 464378
rect 210954 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 211574 464294
rect 210954 452356 211574 464058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 452356 218414 470898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 547174 222134 582618
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 511174 222134 546618
rect 221514 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 222134 511174
rect 221514 510854 222134 510938
rect 221514 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 222134 510854
rect 221514 475174 222134 510618
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 221514 452356 222134 474618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 550894 225854 586338
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 514894 225854 550338
rect 225234 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 225854 514894
rect 225234 514574 225854 514658
rect 225234 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 225854 514574
rect 225234 478894 225854 514338
rect 225234 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 225854 478894
rect 225234 478574 225854 478658
rect 225234 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 225854 478574
rect 225234 452356 225854 478338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 554614 229574 590058
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 518614 229574 554058
rect 228954 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 229574 518614
rect 228954 518294 229574 518378
rect 228954 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 229574 518294
rect 228954 482614 229574 518058
rect 228954 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 229574 482614
rect 228954 482294 229574 482378
rect 228954 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 229574 482294
rect 228954 452356 229574 482058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 452356 236414 452898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 601174 240134 636618
rect 239514 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 240134 601174
rect 239514 600854 240134 600938
rect 239514 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 240134 600854
rect 239514 565174 240134 600618
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 239514 529174 240134 564618
rect 239514 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 240134 529174
rect 239514 528854 240134 528938
rect 239514 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 240134 528854
rect 239514 493174 240134 528618
rect 239514 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 240134 493174
rect 239514 492854 240134 492938
rect 239514 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 240134 492854
rect 239514 457174 240134 492618
rect 239514 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 240134 457174
rect 239514 456854 240134 456938
rect 239514 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 240134 456854
rect 239514 452356 240134 456618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 604894 243854 640338
rect 243234 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 243854 604894
rect 243234 604574 243854 604658
rect 243234 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 243854 604574
rect 243234 568894 243854 604338
rect 243234 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 243854 568894
rect 243234 568574 243854 568658
rect 243234 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 243854 568574
rect 243234 532894 243854 568338
rect 243234 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 243854 532894
rect 243234 532574 243854 532658
rect 243234 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 243854 532574
rect 243234 496894 243854 532338
rect 243234 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 243854 496894
rect 243234 496574 243854 496658
rect 243234 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 243854 496574
rect 243234 460894 243854 496338
rect 243234 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 243854 460894
rect 243234 460574 243854 460658
rect 243234 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 243854 460574
rect 241651 452980 241717 452981
rect 241651 452916 241652 452980
rect 241716 452916 241717 452980
rect 241651 452915 241717 452916
rect 197776 435454 198096 435486
rect 197776 435218 197818 435454
rect 198054 435218 198096 435454
rect 197776 435134 198096 435218
rect 197776 434898 197818 435134
rect 198054 434898 198096 435134
rect 197776 434866 198096 434898
rect 228496 435454 228816 435486
rect 228496 435218 228538 435454
rect 228774 435218 228816 435454
rect 228496 435134 228816 435218
rect 228496 434898 228538 435134
rect 228774 434898 228816 435134
rect 228496 434866 228816 434898
rect 213136 417454 213456 417486
rect 213136 417218 213178 417454
rect 213414 417218 213456 417454
rect 213136 417134 213456 417218
rect 213136 416898 213178 417134
rect 213414 416898 213456 417134
rect 213136 416866 213456 416898
rect 197776 399454 198096 399486
rect 197776 399218 197818 399454
rect 198054 399218 198096 399454
rect 197776 399134 198096 399218
rect 197776 398898 197818 399134
rect 198054 398898 198096 399134
rect 197776 398866 198096 398898
rect 228496 399454 228816 399486
rect 228496 399218 228538 399454
rect 228774 399218 228816 399454
rect 228496 399134 228816 399218
rect 228496 398898 228538 399134
rect 228774 398898 228816 399134
rect 228496 398866 228816 398898
rect 199794 381454 200414 388356
rect 201539 387020 201605 387021
rect 201539 386956 201540 387020
rect 201604 386956 201605 387020
rect 201539 386955 201605 386956
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 197123 376004 197189 376005
rect 197123 375940 197124 376004
rect 197188 375940 197189 376004
rect 197123 375939 197189 375940
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199331 323100 199397 323101
rect 199331 323036 199332 323100
rect 199396 323036 199397 323100
rect 199331 323035 199397 323036
rect 192707 302292 192773 302293
rect 192707 302228 192708 302292
rect 192772 302228 192773 302292
rect 192707 302227 192773 302228
rect 194547 302292 194613 302293
rect 194547 302228 194548 302292
rect 194612 302228 194613 302292
rect 194547 302227 194613 302228
rect 191603 301612 191669 301613
rect 191603 301548 191604 301612
rect 191668 301548 191669 301612
rect 191603 301547 191669 301548
rect 191971 299572 192037 299573
rect 191971 299508 191972 299572
rect 192036 299508 192037 299572
rect 191971 299507 192037 299508
rect 189234 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 189854 298894
rect 189234 298574 189854 298658
rect 189234 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 189854 298574
rect 188291 298212 188357 298213
rect 188291 298148 188292 298212
rect 188356 298148 188357 298212
rect 188291 298147 188357 298148
rect 188294 268565 188354 298147
rect 188843 273324 188909 273325
rect 188843 273260 188844 273324
rect 188908 273260 188909 273324
rect 188843 273259 188909 273260
rect 188291 268564 188357 268565
rect 188291 268500 188292 268564
rect 188356 268500 188357 268564
rect 188291 268499 188357 268500
rect 188291 241636 188357 241637
rect 188291 241572 188292 241636
rect 188356 241572 188357 241636
rect 188291 241571 188357 241572
rect 186819 220148 186885 220149
rect 186819 220084 186820 220148
rect 186884 220084 186885 220148
rect 186819 220083 186885 220084
rect 185514 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 186134 187174
rect 185514 186854 186134 186938
rect 185514 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 186134 186854
rect 184243 152420 184309 152421
rect 184243 152356 184244 152420
rect 184308 152356 184309 152420
rect 184243 152355 184309 152356
rect 185514 151174 186134 186618
rect 187555 182884 187621 182885
rect 187555 182820 187556 182884
rect 187620 182820 187621 182884
rect 187555 182819 187621 182820
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 185514 115174 186134 150618
rect 185514 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 186134 115174
rect 185514 114854 186134 114938
rect 185514 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 186134 114854
rect 184059 108084 184125 108085
rect 184059 108020 184060 108084
rect 184124 108020 184125 108084
rect 184059 108019 184125 108020
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 79174 186134 114618
rect 187558 107541 187618 182819
rect 188294 146981 188354 241571
rect 188846 240141 188906 273259
rect 189234 262894 189854 298338
rect 191419 298076 191485 298077
rect 191419 298012 191420 298076
rect 191484 298012 191485 298076
rect 191419 298011 191485 298012
rect 190315 274684 190381 274685
rect 190315 274620 190316 274684
rect 190380 274620 190381 274684
rect 190315 274619 190381 274620
rect 189234 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 189854 262894
rect 189234 262574 189854 262658
rect 189234 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 189854 262574
rect 188843 240140 188909 240141
rect 188843 240076 188844 240140
rect 188908 240076 188909 240140
rect 188843 240075 188909 240076
rect 189234 226894 189854 262338
rect 189234 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 189854 226894
rect 189234 226574 189854 226658
rect 189234 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 189854 226574
rect 188843 201380 188909 201381
rect 188843 201316 188844 201380
rect 188908 201316 188909 201380
rect 188843 201315 188909 201316
rect 188291 146980 188357 146981
rect 188291 146916 188292 146980
rect 188356 146916 188357 146980
rect 188291 146915 188357 146916
rect 188846 135149 188906 201315
rect 189234 190894 189854 226338
rect 190318 215933 190378 274619
rect 190315 215932 190381 215933
rect 190315 215868 190316 215932
rect 190380 215868 190381 215932
rect 190315 215867 190381 215868
rect 189234 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 189854 190894
rect 189234 190574 189854 190658
rect 189234 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 189854 190574
rect 189234 154894 189854 190338
rect 190315 161668 190381 161669
rect 190315 161604 190316 161668
rect 190380 161604 190381 161668
rect 190315 161603 190381 161604
rect 189234 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 189854 154894
rect 189234 154574 189854 154658
rect 189234 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 189854 154574
rect 188843 135148 188909 135149
rect 188843 135084 188844 135148
rect 188908 135084 188909 135148
rect 188843 135083 188909 135084
rect 189234 118894 189854 154338
rect 190318 131205 190378 161603
rect 190315 131204 190381 131205
rect 190315 131140 190316 131204
rect 190380 131140 190381 131204
rect 190315 131139 190381 131140
rect 191422 129301 191482 298011
rect 191974 293181 192034 299507
rect 192710 297397 192770 302227
rect 193259 301612 193325 301613
rect 193259 301548 193260 301612
rect 193324 301548 193325 301612
rect 193259 301547 193325 301548
rect 193262 300117 193322 301547
rect 193259 300116 193325 300117
rect 193259 300052 193260 300116
rect 193324 300052 193325 300116
rect 193259 300051 193325 300052
rect 192707 297396 192773 297397
rect 192707 297332 192708 297396
rect 192772 297332 192773 297396
rect 192707 297331 192773 297332
rect 191971 293180 192037 293181
rect 191971 293116 191972 293180
rect 192036 293116 192037 293180
rect 191971 293115 192037 293116
rect 192707 293180 192773 293181
rect 192707 293116 192708 293180
rect 192772 293116 192773 293180
rect 192707 293115 192773 293116
rect 192710 292637 192770 293115
rect 192707 292636 192773 292637
rect 192707 292572 192708 292636
rect 192772 292572 192773 292636
rect 192707 292571 192773 292572
rect 191603 291276 191669 291277
rect 191603 291212 191604 291276
rect 191668 291212 191669 291276
rect 191603 291211 191669 291212
rect 191419 129300 191485 129301
rect 191419 129236 191420 129300
rect 191484 129236 191485 129300
rect 191419 129235 191485 129236
rect 189234 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 189854 118894
rect 189234 118574 189854 118658
rect 189234 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 189854 118574
rect 187555 107540 187621 107541
rect 187555 107476 187556 107540
rect 187620 107476 187621 107540
rect 187555 107475 187621 107476
rect 187558 107130 187618 107475
rect 187558 107070 187802 107130
rect 187742 85509 187802 107070
rect 187739 85508 187805 85509
rect 187739 85444 187740 85508
rect 187804 85444 187805 85508
rect 187739 85443 187805 85444
rect 185514 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 186134 79174
rect 185514 78854 186134 78938
rect 185514 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 186134 78854
rect 185514 43174 186134 78618
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 82894 189854 118338
rect 191606 118013 191666 291211
rect 192710 217293 192770 292571
rect 197776 291454 198096 291486
rect 197776 291218 197818 291454
rect 198054 291218 198096 291454
rect 197776 291134 198096 291218
rect 197776 290898 197818 291134
rect 198054 290898 198096 291134
rect 197776 290866 198096 290898
rect 193443 265572 193509 265573
rect 193443 265508 193444 265572
rect 193508 265508 193509 265572
rect 193443 265507 193509 265508
rect 193446 258090 193506 265507
rect 193446 258030 193874 258090
rect 193259 251836 193325 251837
rect 193259 251772 193260 251836
rect 193324 251772 193325 251836
rect 193259 251771 193325 251772
rect 193262 242861 193322 251771
rect 193259 242860 193325 242861
rect 193259 242796 193260 242860
rect 193324 242796 193325 242860
rect 193259 242795 193325 242796
rect 192954 230614 193574 239592
rect 192954 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 193574 230614
rect 192954 230294 193574 230378
rect 192954 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 193574 230294
rect 192707 217292 192773 217293
rect 192707 217228 192708 217292
rect 192772 217228 192773 217292
rect 192707 217227 192773 217228
rect 192954 194614 193574 230058
rect 192954 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 193574 194614
rect 192954 194294 193574 194378
rect 192954 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 193574 194294
rect 192954 158614 193574 194058
rect 192954 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 193574 158614
rect 192954 158294 193574 158378
rect 192954 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 193574 158294
rect 192954 143035 193574 158058
rect 193814 153101 193874 258030
rect 197776 255454 198096 255486
rect 197776 255218 197818 255454
rect 198054 255218 198096 255454
rect 197776 255134 198096 255218
rect 197776 254898 197818 255134
rect 198054 254898 198096 255134
rect 197776 254866 198096 254898
rect 199334 161669 199394 323035
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 303592 200414 308898
rect 200619 303516 200685 303517
rect 200619 303452 200620 303516
rect 200684 303452 200685 303516
rect 200619 303451 200685 303452
rect 199794 237454 200414 239592
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 200622 235789 200682 303451
rect 201542 241501 201602 386955
rect 203514 385174 204134 388356
rect 203514 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 204134 385174
rect 203514 384854 204134 384938
rect 203514 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 204134 384854
rect 203011 376004 203077 376005
rect 203011 375940 203012 376004
rect 203076 375940 203077 376004
rect 203011 375939 203077 375940
rect 201539 241500 201605 241501
rect 201539 241436 201540 241500
rect 201604 241436 201605 241500
rect 201539 241435 201605 241436
rect 203014 240141 203074 375939
rect 203514 349174 204134 384618
rect 203514 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 204134 349174
rect 203514 348854 204134 348938
rect 203514 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 204134 348854
rect 203514 313174 204134 348618
rect 203514 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 204134 313174
rect 203514 312854 204134 312938
rect 203514 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 204134 312854
rect 203514 303592 204134 312618
rect 207234 352894 207854 388356
rect 208347 385660 208413 385661
rect 208347 385596 208348 385660
rect 208412 385596 208413 385660
rect 208347 385595 208413 385596
rect 207234 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 207854 352894
rect 207234 352574 207854 352658
rect 207234 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 207854 352574
rect 207234 316894 207854 352338
rect 207234 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 207854 316894
rect 207234 316574 207854 316658
rect 207234 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 207854 316574
rect 206139 307732 206205 307733
rect 206139 307668 206140 307732
rect 206204 307668 206205 307732
rect 206139 307667 206205 307668
rect 204299 301476 204365 301477
rect 204299 301412 204300 301476
rect 204364 301412 204365 301476
rect 204299 301411 204365 301412
rect 203011 240140 203077 240141
rect 203011 240076 203012 240140
rect 203076 240076 203077 240140
rect 203011 240075 203077 240076
rect 201539 237964 201605 237965
rect 201539 237900 201540 237964
rect 201604 237900 201605 237964
rect 201539 237899 201605 237900
rect 200619 235788 200685 235789
rect 200619 235724 200620 235788
rect 200684 235724 200685 235788
rect 200619 235723 200685 235724
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199331 161668 199397 161669
rect 199331 161604 199332 161668
rect 199396 161604 199397 161668
rect 199331 161603 199397 161604
rect 195835 155276 195901 155277
rect 195835 155212 195836 155276
rect 195900 155212 195901 155276
rect 195835 155211 195901 155212
rect 193811 153100 193877 153101
rect 193811 153036 193812 153100
rect 193876 153036 193877 153100
rect 193811 153035 193877 153036
rect 193814 152693 193874 153035
rect 193811 152692 193877 152693
rect 193811 152628 193812 152692
rect 193876 152628 193877 152692
rect 193811 152627 193877 152628
rect 195838 142170 195898 155211
rect 197859 143172 197925 143173
rect 197859 143108 197860 143172
rect 197924 143108 197925 143172
rect 197859 143107 197925 143108
rect 194550 142110 195898 142170
rect 194179 137732 194245 137733
rect 194179 137668 194180 137732
rect 194244 137730 194245 137732
rect 194550 137730 194610 142110
rect 197862 140589 197922 143107
rect 199794 143035 200414 164898
rect 197859 140588 197925 140589
rect 197859 140524 197860 140588
rect 197924 140524 197925 140588
rect 197859 140523 197925 140524
rect 196571 140452 196637 140453
rect 196571 140388 196572 140452
rect 196636 140388 196637 140452
rect 196571 140387 196637 140388
rect 194244 137670 194610 137730
rect 194244 137668 194245 137670
rect 194179 137667 194245 137668
rect 192707 128484 192773 128485
rect 192707 128420 192708 128484
rect 192772 128420 192773 128484
rect 192707 128419 192773 128420
rect 191603 118012 191669 118013
rect 191603 117948 191604 118012
rect 191668 117948 191669 118012
rect 191603 117947 191669 117948
rect 191051 96932 191117 96933
rect 191051 96868 191052 96932
rect 191116 96868 191117 96932
rect 191051 96867 191117 96868
rect 191054 88093 191114 96867
rect 191051 88092 191117 88093
rect 191051 88028 191052 88092
rect 191116 88028 191117 88092
rect 191051 88027 191117 88028
rect 189234 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 189854 82894
rect 189234 82574 189854 82658
rect 189234 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 189854 82574
rect 189234 46894 189854 82338
rect 192710 80749 192770 128419
rect 193443 94756 193509 94757
rect 193443 94692 193444 94756
rect 193508 94692 193509 94756
rect 193443 94691 193509 94692
rect 193446 92581 193506 94691
rect 193811 94212 193877 94213
rect 193811 94148 193812 94212
rect 193876 94148 193877 94212
rect 193811 94147 193877 94148
rect 193443 92580 193509 92581
rect 193443 92516 193444 92580
rect 193508 92516 193509 92580
rect 193443 92515 193509 92516
rect 192954 86614 193574 90782
rect 192954 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 193574 86614
rect 192954 86294 193574 86378
rect 192954 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 193574 86294
rect 192707 80748 192773 80749
rect 192707 80684 192708 80748
rect 192772 80684 192773 80748
rect 192707 80683 192773 80684
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 50614 193574 86058
rect 193814 63477 193874 94147
rect 196574 76533 196634 140387
rect 196571 76532 196637 76533
rect 196571 76468 196572 76532
rect 196636 76468 196637 76532
rect 196571 76467 196637 76468
rect 193811 63476 193877 63477
rect 193811 63412 193812 63476
rect 193876 63412 193877 63476
rect 193811 63411 193877 63412
rect 193814 60621 193874 63411
rect 193811 60620 193877 60621
rect 193811 60556 193812 60620
rect 193876 60556 193877 60620
rect 193811 60555 193877 60556
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 197862 7581 197922 140523
rect 199388 111454 199708 111486
rect 199388 111218 199430 111454
rect 199666 111218 199708 111454
rect 199388 111134 199708 111218
rect 199388 110898 199430 111134
rect 199666 110898 199708 111134
rect 199388 110866 199708 110898
rect 201542 92853 201602 237899
rect 203011 214708 203077 214709
rect 203011 214644 203012 214708
rect 203076 214644 203077 214708
rect 203011 214643 203077 214644
rect 201539 92852 201605 92853
rect 201539 92788 201540 92852
rect 201604 92788 201605 92852
rect 201539 92787 201605 92788
rect 203014 92445 203074 214643
rect 203514 205174 204134 239592
rect 203514 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 204134 205174
rect 203514 204854 204134 204938
rect 203514 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 204134 204854
rect 203514 169174 204134 204618
rect 204302 202197 204362 301411
rect 205403 237964 205469 237965
rect 205403 237900 205404 237964
rect 205468 237900 205469 237964
rect 205403 237899 205469 237900
rect 204299 202196 204365 202197
rect 204299 202132 204300 202196
rect 204364 202132 204365 202196
rect 204299 202131 204365 202132
rect 203514 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 204134 169174
rect 203514 168854 204134 168938
rect 203514 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 204134 168854
rect 203514 143035 204134 168618
rect 204264 129454 204584 129486
rect 204264 129218 204306 129454
rect 204542 129218 204584 129454
rect 204264 129134 204584 129218
rect 204264 128898 204306 129134
rect 204542 128898 204584 129134
rect 204264 128866 204584 128898
rect 205406 92853 205466 237899
rect 206142 228445 206202 307667
rect 207234 303592 207854 316338
rect 207059 301476 207125 301477
rect 207059 301412 207060 301476
rect 207124 301412 207125 301476
rect 207059 301411 207125 301412
rect 206139 228444 206205 228445
rect 206139 228380 206140 228444
rect 206204 228380 206205 228444
rect 206139 228379 206205 228380
rect 207062 225589 207122 301411
rect 208350 241501 208410 385595
rect 210954 356614 211574 388356
rect 216443 384028 216509 384029
rect 216443 383964 216444 384028
rect 216508 383964 216509 384028
rect 216443 383963 216509 383964
rect 215155 364988 215221 364989
rect 215155 364924 215156 364988
rect 215220 364924 215221 364988
rect 215155 364923 215221 364924
rect 210954 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 211574 356614
rect 210954 356294 211574 356378
rect 210954 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 211574 356294
rect 210954 320614 211574 356058
rect 210954 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 211574 320614
rect 210954 320294 211574 320378
rect 210954 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 211574 320294
rect 210954 303592 211574 320058
rect 213683 303788 213749 303789
rect 213683 303724 213684 303788
rect 213748 303724 213749 303788
rect 213683 303723 213749 303724
rect 211659 303652 211725 303653
rect 211659 303588 211660 303652
rect 211724 303588 211725 303652
rect 211659 303587 211725 303588
rect 210555 301476 210621 301477
rect 210555 301412 210556 301476
rect 210620 301412 210621 301476
rect 210555 301411 210621 301412
rect 208347 241500 208413 241501
rect 208347 241436 208348 241500
rect 208412 241436 208413 241500
rect 208347 241435 208413 241436
rect 210371 240956 210437 240957
rect 210371 240892 210372 240956
rect 210436 240892 210437 240956
rect 210371 240891 210437 240892
rect 207059 225588 207125 225589
rect 207059 225524 207060 225588
rect 207124 225524 207125 225588
rect 207059 225523 207125 225524
rect 207234 208894 207854 239592
rect 208347 232524 208413 232525
rect 208347 232460 208348 232524
rect 208412 232460 208413 232524
rect 208347 232459 208413 232460
rect 207234 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 207854 208894
rect 207234 208574 207854 208658
rect 207234 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 207854 208574
rect 207234 172894 207854 208338
rect 207234 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 207854 172894
rect 207234 172574 207854 172658
rect 207234 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 207854 172574
rect 207234 143035 207854 172338
rect 208350 92853 208410 232459
rect 209140 111454 209460 111486
rect 209140 111218 209182 111454
rect 209418 111218 209460 111454
rect 209140 111134 209460 111218
rect 209140 110898 209182 111134
rect 209418 110898 209460 111134
rect 209140 110866 209460 110898
rect 210374 93870 210434 240891
rect 210558 240141 210618 301411
rect 210555 240140 210621 240141
rect 210555 240076 210556 240140
rect 210620 240076 210621 240140
rect 210555 240075 210621 240076
rect 210954 212614 211574 239592
rect 211662 229125 211722 303587
rect 213136 273454 213456 273486
rect 213136 273218 213178 273454
rect 213414 273218 213456 273454
rect 213136 273134 213456 273218
rect 213136 272898 213178 273134
rect 213414 272898 213456 273134
rect 213136 272866 213456 272898
rect 211659 229124 211725 229125
rect 211659 229060 211660 229124
rect 211724 229060 211725 229124
rect 211659 229059 211725 229060
rect 212579 218108 212645 218109
rect 212579 218044 212580 218108
rect 212644 218044 212645 218108
rect 212579 218043 212645 218044
rect 210954 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 211574 212614
rect 210954 212294 211574 212378
rect 210954 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 211574 212294
rect 210954 176614 211574 212058
rect 210954 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 211574 176614
rect 210954 176294 211574 176378
rect 210954 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 211574 176294
rect 210954 143035 211574 176058
rect 211659 143852 211725 143853
rect 211659 143788 211660 143852
rect 211724 143788 211725 143852
rect 211659 143787 211725 143788
rect 210006 93810 210434 93870
rect 210006 92853 210066 93810
rect 211662 93397 211722 143787
rect 211659 93396 211725 93397
rect 211659 93332 211660 93396
rect 211724 93332 211725 93396
rect 211659 93331 211725 93332
rect 205403 92852 205469 92853
rect 205403 92788 205404 92852
rect 205468 92788 205469 92852
rect 205403 92787 205469 92788
rect 208347 92852 208413 92853
rect 208347 92788 208348 92852
rect 208412 92788 208413 92852
rect 208347 92787 208413 92788
rect 210003 92852 210069 92853
rect 210003 92788 210004 92852
rect 210068 92788 210069 92852
rect 210003 92787 210069 92788
rect 203011 92444 203077 92445
rect 203011 92380 203012 92444
rect 203076 92380 203077 92444
rect 203011 92379 203077 92380
rect 204851 92036 204917 92037
rect 204851 91972 204852 92036
rect 204916 91972 204917 92036
rect 204851 91971 204917 91972
rect 199794 57454 200414 90782
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 197859 7580 197925 7581
rect 197859 7516 197860 7580
rect 197924 7516 197925 7580
rect 197859 7515 197925 7516
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 61174 204134 90782
rect 204854 88093 204914 91971
rect 204851 88092 204917 88093
rect 204851 88028 204852 88092
rect 204916 88028 204917 88092
rect 204851 88027 204917 88028
rect 203514 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 204134 61174
rect 203514 60854 204134 60938
rect 203514 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 204134 60854
rect 203514 25174 204134 60618
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 64894 207854 90782
rect 210006 82517 210066 92787
rect 212582 92445 212642 218043
rect 213686 167653 213746 303723
rect 214419 302292 214485 302293
rect 214419 302228 214420 302292
rect 214484 302228 214485 302292
rect 214419 302227 214485 302228
rect 214422 180029 214482 302227
rect 215158 241501 215218 364923
rect 215891 301476 215957 301477
rect 215891 301412 215892 301476
rect 215956 301412 215957 301476
rect 215891 301411 215957 301412
rect 215155 241500 215221 241501
rect 215155 241436 215156 241500
rect 215220 241436 215221 241500
rect 215155 241435 215221 241436
rect 215894 211853 215954 301411
rect 216446 240005 216506 383963
rect 217794 363454 218414 388356
rect 221514 367174 222134 388356
rect 221514 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 222134 367174
rect 221514 366854 222134 366938
rect 221514 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 222134 366854
rect 218651 366348 218717 366349
rect 218651 366284 218652 366348
rect 218716 366284 218717 366348
rect 218651 366283 218717 366284
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217179 322964 217245 322965
rect 217179 322900 217180 322964
rect 217244 322900 217245 322964
rect 217179 322899 217245 322900
rect 217182 306390 217242 322899
rect 217182 306330 217610 306390
rect 217550 303925 217610 306330
rect 217547 303924 217613 303925
rect 217547 303860 217548 303924
rect 217612 303860 217613 303924
rect 217547 303859 217613 303860
rect 216443 240004 216509 240005
rect 216443 239940 216444 240004
rect 216508 239940 216509 240004
rect 216443 239939 216509 239940
rect 216446 238101 216506 239939
rect 216443 238100 216509 238101
rect 216443 238036 216444 238100
rect 216508 238036 216509 238100
rect 216443 238035 216509 238036
rect 215891 211852 215957 211853
rect 215891 211788 215892 211852
rect 215956 211788 215957 211852
rect 215891 211787 215957 211788
rect 215339 210356 215405 210357
rect 215339 210292 215340 210356
rect 215404 210292 215405 210356
rect 215339 210291 215405 210292
rect 214419 180028 214485 180029
rect 214419 179964 214420 180028
rect 214484 179964 214485 180028
rect 214419 179963 214485 179964
rect 213683 167652 213749 167653
rect 213683 167588 213684 167652
rect 213748 167588 213749 167652
rect 213683 167587 213749 167588
rect 214016 129454 214336 129486
rect 214016 129218 214058 129454
rect 214294 129218 214336 129454
rect 214016 129134 214336 129218
rect 214016 128898 214058 129134
rect 214294 128898 214336 129134
rect 214016 128866 214336 128898
rect 215342 92717 215402 210291
rect 217550 155277 217610 303859
rect 217794 303592 218414 326898
rect 218654 241501 218714 366283
rect 221227 360908 221293 360909
rect 221227 360844 221228 360908
rect 221292 360844 221293 360908
rect 221227 360843 221293 360844
rect 220491 305284 220557 305285
rect 220491 305220 220492 305284
rect 220556 305220 220557 305284
rect 220491 305219 220557 305220
rect 219203 301476 219269 301477
rect 219203 301412 219204 301476
rect 219268 301412 219269 301476
rect 219203 301411 219269 301412
rect 218651 241500 218717 241501
rect 218651 241436 218652 241500
rect 218716 241436 218717 241500
rect 218651 241435 218717 241436
rect 217794 219454 218414 239592
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217547 155276 217613 155277
rect 217547 155212 217548 155276
rect 217612 155212 217613 155276
rect 217547 155211 217613 155212
rect 217794 147454 218414 182898
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 219206 147117 219266 301411
rect 220494 177445 220554 305219
rect 220859 301884 220925 301885
rect 220859 301820 220860 301884
rect 220924 301820 220925 301884
rect 220859 301819 220925 301820
rect 220675 227764 220741 227765
rect 220675 227700 220676 227764
rect 220740 227700 220741 227764
rect 220675 227699 220741 227700
rect 220491 177444 220557 177445
rect 220491 177380 220492 177444
rect 220556 177380 220557 177444
rect 220491 177379 220557 177380
rect 219203 147116 219269 147117
rect 219203 147052 219204 147116
rect 219268 147052 219269 147116
rect 219203 147051 219269 147052
rect 217794 143035 218414 146898
rect 218892 111454 219212 111486
rect 218892 111218 218934 111454
rect 219170 111218 219212 111454
rect 218892 111134 219212 111218
rect 218892 110898 218934 111134
rect 219170 110898 219212 111134
rect 218892 110866 219212 110898
rect 220678 92853 220738 227699
rect 220862 224229 220922 301819
rect 221230 241501 221290 360843
rect 221514 331174 222134 366618
rect 221514 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 222134 331174
rect 221514 330854 222134 330938
rect 221514 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 222134 330854
rect 221514 303592 222134 330618
rect 225234 370894 225854 388356
rect 225234 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 225854 370894
rect 225234 370574 225854 370658
rect 225234 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 225854 370574
rect 225234 334894 225854 370338
rect 225234 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 225854 334894
rect 225234 334574 225854 334658
rect 225234 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 225854 334574
rect 224171 307732 224237 307733
rect 224171 307668 224172 307732
rect 224236 307668 224237 307732
rect 224171 307667 224237 307668
rect 222331 301612 222397 301613
rect 222331 301548 222332 301612
rect 222396 301548 222397 301612
rect 222331 301547 222397 301548
rect 221227 241500 221293 241501
rect 221227 241436 221228 241500
rect 221292 241436 221293 241500
rect 221227 241435 221293 241436
rect 220859 224228 220925 224229
rect 220859 224164 220860 224228
rect 220924 224164 220925 224228
rect 220859 224163 220925 224164
rect 221514 223174 222134 239592
rect 221514 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 222134 223174
rect 221514 222854 222134 222938
rect 221514 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 222134 222854
rect 221514 187174 222134 222618
rect 222334 203557 222394 301547
rect 222699 301476 222765 301477
rect 222699 301412 222700 301476
rect 222764 301412 222765 301476
rect 222699 301411 222765 301412
rect 223619 301476 223685 301477
rect 223619 301412 223620 301476
rect 223684 301412 223685 301476
rect 223619 301411 223685 301412
rect 222702 230349 222762 301411
rect 222699 230348 222765 230349
rect 222699 230284 222700 230348
rect 222764 230284 222765 230348
rect 222699 230283 222765 230284
rect 223435 229940 223501 229941
rect 223435 229876 223436 229940
rect 223500 229876 223501 229940
rect 223435 229875 223501 229876
rect 222331 203556 222397 203557
rect 222331 203492 222332 203556
rect 222396 203492 222397 203556
rect 222331 203491 222397 203492
rect 221514 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 222134 187174
rect 221514 186854 222134 186938
rect 221514 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 222134 186854
rect 221514 151174 222134 186618
rect 221514 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 222134 151174
rect 221514 150854 222134 150938
rect 221514 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 222134 150854
rect 221514 143035 222134 150618
rect 223438 92989 223498 229875
rect 223622 200701 223682 301411
rect 224174 239869 224234 307667
rect 225234 303592 225854 334338
rect 228954 374614 229574 388356
rect 228954 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 229574 374614
rect 228954 374294 229574 374378
rect 228954 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 229574 374294
rect 228954 338614 229574 374058
rect 228954 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 229574 338614
rect 228954 338294 229574 338378
rect 228954 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 229574 338294
rect 226195 305148 226261 305149
rect 226195 305084 226196 305148
rect 226260 305084 226261 305148
rect 226195 305083 226261 305084
rect 224907 301476 224973 301477
rect 224907 301412 224908 301476
rect 224972 301412 224973 301476
rect 224907 301411 224973 301412
rect 224171 239868 224237 239869
rect 224171 239804 224172 239868
rect 224236 239804 224237 239868
rect 224171 239803 224237 239804
rect 223619 200700 223685 200701
rect 223619 200636 223620 200700
rect 223684 200636 223685 200700
rect 223619 200635 223685 200636
rect 224910 197981 224970 301411
rect 226198 241501 226258 305083
rect 228954 303592 229574 338058
rect 235794 381454 236414 388356
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 239514 385174 240134 388356
rect 239514 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 240134 385174
rect 239514 384854 240134 384938
rect 239514 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 240134 384854
rect 236499 370700 236565 370701
rect 236499 370636 236500 370700
rect 236564 370636 236565 370700
rect 236499 370635 236565 370636
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 230243 306508 230309 306509
rect 230243 306444 230244 306508
rect 230308 306444 230309 306508
rect 230243 306443 230309 306444
rect 226563 301612 226629 301613
rect 226563 301548 226564 301612
rect 226628 301548 226629 301612
rect 226563 301547 226629 301548
rect 226195 241500 226261 241501
rect 226195 241436 226196 241500
rect 226260 241436 226261 241500
rect 226195 241435 226261 241436
rect 225234 226894 225854 239592
rect 226566 229805 226626 301547
rect 226747 301476 226813 301477
rect 226747 301412 226748 301476
rect 226812 301412 226813 301476
rect 226747 301411 226813 301412
rect 227667 301476 227733 301477
rect 227667 301412 227668 301476
rect 227732 301412 227733 301476
rect 227667 301411 227733 301412
rect 229691 301476 229757 301477
rect 229691 301412 229692 301476
rect 229756 301412 229757 301476
rect 229691 301411 229757 301412
rect 226563 229804 226629 229805
rect 226563 229740 226564 229804
rect 226628 229740 226629 229804
rect 226563 229739 226629 229740
rect 225234 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 225854 226894
rect 225234 226574 225854 226658
rect 225234 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 225854 226574
rect 224907 197980 224973 197981
rect 224907 197916 224908 197980
rect 224972 197916 224973 197980
rect 224907 197915 224973 197916
rect 225234 190894 225854 226338
rect 226750 204917 226810 301411
rect 226747 204916 226813 204917
rect 226747 204852 226748 204916
rect 226812 204852 226813 204916
rect 226747 204851 226813 204852
rect 225234 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 225854 190894
rect 225234 190574 225854 190658
rect 225234 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 225854 190574
rect 224907 156228 224973 156229
rect 224907 156164 224908 156228
rect 224972 156164 224973 156228
rect 224907 156163 224973 156164
rect 223619 147796 223685 147797
rect 223619 147732 223620 147796
rect 223684 147732 223685 147796
rect 223619 147731 223685 147732
rect 223622 132510 223682 147731
rect 224723 142220 224789 142221
rect 224723 142156 224724 142220
rect 224788 142156 224789 142220
rect 224723 142155 224789 142156
rect 224726 135965 224786 142155
rect 224723 135964 224789 135965
rect 224723 135900 224724 135964
rect 224788 135900 224789 135964
rect 224723 135899 224789 135900
rect 223622 132450 224418 132510
rect 224358 124133 224418 132450
rect 224910 130661 224970 156163
rect 225234 154894 225854 190338
rect 227670 189685 227730 301411
rect 228496 291454 228816 291486
rect 228496 291218 228538 291454
rect 228774 291218 228816 291454
rect 228496 291134 228816 291218
rect 228496 290898 228538 291134
rect 228774 290898 228816 291134
rect 228496 290866 228816 290898
rect 228496 255454 228816 255486
rect 228496 255218 228538 255454
rect 228774 255218 228816 255454
rect 228496 255134 228816 255218
rect 228496 254898 228538 255134
rect 228774 254898 228816 255134
rect 228496 254866 228816 254898
rect 229694 240141 229754 301411
rect 229691 240140 229757 240141
rect 229691 240076 229692 240140
rect 229756 240076 229757 240140
rect 229691 240075 229757 240076
rect 228954 230614 229574 239592
rect 230246 238781 230306 306443
rect 235794 303592 236414 308898
rect 230427 301612 230493 301613
rect 230427 301548 230428 301612
rect 230492 301548 230493 301612
rect 230427 301547 230493 301548
rect 234659 301612 234725 301613
rect 234659 301548 234660 301612
rect 234724 301548 234725 301612
rect 234659 301547 234725 301548
rect 230243 238780 230309 238781
rect 230243 238770 230244 238780
rect 229878 238716 230244 238770
rect 230308 238716 230309 238780
rect 229878 238715 230309 238716
rect 229878 238710 230306 238715
rect 229878 235653 229938 238710
rect 229875 235652 229941 235653
rect 229875 235588 229876 235652
rect 229940 235588 229941 235652
rect 229875 235587 229941 235588
rect 228954 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 229574 230614
rect 228954 230294 229574 230378
rect 228954 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 229574 230294
rect 228954 194614 229574 230058
rect 228954 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 229574 194614
rect 228954 194294 229574 194378
rect 228954 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 229574 194294
rect 227667 189684 227733 189685
rect 227667 189620 227668 189684
rect 227732 189620 227733 189684
rect 227667 189619 227733 189620
rect 228219 189684 228285 189685
rect 228219 189620 228220 189684
rect 228284 189620 228285 189684
rect 228219 189619 228285 189620
rect 225234 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 225854 154894
rect 225234 154574 225854 154658
rect 225234 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 225854 154574
rect 226379 154596 226445 154597
rect 226379 154532 226380 154596
rect 226444 154532 226445 154596
rect 226379 154531 226445 154532
rect 225234 143035 225854 154338
rect 224907 130660 224973 130661
rect 224907 130596 224908 130660
rect 224972 130596 224973 130660
rect 224907 130595 224973 130596
rect 224355 124132 224421 124133
rect 224355 124068 224356 124132
rect 224420 124068 224421 124132
rect 224355 124067 224421 124068
rect 226382 107813 226442 154531
rect 228222 151830 228282 189619
rect 227670 151770 228282 151830
rect 228954 158614 229574 194058
rect 228954 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 229574 158614
rect 228954 158294 229574 158378
rect 228954 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 229574 158294
rect 227670 149293 227730 151770
rect 227667 149292 227733 149293
rect 227667 149228 227668 149292
rect 227732 149228 227733 149292
rect 227667 149227 227733 149228
rect 226931 146300 226997 146301
rect 226931 146236 226932 146300
rect 226996 146236 226997 146300
rect 226931 146235 226997 146236
rect 226934 136373 226994 146235
rect 226931 136372 226997 136373
rect 226931 136308 226932 136372
rect 226996 136308 226997 136372
rect 226931 136307 226997 136308
rect 227670 135557 227730 149227
rect 227667 135556 227733 135557
rect 227667 135492 227668 135556
rect 227732 135492 227733 135556
rect 227667 135491 227733 135492
rect 228954 122614 229574 158058
rect 228954 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 229574 122614
rect 228954 122294 229574 122378
rect 228954 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 229574 122294
rect 226563 108628 226629 108629
rect 226563 108564 226564 108628
rect 226628 108564 226629 108628
rect 226563 108563 226629 108564
rect 226379 107812 226445 107813
rect 226379 107748 226380 107812
rect 226444 107748 226445 107812
rect 226379 107747 226445 107748
rect 226566 103530 226626 108563
rect 226382 103470 226626 103530
rect 224723 97476 224789 97477
rect 224723 97412 224724 97476
rect 224788 97412 224789 97476
rect 224723 97411 224789 97412
rect 224355 94756 224421 94757
rect 224355 94692 224356 94756
rect 224420 94692 224421 94756
rect 224355 94691 224421 94692
rect 223435 92988 223501 92989
rect 223435 92924 223436 92988
rect 223500 92924 223501 92988
rect 223435 92923 223501 92924
rect 224358 92853 224418 94691
rect 224726 93397 224786 97411
rect 224907 95164 224973 95165
rect 224907 95100 224908 95164
rect 224972 95100 224973 95164
rect 224907 95099 224973 95100
rect 224723 93396 224789 93397
rect 224723 93332 224724 93396
rect 224788 93332 224789 93396
rect 224723 93331 224789 93332
rect 220675 92852 220741 92853
rect 220675 92788 220676 92852
rect 220740 92788 220741 92852
rect 220675 92787 220741 92788
rect 224355 92852 224421 92853
rect 224355 92788 224356 92852
rect 224420 92788 224421 92852
rect 224355 92787 224421 92788
rect 215339 92716 215405 92717
rect 215339 92652 215340 92716
rect 215404 92652 215405 92716
rect 215339 92651 215405 92652
rect 212579 92444 212645 92445
rect 212579 92380 212580 92444
rect 212644 92380 212645 92444
rect 212579 92379 212645 92380
rect 212582 92037 212642 92379
rect 212579 92036 212645 92037
rect 212579 91972 212580 92036
rect 212644 91972 212645 92036
rect 212579 91971 212645 91972
rect 210003 82516 210069 82517
rect 210003 82452 210004 82516
rect 210068 82452 210069 82516
rect 210003 82451 210069 82452
rect 207234 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 207854 64894
rect 207234 64574 207854 64658
rect 207234 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 207854 64574
rect 207234 28894 207854 64338
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 68614 211574 90782
rect 210954 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 211574 68614
rect 210954 68294 211574 68378
rect 210954 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 211574 68294
rect 210954 32614 211574 68058
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 75454 218414 90782
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 79174 222134 90782
rect 224910 87957 224970 95099
rect 224907 87956 224973 87957
rect 224907 87892 224908 87956
rect 224972 87892 224973 87956
rect 224907 87891 224973 87892
rect 221514 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 222134 79174
rect 221514 78854 222134 78938
rect 221514 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 222134 78854
rect 221514 43174 222134 78618
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 82894 225854 90782
rect 225234 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 225854 82894
rect 225234 82574 225854 82658
rect 226382 82653 226442 103470
rect 228954 86614 229574 122058
rect 228954 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 229574 86614
rect 228954 86294 229574 86378
rect 228954 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 229574 86294
rect 226379 82652 226445 82653
rect 226379 82588 226380 82652
rect 226444 82588 226445 82652
rect 226379 82587 226445 82588
rect 225234 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 225854 82574
rect 225234 46894 225854 82338
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 50614 229574 86058
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 230430 6221 230490 301547
rect 230611 301476 230677 301477
rect 230611 301412 230612 301476
rect 230676 301412 230677 301476
rect 230611 301411 230677 301412
rect 232083 301476 232149 301477
rect 232083 301412 232084 301476
rect 232148 301412 232149 301476
rect 232083 301411 232149 301412
rect 232267 301476 232333 301477
rect 232267 301412 232268 301476
rect 232332 301412 232333 301476
rect 232267 301411 232333 301412
rect 233187 301476 233253 301477
rect 233187 301412 233188 301476
rect 233252 301412 233253 301476
rect 233187 301411 233253 301412
rect 233555 301476 233621 301477
rect 233555 301412 233556 301476
rect 233620 301412 233621 301476
rect 233555 301411 233621 301412
rect 230614 73813 230674 301411
rect 230611 73812 230677 73813
rect 230611 73748 230612 73812
rect 230676 73748 230677 73812
rect 230611 73747 230677 73748
rect 232086 69597 232146 301411
rect 232083 69596 232149 69597
rect 232083 69532 232084 69596
rect 232148 69532 232149 69596
rect 232083 69531 232149 69532
rect 232270 14517 232330 301411
rect 233190 61437 233250 301411
rect 233187 61436 233253 61437
rect 233187 61372 233188 61436
rect 233252 61372 233253 61436
rect 233187 61371 233253 61372
rect 233558 48925 233618 301411
rect 234662 54501 234722 301547
rect 234843 301476 234909 301477
rect 234843 301412 234844 301476
rect 234908 301412 234909 301476
rect 234843 301411 234909 301412
rect 234846 240141 234906 301411
rect 236502 241501 236562 370635
rect 239514 349174 240134 384618
rect 239514 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 240134 349174
rect 239514 348854 240134 348938
rect 239514 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 240134 348854
rect 238891 337380 238957 337381
rect 238891 337316 238892 337380
rect 238956 337316 238957 337380
rect 238891 337315 238957 337316
rect 237603 301612 237669 301613
rect 237603 301548 237604 301612
rect 237668 301548 237669 301612
rect 237603 301547 237669 301548
rect 236683 301476 236749 301477
rect 236683 301412 236684 301476
rect 236748 301412 236749 301476
rect 236683 301411 236749 301412
rect 236499 241500 236565 241501
rect 236499 241436 236500 241500
rect 236564 241436 236565 241500
rect 236499 241435 236565 241436
rect 234843 240140 234909 240141
rect 234843 240076 234844 240140
rect 234908 240076 234909 240140
rect 234843 240075 234909 240076
rect 235794 237454 236414 239592
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 235794 201454 236414 236898
rect 236686 231165 236746 301411
rect 236683 231164 236749 231165
rect 236683 231100 236684 231164
rect 236748 231100 236749 231164
rect 236683 231099 236749 231100
rect 237606 226949 237666 301547
rect 237787 301476 237853 301477
rect 237787 301412 237788 301476
rect 237852 301412 237853 301476
rect 237787 301411 237853 301412
rect 238523 301476 238589 301477
rect 238523 301412 238524 301476
rect 238588 301412 238589 301476
rect 238523 301411 238589 301412
rect 237603 226948 237669 226949
rect 237603 226884 237604 226948
rect 237668 226884 237669 226948
rect 237603 226883 237669 226884
rect 237790 222733 237850 301411
rect 238526 225725 238586 301411
rect 238894 241501 238954 337315
rect 239514 313174 240134 348618
rect 239514 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 240134 313174
rect 239514 312854 240134 312938
rect 239514 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 240134 312854
rect 239514 303592 240134 312618
rect 241467 305148 241533 305149
rect 241467 305084 241468 305148
rect 241532 305084 241533 305148
rect 241467 305083 241533 305084
rect 241470 305010 241530 305083
rect 241654 305010 241714 452915
rect 243234 452356 243854 460338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 608614 247574 644058
rect 246954 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 247574 608614
rect 246954 608294 247574 608378
rect 246954 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 247574 608294
rect 246954 572614 247574 608058
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 536614 247574 572058
rect 246954 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 247574 536614
rect 246954 536294 247574 536378
rect 246954 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 247574 536294
rect 246954 500614 247574 536058
rect 246954 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 247574 500614
rect 246954 500294 247574 500378
rect 246954 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 247574 500294
rect 246954 464614 247574 500058
rect 246954 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 247574 464614
rect 246954 464294 247574 464378
rect 246954 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 247574 464294
rect 246954 452356 247574 464058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253059 458556 253125 458557
rect 253059 458492 253060 458556
rect 253124 458492 253125 458556
rect 253059 458491 253125 458492
rect 247723 451620 247789 451621
rect 247723 451556 247724 451620
rect 247788 451556 247789 451620
rect 247723 451555 247789 451556
rect 244411 449988 244477 449989
rect 244411 449924 244412 449988
rect 244476 449924 244477 449988
rect 244411 449923 244477 449924
rect 242939 449716 243005 449717
rect 242939 449652 242940 449716
rect 243004 449652 243005 449716
rect 242939 449651 243005 449652
rect 242942 384301 243002 449651
rect 243856 417454 244176 417486
rect 243856 417218 243898 417454
rect 244134 417218 244176 417454
rect 243856 417134 244176 417218
rect 243856 416898 243898 417134
rect 244134 416898 244176 417134
rect 243856 416866 244176 416898
rect 242939 384300 243005 384301
rect 242939 384236 242940 384300
rect 243004 384236 243005 384300
rect 242939 384235 243005 384236
rect 242755 378044 242821 378045
rect 242755 377980 242756 378044
rect 242820 377980 242821 378044
rect 242755 377979 242821 377980
rect 241470 304950 241714 305010
rect 241654 304197 241714 304950
rect 241651 304196 241717 304197
rect 241651 304132 241652 304196
rect 241716 304132 241717 304196
rect 241651 304131 241717 304132
rect 240731 302292 240797 302293
rect 240731 302228 240732 302292
rect 240796 302228 240797 302292
rect 240731 302227 240797 302228
rect 238891 241500 238957 241501
rect 238891 241436 238892 241500
rect 238956 241436 238957 241500
rect 238891 241435 238957 241436
rect 238894 240141 238954 241435
rect 238891 240140 238957 240141
rect 238891 240076 238892 240140
rect 238956 240076 238957 240140
rect 238891 240075 238957 240076
rect 238523 225724 238589 225725
rect 238523 225660 238524 225724
rect 238588 225660 238589 225724
rect 238523 225659 238589 225660
rect 237787 222732 237853 222733
rect 237787 222668 237788 222732
rect 237852 222668 237853 222732
rect 237787 222667 237853 222668
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 165454 236414 200898
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 235794 129454 236414 164898
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 234659 54500 234725 54501
rect 234659 54436 234660 54500
rect 234724 54436 234725 54500
rect 234659 54435 234725 54436
rect 233555 48924 233621 48925
rect 233555 48860 233556 48924
rect 233620 48860 233621 48924
rect 233555 48859 233621 48860
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 232267 14516 232333 14517
rect 232267 14452 232268 14516
rect 232332 14452 232333 14516
rect 232267 14451 232333 14452
rect 230427 6220 230493 6221
rect 230427 6156 230428 6220
rect 230492 6156 230493 6220
rect 230427 6155 230493 6156
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 205174 240134 239592
rect 240734 226949 240794 302227
rect 242758 241501 242818 377979
rect 243234 352894 243854 388356
rect 244414 384437 244474 449923
rect 244411 384436 244477 384437
rect 244411 384372 244412 384436
rect 244476 384372 244477 384436
rect 244411 384371 244477 384372
rect 243234 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 243854 352894
rect 243234 352574 243854 352658
rect 243234 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 243854 352574
rect 243234 316894 243854 352338
rect 243234 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 243854 316894
rect 243234 316574 243854 316658
rect 243234 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 243854 316574
rect 243234 303592 243854 316338
rect 246954 356614 247574 388356
rect 247726 370701 247786 451555
rect 249747 449988 249813 449989
rect 249747 449924 249748 449988
rect 249812 449924 249813 449988
rect 249747 449923 249813 449924
rect 247723 370700 247789 370701
rect 247723 370636 247724 370700
rect 247788 370636 247789 370700
rect 247723 370635 247789 370636
rect 249750 366349 249810 449923
rect 252875 440332 252941 440333
rect 252875 440268 252876 440332
rect 252940 440268 252941 440332
rect 252875 440267 252941 440268
rect 252878 431970 252938 440267
rect 253062 436797 253122 458491
rect 253794 452356 254414 470898
rect 257514 691174 258134 706202
rect 258579 702540 258645 702541
rect 258579 702476 258580 702540
rect 258644 702476 258645 702540
rect 258579 702475 258645 702476
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 547174 258134 582618
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257514 511174 258134 546618
rect 257514 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 258134 511174
rect 257514 510854 258134 510938
rect 257514 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 258134 510854
rect 257514 475174 258134 510618
rect 257514 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 258134 475174
rect 257514 474854 258134 474938
rect 257514 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 258134 474854
rect 256739 450124 256805 450125
rect 256739 450060 256740 450124
rect 256804 450060 256805 450124
rect 256739 450059 256805 450060
rect 253059 436796 253125 436797
rect 253059 436732 253060 436796
rect 253124 436732 253125 436796
rect 253059 436731 253125 436732
rect 252510 431910 252938 431970
rect 249747 366348 249813 366349
rect 249747 366284 249748 366348
rect 249812 366284 249813 366348
rect 249747 366283 249813 366284
rect 246954 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 247574 356614
rect 246954 356294 247574 356378
rect 246954 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 247574 356294
rect 246954 320614 247574 356058
rect 252510 338061 252570 431910
rect 252875 404836 252941 404837
rect 252875 404772 252876 404836
rect 252940 404772 252941 404836
rect 252875 404771 252941 404772
rect 252878 393330 252938 404771
rect 253979 395588 254045 395589
rect 253979 395524 253980 395588
rect 254044 395524 254045 395588
rect 253979 395523 254045 395524
rect 252694 393270 252938 393330
rect 252694 368389 252754 393270
rect 253982 389197 254042 395523
rect 253979 389196 254045 389197
rect 253979 389132 253980 389196
rect 254044 389132 254045 389196
rect 253979 389131 254045 389132
rect 252691 368388 252757 368389
rect 252691 368324 252692 368388
rect 252756 368324 252757 368388
rect 252691 368323 252757 368324
rect 252507 338060 252573 338061
rect 252507 337996 252508 338060
rect 252572 337996 252573 338060
rect 252507 337995 252573 337996
rect 252694 336701 252754 368323
rect 253794 363454 254414 388356
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 252691 336700 252757 336701
rect 252691 336636 252692 336700
rect 252756 336636 252757 336700
rect 252691 336635 252757 336636
rect 252507 334660 252573 334661
rect 252507 334596 252508 334660
rect 252572 334596 252573 334660
rect 252507 334595 252573 334596
rect 252323 328404 252389 328405
rect 252323 328340 252324 328404
rect 252388 328340 252389 328404
rect 252323 328339 252389 328340
rect 252326 327181 252386 328339
rect 252323 327180 252389 327181
rect 252323 327116 252324 327180
rect 252388 327116 252389 327180
rect 252323 327115 252389 327116
rect 246954 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 247574 320614
rect 246954 320294 247574 320378
rect 246954 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 247574 320294
rect 246954 303592 247574 320058
rect 252326 302250 252386 327115
rect 252510 306390 252570 334595
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 252510 306330 252938 306390
rect 252878 302250 252938 306330
rect 253794 303592 254414 326898
rect 256742 309501 256802 450059
rect 257514 439174 258134 474618
rect 258582 462909 258642 702475
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 550894 261854 586338
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 514894 261854 550338
rect 261234 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 261854 514894
rect 261234 514574 261854 514658
rect 261234 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 261854 514574
rect 261234 478894 261854 514338
rect 261234 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 261854 478894
rect 261234 478574 261854 478658
rect 261234 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 261854 478574
rect 258579 462908 258645 462909
rect 258579 462844 258580 462908
rect 258644 462844 258645 462908
rect 258579 462843 258645 462844
rect 258582 451290 258642 462843
rect 258398 451230 258642 451290
rect 258398 442101 258458 451230
rect 261234 442894 261854 478338
rect 261234 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 261854 442894
rect 261234 442574 261854 442658
rect 261234 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 261854 442574
rect 258395 442100 258461 442101
rect 258395 442036 258396 442100
rect 258460 442036 258461 442100
rect 258395 442035 258461 442036
rect 257514 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 258134 439174
rect 257514 438854 258134 438938
rect 257514 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 258134 438854
rect 257514 403174 258134 438618
rect 257514 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 258134 403174
rect 257514 402854 258134 402938
rect 257514 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 258134 402854
rect 257514 367174 258134 402618
rect 261234 406894 261854 442338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 554614 265574 590058
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 518614 265574 554058
rect 264954 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 265574 518614
rect 264954 518294 265574 518378
rect 264954 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 265574 518294
rect 264954 482614 265574 518058
rect 264954 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 265574 482614
rect 264954 482294 265574 482378
rect 264954 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 265574 482294
rect 264954 446614 265574 482058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 269067 465220 269133 465221
rect 269067 465156 269068 465220
rect 269132 465156 269133 465220
rect 269067 465155 269133 465156
rect 267779 455700 267845 455701
rect 267779 455636 267780 455700
rect 267844 455636 267845 455700
rect 267779 455635 267845 455636
rect 266491 454204 266557 454205
rect 266491 454140 266492 454204
rect 266556 454140 266557 454204
rect 266491 454139 266557 454140
rect 264954 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 265574 446614
rect 264954 446294 265574 446378
rect 264954 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 265574 446294
rect 262259 424284 262325 424285
rect 262259 424220 262260 424284
rect 262324 424220 262325 424284
rect 262259 424219 262325 424220
rect 261234 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 261854 406894
rect 261234 406574 261854 406658
rect 261234 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 261854 406574
rect 258395 375324 258461 375325
rect 258395 375260 258396 375324
rect 258460 375260 258461 375324
rect 258395 375259 258461 375260
rect 257514 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 258134 367174
rect 257514 366854 258134 366938
rect 257514 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 258134 366854
rect 257514 331174 258134 366618
rect 257514 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 258134 331174
rect 257514 330854 258134 330938
rect 257514 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 258134 330854
rect 256739 309500 256805 309501
rect 256739 309436 256740 309500
rect 256804 309436 256805 309500
rect 256739 309435 256805 309436
rect 255267 307052 255333 307053
rect 255267 306988 255268 307052
rect 255332 306988 255333 307052
rect 255267 306987 255333 306988
rect 252326 302190 252570 302250
rect 252878 302190 253122 302250
rect 245883 301612 245949 301613
rect 245883 301548 245884 301612
rect 245948 301548 245949 301612
rect 245883 301547 245949 301548
rect 242939 301476 243005 301477
rect 242939 301412 242940 301476
rect 243004 301412 243005 301476
rect 242939 301411 243005 301412
rect 245515 301476 245581 301477
rect 245515 301412 245516 301476
rect 245580 301412 245581 301476
rect 245515 301411 245581 301412
rect 242755 241500 242821 241501
rect 242755 241436 242756 241500
rect 242820 241436 242821 241500
rect 242755 241435 242821 241436
rect 240731 226948 240797 226949
rect 240731 226884 240732 226948
rect 240796 226884 240797 226948
rect 240731 226883 240797 226884
rect 239514 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 240134 205174
rect 239514 204854 240134 204938
rect 239514 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 240134 204854
rect 239514 169174 240134 204618
rect 242942 178669 243002 301411
rect 243856 273454 244176 273486
rect 243856 273218 243898 273454
rect 244134 273218 244176 273454
rect 243856 273134 244176 273218
rect 243856 272898 243898 273134
rect 244134 272898 244176 273134
rect 243856 272866 244176 272898
rect 245518 241501 245578 301411
rect 245886 292590 245946 301547
rect 247723 301476 247789 301477
rect 247723 301412 247724 301476
rect 247788 301412 247789 301476
rect 247723 301411 247789 301412
rect 245702 292530 245946 292590
rect 245515 241500 245581 241501
rect 245515 241436 245516 241500
rect 245580 241436 245581 241500
rect 245515 241435 245581 241436
rect 243234 208894 243854 239592
rect 245702 237965 245762 292530
rect 245699 237964 245765 237965
rect 245699 237900 245700 237964
rect 245764 237900 245765 237964
rect 245699 237899 245765 237900
rect 243234 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 243854 208894
rect 243234 208574 243854 208658
rect 243234 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 243854 208574
rect 242939 178668 243005 178669
rect 242939 178604 242940 178668
rect 243004 178604 243005 178668
rect 242939 178603 243005 178604
rect 239514 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 240134 169174
rect 239514 168854 240134 168938
rect 239514 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 240134 168854
rect 239514 133174 240134 168618
rect 239514 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 240134 133174
rect 239514 132854 240134 132938
rect 239514 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 240134 132854
rect 239514 97174 240134 132618
rect 239514 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 240134 97174
rect 239514 96854 240134 96938
rect 239514 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 240134 96854
rect 239514 61174 240134 96618
rect 239514 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 240134 61174
rect 239514 60854 240134 60938
rect 239514 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 240134 60854
rect 239514 25174 240134 60618
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 172894 243854 208338
rect 243234 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 243854 172894
rect 243234 172574 243854 172658
rect 243234 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 243854 172574
rect 243234 136894 243854 172338
rect 243234 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 243854 136894
rect 243234 136574 243854 136658
rect 243234 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 243854 136574
rect 243234 100894 243854 136338
rect 243234 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 243854 100894
rect 243234 100574 243854 100658
rect 243234 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 243854 100574
rect 243234 64894 243854 100338
rect 243234 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 243854 64894
rect 243234 64574 243854 64658
rect 243234 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 243854 64574
rect 243234 28894 243854 64338
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 212614 247574 239592
rect 246954 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 247574 212614
rect 246954 212294 247574 212378
rect 246954 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 247574 212294
rect 246954 176614 247574 212058
rect 246954 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 247574 176614
rect 246954 176294 247574 176378
rect 246954 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 247574 176294
rect 246954 140614 247574 176058
rect 246954 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 247574 140614
rect 246954 140294 247574 140378
rect 246954 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 247574 140294
rect 246954 104614 247574 140058
rect 246954 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 247574 104614
rect 246954 104294 247574 104378
rect 246954 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 247574 104294
rect 246954 68614 247574 104058
rect 246954 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 247574 68614
rect 246954 68294 247574 68378
rect 246954 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 247574 68294
rect 246954 32614 247574 68058
rect 247726 66197 247786 301411
rect 252510 300930 252570 302190
rect 252510 300870 252938 300930
rect 252878 300661 252938 300870
rect 252875 300660 252941 300661
rect 252875 300596 252876 300660
rect 252940 300596 252941 300660
rect 252875 300595 252941 300596
rect 253062 292590 253122 302190
rect 255270 295901 255330 306987
rect 255267 295900 255333 295901
rect 255267 295836 255268 295900
rect 255332 295836 255333 295900
rect 255267 295835 255333 295836
rect 252878 292530 253122 292590
rect 252878 289509 252938 292530
rect 252875 289508 252941 289509
rect 252875 289444 252876 289508
rect 252940 289444 252941 289508
rect 252875 289443 252941 289444
rect 256742 275637 256802 309435
rect 257514 295174 258134 330618
rect 258398 306390 258458 375259
rect 261234 370894 261854 406338
rect 261234 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 261854 370894
rect 261234 370574 261854 370658
rect 261234 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 261854 370574
rect 261234 334894 261854 370338
rect 261234 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 261854 334894
rect 261234 334574 261854 334658
rect 261234 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 261854 334574
rect 260971 331804 261037 331805
rect 260971 331740 260972 331804
rect 261036 331740 261037 331804
rect 260971 331739 261037 331740
rect 260051 316572 260117 316573
rect 260051 316508 260052 316572
rect 260116 316508 260117 316572
rect 260051 316507 260117 316508
rect 259499 313988 259565 313989
rect 259499 313924 259500 313988
rect 259564 313924 259565 313988
rect 259499 313923 259565 313924
rect 258398 306330 258826 306390
rect 258395 301476 258461 301477
rect 258395 301412 258396 301476
rect 258460 301412 258461 301476
rect 258395 301411 258461 301412
rect 258398 300930 258458 301411
rect 257514 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 258134 295174
rect 257514 294854 258134 294938
rect 257514 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 258134 294854
rect 256739 275636 256805 275637
rect 256739 275572 256740 275636
rect 256804 275572 256805 275636
rect 256739 275571 256805 275572
rect 254531 261084 254597 261085
rect 254531 261020 254532 261084
rect 254596 261020 254597 261084
rect 254531 261019 254597 261020
rect 252875 248164 252941 248165
rect 252875 248100 252876 248164
rect 252940 248100 252941 248164
rect 252875 248099 252941 248100
rect 252878 238770 252938 248099
rect 252510 238710 252938 238770
rect 252510 229110 252570 238710
rect 252510 229050 253122 229110
rect 253062 224773 253122 229050
rect 253059 224772 253125 224773
rect 253059 224708 253060 224772
rect 253124 224708 253125 224772
rect 253059 224707 253125 224708
rect 253062 219197 253122 224707
rect 253794 219454 254414 239592
rect 254534 238645 254594 261019
rect 255267 260676 255333 260677
rect 255267 260612 255268 260676
rect 255332 260612 255333 260676
rect 255267 260611 255333 260612
rect 254531 238644 254597 238645
rect 254531 238580 254532 238644
rect 254596 238580 254597 238644
rect 254531 238579 254597 238580
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253059 219196 253125 219197
rect 253059 219132 253060 219196
rect 253124 219132 253125 219196
rect 253059 219131 253125 219132
rect 253794 219134 254414 219218
rect 253062 206277 253122 219131
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253059 206276 253125 206277
rect 253059 206212 253060 206276
rect 253124 206212 253125 206276
rect 253059 206211 253125 206212
rect 253794 183454 254414 218898
rect 254534 211989 254594 238579
rect 255270 214573 255330 260611
rect 257514 259174 258134 294618
rect 257514 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 258134 259174
rect 257514 258854 258134 258938
rect 257514 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 258134 258854
rect 257514 223174 258134 258618
rect 257514 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 258134 223174
rect 257514 222854 258134 222938
rect 257514 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 258134 222854
rect 255267 214572 255333 214573
rect 255267 214508 255268 214572
rect 255332 214508 255333 214572
rect 255267 214507 255333 214508
rect 254531 211988 254597 211989
rect 254531 211924 254532 211988
rect 254596 211924 254597 211988
rect 254531 211923 254597 211924
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 247723 66196 247789 66197
rect 247723 66132 247724 66196
rect 247788 66132 247789 66196
rect 247723 66131 247789 66132
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 187174 258134 222618
rect 258214 300870 258458 300930
rect 258214 209790 258274 300870
rect 258766 292590 258826 306330
rect 258398 292530 258826 292590
rect 258398 270605 258458 292530
rect 258395 270604 258461 270605
rect 258395 270540 258396 270604
rect 258460 270540 258461 270604
rect 258395 270539 258461 270540
rect 259502 269381 259562 313923
rect 260054 273189 260114 316507
rect 260974 276861 261034 331739
rect 261234 298894 261854 334338
rect 261234 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 261854 298894
rect 261234 298574 261854 298658
rect 261234 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 261854 298574
rect 260971 276860 261037 276861
rect 260971 276796 260972 276860
rect 261036 276796 261037 276860
rect 260971 276795 261037 276796
rect 260051 273188 260117 273189
rect 260051 273124 260052 273188
rect 260116 273124 260117 273188
rect 260051 273123 260117 273124
rect 259499 269380 259565 269381
rect 259499 269316 259500 269380
rect 259564 269316 259565 269380
rect 259499 269315 259565 269316
rect 261234 262894 261854 298338
rect 261234 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 261854 262894
rect 261234 262574 261854 262658
rect 261234 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 261854 262574
rect 259499 259860 259565 259861
rect 259499 259796 259500 259860
rect 259564 259796 259565 259860
rect 259499 259795 259565 259796
rect 258395 253740 258461 253741
rect 258395 253676 258396 253740
rect 258460 253676 258461 253740
rect 258395 253675 258461 253676
rect 258398 236741 258458 253675
rect 258395 236740 258461 236741
rect 258395 236676 258396 236740
rect 258460 236676 258461 236740
rect 258395 236675 258461 236676
rect 259502 231845 259562 259795
rect 259683 242316 259749 242317
rect 259683 242252 259684 242316
rect 259748 242252 259749 242316
rect 259683 242251 259749 242252
rect 259499 231844 259565 231845
rect 259499 231780 259500 231844
rect 259564 231780 259565 231844
rect 259499 231779 259565 231780
rect 259686 223005 259746 242251
rect 261234 226894 261854 262338
rect 262262 259453 262322 424219
rect 264954 410614 265574 446058
rect 264954 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 265574 410614
rect 264954 410294 265574 410378
rect 264954 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 265574 410294
rect 263547 386340 263613 386341
rect 263547 386276 263548 386340
rect 263612 386276 263613 386340
rect 263547 386275 263613 386276
rect 262443 332620 262509 332621
rect 262443 332556 262444 332620
rect 262508 332556 262509 332620
rect 262443 332555 262509 332556
rect 262446 290733 262506 332555
rect 263550 302250 263610 386275
rect 264954 374614 265574 410058
rect 266307 387700 266373 387701
rect 266307 387636 266308 387700
rect 266372 387636 266373 387700
rect 266307 387635 266373 387636
rect 264954 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 265574 374614
rect 264954 374294 265574 374378
rect 264954 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 265574 374294
rect 264954 338614 265574 374058
rect 264954 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 265574 338614
rect 264954 338294 265574 338378
rect 264954 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 265574 338294
rect 263731 316708 263797 316709
rect 263731 316644 263732 316708
rect 263796 316644 263797 316708
rect 263731 316643 263797 316644
rect 263366 302190 263610 302250
rect 263366 292590 263426 302190
rect 263366 292530 263610 292590
rect 262443 290732 262509 290733
rect 262443 290668 262444 290732
rect 262508 290668 262509 290732
rect 262443 290667 262509 290668
rect 262443 263668 262509 263669
rect 262443 263604 262444 263668
rect 262508 263604 262509 263668
rect 262443 263603 262509 263604
rect 262259 259452 262325 259453
rect 262259 259388 262260 259452
rect 262324 259388 262325 259452
rect 262259 259387 262325 259388
rect 262075 249796 262141 249797
rect 262075 249732 262076 249796
rect 262140 249732 262141 249796
rect 262075 249731 262141 249732
rect 262078 240821 262138 249731
rect 262075 240820 262141 240821
rect 262075 240756 262076 240820
rect 262140 240756 262141 240820
rect 262075 240755 262141 240756
rect 262262 228445 262322 259387
rect 262446 249797 262506 263603
rect 263550 261765 263610 292530
rect 263547 261764 263613 261765
rect 263547 261700 263548 261764
rect 263612 261700 263613 261764
rect 263547 261699 263613 261700
rect 262443 249796 262509 249797
rect 262443 249732 262444 249796
rect 262508 249732 262509 249796
rect 262443 249731 262509 249732
rect 262811 247892 262877 247893
rect 262811 247828 262812 247892
rect 262876 247828 262877 247892
rect 262811 247827 262877 247828
rect 262259 228444 262325 228445
rect 262259 228380 262260 228444
rect 262324 228380 262325 228444
rect 262259 228379 262325 228380
rect 261234 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 261854 226894
rect 261234 226574 261854 226658
rect 261234 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 261854 226574
rect 259683 223004 259749 223005
rect 259683 222940 259684 223004
rect 259748 222940 259749 223004
rect 259683 222939 259749 222940
rect 258214 209730 258458 209790
rect 257514 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 258134 187174
rect 257514 186854 258134 186938
rect 257514 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 258134 186854
rect 257514 151174 258134 186618
rect 258398 184245 258458 209730
rect 261234 190894 261854 226338
rect 262814 222869 262874 247827
rect 263550 235789 263610 261699
rect 263734 261357 263794 316643
rect 264954 302614 265574 338058
rect 264954 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 265574 302614
rect 264954 302294 265574 302378
rect 264954 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 265574 302294
rect 264954 266614 265574 302058
rect 265755 298756 265821 298757
rect 265755 298692 265756 298756
rect 265820 298692 265821 298756
rect 265755 298691 265821 298692
rect 264954 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 265574 266614
rect 264954 266294 265574 266378
rect 264954 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 265574 266294
rect 263731 261356 263797 261357
rect 263731 261292 263732 261356
rect 263796 261292 263797 261356
rect 263731 261291 263797 261292
rect 263731 259588 263797 259589
rect 263731 259524 263732 259588
rect 263796 259524 263797 259588
rect 263731 259523 263797 259524
rect 263734 240141 263794 259523
rect 263731 240140 263797 240141
rect 263731 240076 263732 240140
rect 263796 240076 263797 240140
rect 263731 240075 263797 240076
rect 263547 235788 263613 235789
rect 263547 235724 263548 235788
rect 263612 235724 263613 235788
rect 263547 235723 263613 235724
rect 264954 230614 265574 266058
rect 265758 237965 265818 298691
rect 266310 247893 266370 387635
rect 266494 339557 266554 454139
rect 266491 339556 266557 339557
rect 266491 339492 266492 339556
rect 266556 339492 266557 339556
rect 266491 339491 266557 339492
rect 266494 335370 266554 339491
rect 266494 335310 266922 335370
rect 266862 267069 266922 335310
rect 267782 298077 267842 455635
rect 267963 358052 268029 358053
rect 267963 357988 267964 358052
rect 268028 357988 268029 358052
rect 267963 357987 268029 357988
rect 267779 298076 267845 298077
rect 267779 298012 267780 298076
rect 267844 298012 267845 298076
rect 267779 298011 267845 298012
rect 266859 267068 266925 267069
rect 266859 267004 266860 267068
rect 266924 267004 266925 267068
rect 266859 267003 266925 267004
rect 266491 262716 266557 262717
rect 266491 262652 266492 262716
rect 266556 262652 266557 262716
rect 266491 262651 266557 262652
rect 266307 247892 266373 247893
rect 266307 247828 266308 247892
rect 266372 247828 266373 247892
rect 266307 247827 266373 247828
rect 265755 237964 265821 237965
rect 265755 237900 265756 237964
rect 265820 237900 265821 237964
rect 265755 237899 265821 237900
rect 264954 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 265574 230614
rect 264954 230294 265574 230378
rect 264954 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 265574 230294
rect 262811 222868 262877 222869
rect 262811 222804 262812 222868
rect 262876 222804 262877 222868
rect 262811 222803 262877 222804
rect 261234 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 261854 190894
rect 261234 190574 261854 190658
rect 261234 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 261854 190574
rect 258395 184244 258461 184245
rect 258395 184180 258396 184244
rect 258460 184180 258461 184244
rect 258395 184179 258461 184180
rect 257514 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 258134 151174
rect 257514 150854 258134 150938
rect 257514 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 258134 150854
rect 257514 115174 258134 150618
rect 257514 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 258134 115174
rect 257514 114854 258134 114938
rect 257514 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 258134 114854
rect 257514 79174 258134 114618
rect 257514 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 258134 79174
rect 257514 78854 258134 78938
rect 257514 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 258134 78854
rect 257514 43174 258134 78618
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 154894 261854 190338
rect 261234 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 261854 154894
rect 261234 154574 261854 154658
rect 261234 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 261854 154574
rect 261234 118894 261854 154338
rect 261234 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 261854 118894
rect 261234 118574 261854 118658
rect 261234 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 261854 118574
rect 261234 82894 261854 118338
rect 261234 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 261854 82894
rect 261234 82574 261854 82658
rect 261234 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 261854 82574
rect 261234 46894 261854 82338
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 194614 265574 230058
rect 266494 228309 266554 262651
rect 267966 256869 268026 357987
rect 268331 295356 268397 295357
rect 268331 295292 268332 295356
rect 268396 295292 268397 295356
rect 268331 295291 268397 295292
rect 268334 280941 268394 295291
rect 268331 280940 268397 280941
rect 268331 280876 268332 280940
rect 268396 280876 268397 280940
rect 268331 280875 268397 280876
rect 269070 264893 269130 465155
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 270539 403612 270605 403613
rect 270539 403548 270540 403612
rect 270604 403548 270605 403612
rect 270539 403547 270605 403548
rect 269251 363084 269317 363085
rect 269251 363020 269252 363084
rect 269316 363020 269317 363084
rect 269251 363019 269317 363020
rect 269067 264892 269133 264893
rect 269067 264828 269068 264892
rect 269132 264828 269133 264892
rect 269067 264827 269133 264828
rect 267963 256868 268029 256869
rect 267963 256804 267964 256868
rect 268028 256804 268029 256868
rect 267963 256803 268029 256804
rect 269254 255237 269314 363019
rect 270542 258909 270602 403547
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 270723 318068 270789 318069
rect 270723 318004 270724 318068
rect 270788 318004 270789 318068
rect 270723 318003 270789 318004
rect 270726 263669 270786 318003
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 601174 276134 636618
rect 275514 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 276134 601174
rect 275514 600854 276134 600938
rect 275514 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 276134 600854
rect 275514 565174 276134 600618
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 529174 276134 564618
rect 275514 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 276134 529174
rect 275514 528854 276134 528938
rect 275514 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 276134 528854
rect 275514 493174 276134 528618
rect 275514 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 276134 493174
rect 275514 492854 276134 492938
rect 275514 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 276134 492854
rect 275514 457174 276134 492618
rect 275514 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 276134 457174
rect 275514 456854 276134 456938
rect 275514 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 276134 456854
rect 275514 421174 276134 456618
rect 275514 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 276134 421174
rect 275514 420854 276134 420938
rect 275514 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 276134 420854
rect 275514 385174 276134 420618
rect 275514 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 276134 385174
rect 275514 384854 276134 384938
rect 275514 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 276134 384854
rect 275514 349174 276134 384618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 604894 279854 640338
rect 279234 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 279854 604894
rect 279234 604574 279854 604658
rect 279234 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 279854 604574
rect 279234 568894 279854 604338
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 279234 532894 279854 568338
rect 279234 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 279854 532894
rect 279234 532574 279854 532658
rect 279234 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 279854 532574
rect 279234 496894 279854 532338
rect 279234 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 279854 496894
rect 279234 496574 279854 496658
rect 279234 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 279854 496574
rect 279234 460894 279854 496338
rect 279234 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 279854 460894
rect 279234 460574 279854 460658
rect 279234 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 279854 460574
rect 279234 424894 279854 460338
rect 279234 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 279854 424894
rect 279234 424574 279854 424658
rect 279234 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 279854 424574
rect 279234 388894 279854 424338
rect 279234 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 279854 388894
rect 279234 388574 279854 388658
rect 279234 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 279854 388574
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 608614 283574 644058
rect 282954 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 283574 608614
rect 282954 608294 283574 608378
rect 282954 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 283574 608294
rect 282954 572614 283574 608058
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 536614 283574 572058
rect 282954 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 283574 536614
rect 282954 536294 283574 536378
rect 282954 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 283574 536294
rect 282954 500614 283574 536058
rect 282954 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 283574 500614
rect 282954 500294 283574 500378
rect 282954 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 283574 500294
rect 282954 464614 283574 500058
rect 282954 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 283574 464614
rect 282954 464294 283574 464378
rect 282954 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 283574 464294
rect 282954 428614 283574 464058
rect 282954 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 283574 428614
rect 282954 428294 283574 428378
rect 282954 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 283574 428294
rect 282954 392614 283574 428058
rect 282954 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 283574 392614
rect 282954 392294 283574 392378
rect 282954 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 283574 392294
rect 276243 379540 276309 379541
rect 276243 379476 276244 379540
rect 276308 379476 276309 379540
rect 276243 379475 276309 379476
rect 275514 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 276134 349174
rect 275514 348854 276134 348938
rect 275514 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 276134 348854
rect 275514 313174 276134 348618
rect 275514 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 276134 313174
rect 275514 312854 276134 312938
rect 275514 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 276134 312854
rect 273299 305828 273365 305829
rect 273299 305764 273300 305828
rect 273364 305764 273365 305828
rect 273299 305763 273365 305764
rect 272563 299436 272629 299437
rect 272563 299372 272564 299436
rect 272628 299372 272629 299436
rect 272563 299371 272629 299372
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 270723 263668 270789 263669
rect 270723 263604 270724 263668
rect 270788 263604 270789 263668
rect 270723 263603 270789 263604
rect 270723 259588 270789 259589
rect 270723 259524 270724 259588
rect 270788 259524 270789 259588
rect 270723 259523 270789 259524
rect 270539 258908 270605 258909
rect 270539 258844 270540 258908
rect 270604 258844 270605 258908
rect 270539 258843 270605 258844
rect 269251 255236 269317 255237
rect 269251 255172 269252 255236
rect 269316 255172 269317 255236
rect 269251 255171 269317 255172
rect 269067 252652 269133 252653
rect 269067 252588 269068 252652
rect 269132 252588 269133 252652
rect 269067 252587 269133 252588
rect 267779 248436 267845 248437
rect 267779 248372 267780 248436
rect 267844 248372 267845 248436
rect 267779 248371 267845 248372
rect 266491 228308 266557 228309
rect 266491 228244 266492 228308
rect 266556 228244 266557 228308
rect 266491 228243 266557 228244
rect 267782 217973 267842 248371
rect 267779 217972 267845 217973
rect 267779 217908 267780 217972
rect 267844 217908 267845 217972
rect 267779 217907 267845 217908
rect 264954 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 265574 194614
rect 264954 194294 265574 194378
rect 264954 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 265574 194294
rect 264954 158614 265574 194058
rect 269070 181389 269130 252587
rect 270726 219333 270786 259523
rect 271794 237454 272414 272898
rect 272566 251157 272626 299371
rect 272563 251156 272629 251157
rect 272563 251092 272564 251156
rect 272628 251092 272629 251156
rect 272563 251091 272629 251092
rect 273302 242861 273362 305763
rect 274587 303788 274653 303789
rect 274587 303724 274588 303788
rect 274652 303724 274653 303788
rect 274587 303723 274653 303724
rect 273299 242860 273365 242861
rect 273299 242796 273300 242860
rect 273364 242796 273365 242860
rect 273299 242795 273365 242796
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 270723 219332 270789 219333
rect 270723 219268 270724 219332
rect 270788 219268 270789 219332
rect 270723 219267 270789 219268
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 269067 181388 269133 181389
rect 269067 181324 269068 181388
rect 269132 181324 269133 181388
rect 269067 181323 269133 181324
rect 264954 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 265574 158614
rect 264954 158294 265574 158378
rect 264954 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 265574 158294
rect 264954 122614 265574 158058
rect 264954 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 265574 122614
rect 264954 122294 265574 122378
rect 264954 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 265574 122294
rect 264954 86614 265574 122058
rect 264954 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 265574 86614
rect 264954 86294 265574 86378
rect 264954 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 265574 86294
rect 264954 50614 265574 86058
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 274590 71773 274650 303723
rect 275514 277174 276134 312618
rect 275514 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 276134 277174
rect 275514 276854 276134 276938
rect 275514 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 276134 276854
rect 275514 241174 276134 276618
rect 276246 266797 276306 379475
rect 279234 352894 279854 388338
rect 281579 388380 281645 388381
rect 281579 388316 281580 388380
rect 281644 388316 281645 388380
rect 281579 388315 281645 388316
rect 279234 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 279854 352894
rect 279234 352574 279854 352658
rect 279234 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 279854 352574
rect 279234 316894 279854 352338
rect 279234 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 279854 316894
rect 279234 316574 279854 316658
rect 279234 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 279854 316574
rect 277163 313988 277229 313989
rect 277163 313924 277164 313988
rect 277228 313924 277229 313988
rect 277163 313923 277229 313924
rect 276243 266796 276309 266797
rect 276243 266732 276244 266796
rect 276308 266732 276309 266796
rect 276243 266731 276309 266732
rect 276243 263668 276309 263669
rect 276243 263604 276244 263668
rect 276308 263604 276309 263668
rect 276243 263603 276309 263604
rect 275514 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 276134 241174
rect 275514 240854 276134 240938
rect 275514 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 276134 240854
rect 275514 205174 276134 240618
rect 276246 214573 276306 263603
rect 277166 242317 277226 313923
rect 279234 280894 279854 316338
rect 279234 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 279854 280894
rect 279234 280574 279854 280658
rect 279234 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 279854 280574
rect 279234 244894 279854 280338
rect 281582 264213 281642 388315
rect 282954 356614 283574 392058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 285627 386340 285693 386341
rect 285627 386276 285628 386340
rect 285692 386276 285693 386340
rect 285627 386275 285693 386276
rect 285630 385661 285690 386275
rect 285627 385660 285693 385661
rect 285627 385596 285628 385660
rect 285692 385596 285693 385660
rect 285627 385595 285693 385596
rect 282954 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 283574 356614
rect 282954 356294 283574 356378
rect 282954 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 283574 356294
rect 282954 320614 283574 356058
rect 282954 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 283574 320614
rect 282954 320294 283574 320378
rect 282954 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 283574 320294
rect 282954 284614 283574 320058
rect 282954 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 283574 284614
rect 282954 284294 283574 284378
rect 282954 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 283574 284294
rect 281579 264212 281645 264213
rect 281579 264148 281580 264212
rect 281644 264148 281645 264212
rect 281579 264147 281645 264148
rect 279234 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 279854 244894
rect 279234 244574 279854 244658
rect 279234 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 279854 244574
rect 277163 242316 277229 242317
rect 277163 242252 277164 242316
rect 277228 242252 277229 242316
rect 277163 242251 277229 242252
rect 276243 214572 276309 214573
rect 276243 214508 276244 214572
rect 276308 214508 276309 214572
rect 276243 214507 276309 214508
rect 275514 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 276134 205174
rect 275514 204854 276134 204938
rect 275514 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 276134 204854
rect 275514 169174 276134 204618
rect 275514 168938 275546 169174
rect 275782 168938 275866 169174
rect 276102 168938 276134 169174
rect 275514 168854 276134 168938
rect 275514 168618 275546 168854
rect 275782 168618 275866 168854
rect 276102 168618 276134 168854
rect 275514 133174 276134 168618
rect 275514 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 276134 133174
rect 275514 132854 276134 132938
rect 275514 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 276134 132854
rect 275514 97174 276134 132618
rect 275514 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 276134 97174
rect 275514 96854 276134 96938
rect 275514 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 276134 96854
rect 274587 71772 274653 71773
rect 274587 71708 274588 71772
rect 274652 71708 274653 71772
rect 274587 71707 274653 71708
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 61174 276134 96618
rect 275514 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 276134 61174
rect 275514 60854 276134 60938
rect 275514 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 276134 60854
rect 275514 25174 276134 60618
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 208894 279854 244338
rect 279234 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 279854 208894
rect 279234 208574 279854 208658
rect 279234 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 279854 208574
rect 279234 172894 279854 208338
rect 279234 172658 279266 172894
rect 279502 172658 279586 172894
rect 279822 172658 279854 172894
rect 279234 172574 279854 172658
rect 279234 172338 279266 172574
rect 279502 172338 279586 172574
rect 279822 172338 279854 172574
rect 279234 136894 279854 172338
rect 279234 136658 279266 136894
rect 279502 136658 279586 136894
rect 279822 136658 279854 136894
rect 279234 136574 279854 136658
rect 279234 136338 279266 136574
rect 279502 136338 279586 136574
rect 279822 136338 279854 136574
rect 279234 100894 279854 136338
rect 279234 100658 279266 100894
rect 279502 100658 279586 100894
rect 279822 100658 279854 100894
rect 279234 100574 279854 100658
rect 279234 100338 279266 100574
rect 279502 100338 279586 100574
rect 279822 100338 279854 100574
rect 279234 64894 279854 100338
rect 279234 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 279854 64894
rect 279234 64574 279854 64658
rect 279234 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 279854 64574
rect 279234 28894 279854 64338
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 248614 283574 284058
rect 285630 254557 285690 385595
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 285627 254556 285693 254557
rect 285627 254492 285628 254556
rect 285692 254492 285693 254556
rect 285627 254491 285693 254492
rect 282954 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 283574 248614
rect 282954 248294 283574 248378
rect 282954 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 283574 248294
rect 282954 212614 283574 248058
rect 282954 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 283574 212614
rect 282954 212294 283574 212378
rect 282954 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 283574 212294
rect 282954 176614 283574 212058
rect 282954 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 283574 176614
rect 282954 176294 283574 176378
rect 282954 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 283574 176294
rect 282954 140614 283574 176058
rect 282954 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 283574 140614
rect 282954 140294 283574 140378
rect 282954 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 283574 140294
rect 282954 104614 283574 140058
rect 282954 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 283574 104614
rect 282954 104294 283574 104378
rect 282954 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 283574 104294
rect 282954 68614 283574 104058
rect 282954 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 283574 68614
rect 282954 68294 283574 68378
rect 282954 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 283574 68294
rect 282954 32614 283574 68058
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 511174 294134 546618
rect 293514 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 294134 511174
rect 293514 510854 294134 510938
rect 293514 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 294134 510854
rect 293514 475174 294134 510618
rect 293514 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 294134 475174
rect 293514 474854 294134 474938
rect 293514 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 294134 474854
rect 293514 439174 294134 474618
rect 293514 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 294134 439174
rect 293514 438854 294134 438938
rect 293514 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 294134 438854
rect 293514 403174 294134 438618
rect 293514 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 294134 403174
rect 293514 402854 294134 402938
rect 293514 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 294134 402854
rect 293514 367174 294134 402618
rect 293514 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 294134 367174
rect 293514 366854 294134 366938
rect 293514 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 294134 366854
rect 293514 331174 294134 366618
rect 293514 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 294134 331174
rect 293514 330854 294134 330938
rect 293514 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 294134 330854
rect 293514 295174 294134 330618
rect 293514 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 294134 295174
rect 293514 294854 294134 294938
rect 293514 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 294134 294854
rect 293514 259174 294134 294618
rect 293514 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 294134 259174
rect 293514 258854 294134 258938
rect 293514 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 294134 258854
rect 293514 223174 294134 258618
rect 293514 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 294134 223174
rect 293514 222854 294134 222938
rect 293514 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 294134 222854
rect 293514 187174 294134 222618
rect 293514 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 294134 187174
rect 293514 186854 294134 186938
rect 293514 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 294134 186854
rect 293514 151174 294134 186618
rect 293514 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 294134 151174
rect 293514 150854 294134 150938
rect 293514 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 294134 150854
rect 293514 115174 294134 150618
rect 293514 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 294134 115174
rect 293514 114854 294134 114938
rect 293514 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 294134 114854
rect 293514 79174 294134 114618
rect 293514 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 294134 79174
rect 293514 78854 294134 78938
rect 293514 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 294134 78854
rect 293514 43174 294134 78618
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 514894 297854 550338
rect 297234 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 297854 514894
rect 297234 514574 297854 514658
rect 297234 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 297854 514574
rect 297234 478894 297854 514338
rect 297234 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 297854 478894
rect 297234 478574 297854 478658
rect 297234 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 297854 478574
rect 297234 442894 297854 478338
rect 297234 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 297854 442894
rect 297234 442574 297854 442658
rect 297234 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 297854 442574
rect 297234 406894 297854 442338
rect 297234 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 297854 406894
rect 297234 406574 297854 406658
rect 297234 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 297854 406574
rect 297234 370894 297854 406338
rect 297234 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 297854 370894
rect 297234 370574 297854 370658
rect 297234 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 297854 370574
rect 297234 334894 297854 370338
rect 297234 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 297854 334894
rect 297234 334574 297854 334658
rect 297234 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 297854 334574
rect 297234 298894 297854 334338
rect 297234 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 297854 298894
rect 297234 298574 297854 298658
rect 297234 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 297854 298574
rect 297234 262894 297854 298338
rect 297234 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 297854 262894
rect 297234 262574 297854 262658
rect 297234 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 297854 262574
rect 297234 226894 297854 262338
rect 297234 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 297854 226894
rect 297234 226574 297854 226658
rect 297234 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 297854 226574
rect 297234 190894 297854 226338
rect 297234 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 297854 190894
rect 297234 190574 297854 190658
rect 297234 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 297854 190574
rect 297234 154894 297854 190338
rect 297234 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 297854 154894
rect 297234 154574 297854 154658
rect 297234 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 297854 154574
rect 297234 118894 297854 154338
rect 297234 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 297854 118894
rect 297234 118574 297854 118658
rect 297234 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 297854 118574
rect 297234 82894 297854 118338
rect 297234 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 297854 82894
rect 297234 82574 297854 82658
rect 297234 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 297854 82574
rect 297234 46894 297854 82338
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 518614 301574 554058
rect 300954 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 301574 518614
rect 300954 518294 301574 518378
rect 300954 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 301574 518294
rect 300954 482614 301574 518058
rect 300954 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 301574 482614
rect 300954 482294 301574 482378
rect 300954 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 301574 482294
rect 300954 446614 301574 482058
rect 300954 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 301574 446614
rect 300954 446294 301574 446378
rect 300954 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 301574 446294
rect 300954 410614 301574 446058
rect 300954 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 301574 410614
rect 300954 410294 301574 410378
rect 300954 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 301574 410294
rect 300954 374614 301574 410058
rect 300954 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 301574 374614
rect 300954 374294 301574 374378
rect 300954 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 301574 374294
rect 300954 338614 301574 374058
rect 300954 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 301574 338614
rect 300954 338294 301574 338378
rect 300954 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 301574 338294
rect 300954 302614 301574 338058
rect 300954 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 301574 302614
rect 300954 302294 301574 302378
rect 300954 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 301574 302294
rect 300954 266614 301574 302058
rect 300954 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 301574 266614
rect 300954 266294 301574 266378
rect 300954 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 301574 266294
rect 300954 230614 301574 266058
rect 300954 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 301574 230614
rect 300954 230294 301574 230378
rect 300954 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 301574 230294
rect 300954 194614 301574 230058
rect 300954 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 301574 194614
rect 300954 194294 301574 194378
rect 300954 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 301574 194294
rect 300954 158614 301574 194058
rect 300954 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 301574 158614
rect 300954 158294 301574 158378
rect 300954 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 301574 158294
rect 300954 122614 301574 158058
rect 300954 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 301574 122614
rect 300954 122294 301574 122378
rect 300954 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 301574 122294
rect 300954 86614 301574 122058
rect 300954 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 301574 86614
rect 300954 86294 301574 86378
rect 300954 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 301574 86294
rect 300954 50614 301574 86058
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 529174 312134 564618
rect 311514 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 312134 529174
rect 311514 528854 312134 528938
rect 311514 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 312134 528854
rect 311514 493174 312134 528618
rect 311514 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 312134 493174
rect 311514 492854 312134 492938
rect 311514 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 312134 492854
rect 311514 457174 312134 492618
rect 311514 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 312134 457174
rect 311514 456854 312134 456938
rect 311514 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 312134 456854
rect 311514 421174 312134 456618
rect 311514 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 312134 421174
rect 311514 420854 312134 420938
rect 311514 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 312134 420854
rect 311514 385174 312134 420618
rect 311514 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 312134 385174
rect 311514 384854 312134 384938
rect 311514 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 312134 384854
rect 311514 349174 312134 384618
rect 311514 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 312134 349174
rect 311514 348854 312134 348938
rect 311514 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 312134 348854
rect 311514 313174 312134 348618
rect 311514 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 312134 313174
rect 311514 312854 312134 312938
rect 311514 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 312134 312854
rect 311514 277174 312134 312618
rect 311514 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 312134 277174
rect 311514 276854 312134 276938
rect 311514 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 312134 276854
rect 311514 241174 312134 276618
rect 311514 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 312134 241174
rect 311514 240854 312134 240938
rect 311514 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 312134 240854
rect 311514 205174 312134 240618
rect 311514 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 312134 205174
rect 311514 204854 312134 204938
rect 311514 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 312134 204854
rect 311514 169174 312134 204618
rect 311514 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 312134 169174
rect 311514 168854 312134 168938
rect 311514 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 312134 168854
rect 311514 133174 312134 168618
rect 311514 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 312134 133174
rect 311514 132854 312134 132938
rect 311514 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 312134 132854
rect 311514 97174 312134 132618
rect 311514 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 312134 97174
rect 311514 96854 312134 96938
rect 311514 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 312134 96854
rect 311514 61174 312134 96618
rect 311514 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 312134 61174
rect 311514 60854 312134 60938
rect 311514 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 312134 60854
rect 311514 25174 312134 60618
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 532894 315854 568338
rect 315234 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 315854 532894
rect 315234 532574 315854 532658
rect 315234 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 315854 532574
rect 315234 496894 315854 532338
rect 315234 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 315854 496894
rect 315234 496574 315854 496658
rect 315234 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 315854 496574
rect 315234 460894 315854 496338
rect 315234 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 315854 460894
rect 315234 460574 315854 460658
rect 315234 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 315854 460574
rect 315234 424894 315854 460338
rect 315234 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 315854 424894
rect 315234 424574 315854 424658
rect 315234 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 315854 424574
rect 315234 388894 315854 424338
rect 315234 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 315854 388894
rect 315234 388574 315854 388658
rect 315234 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 315854 388574
rect 315234 352894 315854 388338
rect 315234 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 315854 352894
rect 315234 352574 315854 352658
rect 315234 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 315854 352574
rect 315234 316894 315854 352338
rect 315234 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 315854 316894
rect 315234 316574 315854 316658
rect 315234 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 315854 316574
rect 315234 280894 315854 316338
rect 315234 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 315854 280894
rect 315234 280574 315854 280658
rect 315234 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 315854 280574
rect 315234 244894 315854 280338
rect 315234 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 315854 244894
rect 315234 244574 315854 244658
rect 315234 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 315854 244574
rect 315234 208894 315854 244338
rect 315234 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 315854 208894
rect 315234 208574 315854 208658
rect 315234 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 315854 208574
rect 315234 172894 315854 208338
rect 315234 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 315854 172894
rect 315234 172574 315854 172658
rect 315234 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 315854 172574
rect 315234 136894 315854 172338
rect 315234 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 315854 136894
rect 315234 136574 315854 136658
rect 315234 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 315854 136574
rect 315234 100894 315854 136338
rect 315234 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 315854 100894
rect 315234 100574 315854 100658
rect 315234 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 315854 100574
rect 315234 64894 315854 100338
rect 315234 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 315854 64894
rect 315234 64574 315854 64658
rect 315234 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 315854 64574
rect 315234 28894 315854 64338
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 536614 319574 572058
rect 318954 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 319574 536614
rect 318954 536294 319574 536378
rect 318954 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 319574 536294
rect 318954 500614 319574 536058
rect 318954 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 319574 500614
rect 318954 500294 319574 500378
rect 318954 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 319574 500294
rect 318954 464614 319574 500058
rect 318954 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 319574 464614
rect 318954 464294 319574 464378
rect 318954 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 319574 464294
rect 318954 428614 319574 464058
rect 318954 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 319574 428614
rect 318954 428294 319574 428378
rect 318954 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 319574 428294
rect 318954 392614 319574 428058
rect 318954 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 319574 392614
rect 318954 392294 319574 392378
rect 318954 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 319574 392294
rect 318954 356614 319574 392058
rect 318954 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 319574 356614
rect 318954 356294 319574 356378
rect 318954 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 319574 356294
rect 318954 320614 319574 356058
rect 318954 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 319574 320614
rect 318954 320294 319574 320378
rect 318954 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 319574 320294
rect 318954 284614 319574 320058
rect 318954 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 319574 284614
rect 318954 284294 319574 284378
rect 318954 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 319574 284294
rect 318954 248614 319574 284058
rect 318954 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 319574 248614
rect 318954 248294 319574 248378
rect 318954 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 319574 248294
rect 318954 212614 319574 248058
rect 318954 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 319574 212614
rect 318954 212294 319574 212378
rect 318954 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 319574 212294
rect 318954 176614 319574 212058
rect 318954 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 319574 176614
rect 318954 176294 319574 176378
rect 318954 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 319574 176294
rect 318954 140614 319574 176058
rect 318954 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 319574 140614
rect 318954 140294 319574 140378
rect 318954 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 319574 140294
rect 318954 104614 319574 140058
rect 318954 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 319574 104614
rect 318954 104294 319574 104378
rect 318954 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 319574 104294
rect 318954 68614 319574 104058
rect 318954 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 319574 68614
rect 318954 68294 319574 68378
rect 318954 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 319574 68294
rect 318954 32614 319574 68058
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547174 330134 582618
rect 329514 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 330134 547174
rect 329514 546854 330134 546938
rect 329514 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 330134 546854
rect 329514 511174 330134 546618
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 475174 330134 510618
rect 329514 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 330134 475174
rect 329514 474854 330134 474938
rect 329514 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 330134 474854
rect 329514 439174 330134 474618
rect 329514 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 330134 439174
rect 329514 438854 330134 438938
rect 329514 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 330134 438854
rect 329514 403174 330134 438618
rect 329514 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 330134 403174
rect 329514 402854 330134 402938
rect 329514 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 330134 402854
rect 329514 367174 330134 402618
rect 329514 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 330134 367174
rect 329514 366854 330134 366938
rect 329514 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 330134 366854
rect 329514 331174 330134 366618
rect 329514 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 330134 331174
rect 329514 330854 330134 330938
rect 329514 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 330134 330854
rect 329514 295174 330134 330618
rect 329514 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 330134 295174
rect 329514 294854 330134 294938
rect 329514 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 330134 294854
rect 329514 259174 330134 294618
rect 329514 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 330134 259174
rect 329514 258854 330134 258938
rect 329514 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 330134 258854
rect 329514 223174 330134 258618
rect 329514 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 330134 223174
rect 329514 222854 330134 222938
rect 329514 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 330134 222854
rect 329514 187174 330134 222618
rect 329514 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 330134 187174
rect 329514 186854 330134 186938
rect 329514 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 330134 186854
rect 329514 151174 330134 186618
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 115174 330134 150618
rect 329514 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 330134 115174
rect 329514 114854 330134 114938
rect 329514 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 330134 114854
rect 329514 79174 330134 114618
rect 329514 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 330134 79174
rect 329514 78854 330134 78938
rect 329514 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 330134 78854
rect 329514 43174 330134 78618
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 550894 333854 586338
rect 333234 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 333854 550894
rect 333234 550574 333854 550658
rect 333234 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 333854 550574
rect 333234 514894 333854 550338
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 478894 333854 514338
rect 333234 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 333854 478894
rect 333234 478574 333854 478658
rect 333234 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 333854 478574
rect 333234 442894 333854 478338
rect 333234 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 333854 442894
rect 333234 442574 333854 442658
rect 333234 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 333854 442574
rect 333234 406894 333854 442338
rect 333234 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 333854 406894
rect 333234 406574 333854 406658
rect 333234 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 333854 406574
rect 333234 370894 333854 406338
rect 333234 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 333854 370894
rect 333234 370574 333854 370658
rect 333234 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 333854 370574
rect 333234 334894 333854 370338
rect 333234 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 333854 334894
rect 333234 334574 333854 334658
rect 333234 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 333854 334574
rect 333234 298894 333854 334338
rect 333234 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 333854 298894
rect 333234 298574 333854 298658
rect 333234 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 333854 298574
rect 333234 262894 333854 298338
rect 333234 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 333854 262894
rect 333234 262574 333854 262658
rect 333234 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 333854 262574
rect 333234 226894 333854 262338
rect 333234 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 333854 226894
rect 333234 226574 333854 226658
rect 333234 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 333854 226574
rect 333234 190894 333854 226338
rect 333234 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 333854 190894
rect 333234 190574 333854 190658
rect 333234 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 333854 190574
rect 333234 154894 333854 190338
rect 333234 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 333854 154894
rect 333234 154574 333854 154658
rect 333234 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 333854 154574
rect 333234 118894 333854 154338
rect 333234 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 333854 118894
rect 333234 118574 333854 118658
rect 333234 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 333854 118574
rect 333234 82894 333854 118338
rect 333234 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 333854 82894
rect 333234 82574 333854 82658
rect 333234 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 333854 82574
rect 333234 46894 333854 82338
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 336954 518614 337574 554058
rect 336954 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 337574 518614
rect 336954 518294 337574 518378
rect 336954 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 337574 518294
rect 336954 482614 337574 518058
rect 336954 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 337574 482614
rect 336954 482294 337574 482378
rect 336954 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 337574 482294
rect 336954 446614 337574 482058
rect 336954 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 337574 446614
rect 336954 446294 337574 446378
rect 336954 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 337574 446294
rect 336954 410614 337574 446058
rect 336954 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 337574 410614
rect 336954 410294 337574 410378
rect 336954 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 337574 410294
rect 336954 374614 337574 410058
rect 336954 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 337574 374614
rect 336954 374294 337574 374378
rect 336954 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 337574 374294
rect 336954 338614 337574 374058
rect 336954 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 337574 338614
rect 336954 338294 337574 338378
rect 336954 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 337574 338294
rect 336954 302614 337574 338058
rect 336954 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 337574 302614
rect 336954 302294 337574 302378
rect 336954 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 337574 302294
rect 336954 266614 337574 302058
rect 336954 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 337574 266614
rect 336954 266294 337574 266378
rect 336954 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 337574 266294
rect 336954 230614 337574 266058
rect 336954 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 337574 230614
rect 336954 230294 337574 230378
rect 336954 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 337574 230294
rect 336954 194614 337574 230058
rect 336954 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 337574 194614
rect 336954 194294 337574 194378
rect 336954 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 337574 194294
rect 336954 158614 337574 194058
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 336954 122614 337574 158058
rect 336954 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 337574 122614
rect 336954 122294 337574 122378
rect 336954 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 337574 122294
rect 336954 86614 337574 122058
rect 336954 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 337574 86614
rect 336954 86294 337574 86378
rect 336954 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 337574 86294
rect 336954 50614 337574 86058
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 565174 348134 600618
rect 347514 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 348134 565174
rect 347514 564854 348134 564938
rect 347514 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 348134 564854
rect 347514 529174 348134 564618
rect 347514 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 348134 529174
rect 347514 528854 348134 528938
rect 347514 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 348134 528854
rect 347514 493174 348134 528618
rect 347514 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 348134 493174
rect 347514 492854 348134 492938
rect 347514 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 348134 492854
rect 347514 457174 348134 492618
rect 347514 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 348134 457174
rect 347514 456854 348134 456938
rect 347514 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 348134 456854
rect 347514 421174 348134 456618
rect 347514 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 348134 421174
rect 347514 420854 348134 420938
rect 347514 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 348134 420854
rect 347514 385174 348134 420618
rect 347514 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 348134 385174
rect 347514 384854 348134 384938
rect 347514 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 348134 384854
rect 347514 349174 348134 384618
rect 347514 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 348134 349174
rect 347514 348854 348134 348938
rect 347514 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 348134 348854
rect 347514 313174 348134 348618
rect 347514 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 348134 313174
rect 347514 312854 348134 312938
rect 347514 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 348134 312854
rect 347514 277174 348134 312618
rect 347514 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 348134 277174
rect 347514 276854 348134 276938
rect 347514 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 348134 276854
rect 347514 241174 348134 276618
rect 347514 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 348134 241174
rect 347514 240854 348134 240938
rect 347514 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 348134 240854
rect 347514 205174 348134 240618
rect 347514 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 348134 205174
rect 347514 204854 348134 204938
rect 347514 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 348134 204854
rect 347514 169174 348134 204618
rect 347514 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 348134 169174
rect 347514 168854 348134 168938
rect 347514 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 348134 168854
rect 347514 133174 348134 168618
rect 347514 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 348134 133174
rect 347514 132854 348134 132938
rect 347514 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 348134 132854
rect 347514 97174 348134 132618
rect 347514 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 348134 97174
rect 347514 96854 348134 96938
rect 347514 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 348134 96854
rect 347514 61174 348134 96618
rect 347514 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 348134 61174
rect 347514 60854 348134 60938
rect 347514 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 348134 60854
rect 347514 25174 348134 60618
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 568894 351854 604338
rect 351234 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 351854 568894
rect 351234 568574 351854 568658
rect 351234 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 351854 568574
rect 351234 532894 351854 568338
rect 351234 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 351854 532894
rect 351234 532574 351854 532658
rect 351234 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 351854 532574
rect 351234 496894 351854 532338
rect 351234 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 351854 496894
rect 351234 496574 351854 496658
rect 351234 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 351854 496574
rect 351234 460894 351854 496338
rect 351234 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 351854 460894
rect 351234 460574 351854 460658
rect 351234 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 351854 460574
rect 351234 424894 351854 460338
rect 351234 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 351854 424894
rect 351234 424574 351854 424658
rect 351234 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 351854 424574
rect 351234 388894 351854 424338
rect 351234 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 351854 388894
rect 351234 388574 351854 388658
rect 351234 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 351854 388574
rect 351234 352894 351854 388338
rect 351234 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 351854 352894
rect 351234 352574 351854 352658
rect 351234 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 351854 352574
rect 351234 316894 351854 352338
rect 351234 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 351854 316894
rect 351234 316574 351854 316658
rect 351234 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 351854 316574
rect 351234 280894 351854 316338
rect 351234 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 351854 280894
rect 351234 280574 351854 280658
rect 351234 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 351854 280574
rect 351234 244894 351854 280338
rect 351234 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 351854 244894
rect 351234 244574 351854 244658
rect 351234 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 351854 244574
rect 351234 208894 351854 244338
rect 351234 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 351854 208894
rect 351234 208574 351854 208658
rect 351234 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 351854 208574
rect 351234 172894 351854 208338
rect 351234 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 351854 172894
rect 351234 172574 351854 172658
rect 351234 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 351854 172574
rect 351234 136894 351854 172338
rect 351234 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 351854 136894
rect 351234 136574 351854 136658
rect 351234 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 351854 136574
rect 351234 100894 351854 136338
rect 351234 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 351854 100894
rect 351234 100574 351854 100658
rect 351234 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 351854 100574
rect 351234 64894 351854 100338
rect 351234 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 351854 64894
rect 351234 64574 351854 64658
rect 351234 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 351854 64574
rect 351234 28894 351854 64338
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 354954 536614 355574 572058
rect 354954 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 355574 536614
rect 354954 536294 355574 536378
rect 354954 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 355574 536294
rect 354954 500614 355574 536058
rect 354954 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 355574 500614
rect 354954 500294 355574 500378
rect 354954 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 355574 500294
rect 354954 464614 355574 500058
rect 354954 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 355574 464614
rect 354954 464294 355574 464378
rect 354954 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 355574 464294
rect 354954 428614 355574 464058
rect 354954 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 355574 428614
rect 354954 428294 355574 428378
rect 354954 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 355574 428294
rect 354954 392614 355574 428058
rect 354954 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 355574 392614
rect 354954 392294 355574 392378
rect 354954 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 355574 392294
rect 354954 356614 355574 392058
rect 354954 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 355574 356614
rect 354954 356294 355574 356378
rect 354954 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 355574 356294
rect 354954 320614 355574 356058
rect 354954 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 355574 320614
rect 354954 320294 355574 320378
rect 354954 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 355574 320294
rect 354954 284614 355574 320058
rect 354954 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 355574 284614
rect 354954 284294 355574 284378
rect 354954 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 355574 284294
rect 354954 248614 355574 284058
rect 354954 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 355574 248614
rect 354954 248294 355574 248378
rect 354954 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 355574 248294
rect 354954 212614 355574 248058
rect 354954 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 355574 212614
rect 354954 212294 355574 212378
rect 354954 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 355574 212294
rect 354954 176614 355574 212058
rect 354954 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 355574 176614
rect 354954 176294 355574 176378
rect 354954 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 355574 176294
rect 354954 140614 355574 176058
rect 354954 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 355574 140614
rect 354954 140294 355574 140378
rect 354954 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 355574 140294
rect 354954 104614 355574 140058
rect 354954 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 355574 104614
rect 354954 104294 355574 104378
rect 354954 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 355574 104294
rect 354954 68614 355574 104058
rect 354954 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 355574 68614
rect 354954 68294 355574 68378
rect 354954 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 355574 68294
rect 354954 32614 355574 68058
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 365514 367174 366134 402618
rect 365514 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 366134 367174
rect 365514 366854 366134 366938
rect 365514 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 366134 366854
rect 365514 331174 366134 366618
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 295174 366134 330618
rect 365514 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 366134 295174
rect 365514 294854 366134 294938
rect 365514 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 366134 294854
rect 365514 259174 366134 294618
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 223174 366134 258618
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 370894 369854 406338
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 369234 334894 369854 370338
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 369234 298894 369854 334338
rect 369234 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 369854 298894
rect 369234 298574 369854 298658
rect 369234 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 369854 298574
rect 369234 262894 369854 298338
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 226894 369854 262338
rect 369234 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 369854 226894
rect 369234 226574 369854 226658
rect 369234 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 369854 226574
rect 369234 190894 369854 226338
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 154894 369854 190338
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 338614 373574 374058
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 230614 373574 266058
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 565174 384134 600618
rect 383514 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 384134 565174
rect 383514 564854 384134 564938
rect 383514 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 384134 564854
rect 383514 529174 384134 564618
rect 383514 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 384134 529174
rect 383514 528854 384134 528938
rect 383514 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 384134 528854
rect 383514 493174 384134 528618
rect 383514 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 384134 493174
rect 383514 492854 384134 492938
rect 383514 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 384134 492854
rect 383514 457174 384134 492618
rect 383514 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 384134 457174
rect 383514 456854 384134 456938
rect 383514 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 384134 456854
rect 383514 421174 384134 456618
rect 383514 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 384134 421174
rect 383514 420854 384134 420938
rect 383514 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 384134 420854
rect 383514 385174 384134 420618
rect 383514 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 384134 385174
rect 383514 384854 384134 384938
rect 383514 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 384134 384854
rect 383514 349174 384134 384618
rect 383514 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 384134 349174
rect 383514 348854 384134 348938
rect 383514 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 384134 348854
rect 383514 313174 384134 348618
rect 383514 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 384134 313174
rect 383514 312854 384134 312938
rect 383514 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 384134 312854
rect 383514 277174 384134 312618
rect 383514 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 384134 277174
rect 383514 276854 384134 276938
rect 383514 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 384134 276854
rect 383514 241174 384134 276618
rect 383514 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 384134 241174
rect 383514 240854 384134 240938
rect 383514 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 384134 240854
rect 383514 205174 384134 240618
rect 383514 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 384134 205174
rect 383514 204854 384134 204938
rect 383514 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 384134 204854
rect 383514 169174 384134 204618
rect 383514 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 384134 169174
rect 383514 168854 384134 168938
rect 383514 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 384134 168854
rect 383514 133174 384134 168618
rect 383514 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 384134 133174
rect 383514 132854 384134 132938
rect 383514 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 384134 132854
rect 383514 97174 384134 132618
rect 383514 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 384134 97174
rect 383514 96854 384134 96938
rect 383514 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 384134 96854
rect 383514 61174 384134 96618
rect 383514 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 384134 61174
rect 383514 60854 384134 60938
rect 383514 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 384134 60854
rect 383514 25174 384134 60618
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 568894 387854 604338
rect 387234 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 387854 568894
rect 387234 568574 387854 568658
rect 387234 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 387854 568574
rect 387234 532894 387854 568338
rect 387234 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 387854 532894
rect 387234 532574 387854 532658
rect 387234 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 387854 532574
rect 387234 496894 387854 532338
rect 387234 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 387854 496894
rect 387234 496574 387854 496658
rect 387234 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 387854 496574
rect 387234 460894 387854 496338
rect 387234 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 387854 460894
rect 387234 460574 387854 460658
rect 387234 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 387854 460574
rect 387234 424894 387854 460338
rect 387234 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 387854 424894
rect 387234 424574 387854 424658
rect 387234 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 387854 424574
rect 387234 388894 387854 424338
rect 387234 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 387854 388894
rect 387234 388574 387854 388658
rect 387234 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 387854 388574
rect 387234 352894 387854 388338
rect 387234 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 387854 352894
rect 387234 352574 387854 352658
rect 387234 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 387854 352574
rect 387234 316894 387854 352338
rect 387234 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 387854 316894
rect 387234 316574 387854 316658
rect 387234 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 387854 316574
rect 387234 280894 387854 316338
rect 387234 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 387854 280894
rect 387234 280574 387854 280658
rect 387234 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 387854 280574
rect 387234 244894 387854 280338
rect 387234 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 387854 244894
rect 387234 244574 387854 244658
rect 387234 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 387854 244574
rect 387234 208894 387854 244338
rect 387234 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 387854 208894
rect 387234 208574 387854 208658
rect 387234 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 387854 208574
rect 387234 172894 387854 208338
rect 387234 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 387854 172894
rect 387234 172574 387854 172658
rect 387234 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 387854 172574
rect 387234 136894 387854 172338
rect 387234 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 387854 136894
rect 387234 136574 387854 136658
rect 387234 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 387854 136574
rect 387234 100894 387854 136338
rect 387234 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 387854 100894
rect 387234 100574 387854 100658
rect 387234 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 387854 100574
rect 387234 64894 387854 100338
rect 387234 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 387854 64894
rect 387234 64574 387854 64658
rect 387234 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 387854 64574
rect 387234 28894 387854 64338
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 390954 536614 391574 572058
rect 390954 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 391574 536614
rect 390954 536294 391574 536378
rect 390954 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 391574 536294
rect 390954 500614 391574 536058
rect 390954 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 391574 500614
rect 390954 500294 391574 500378
rect 390954 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 391574 500294
rect 390954 464614 391574 500058
rect 390954 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 391574 464614
rect 390954 464294 391574 464378
rect 390954 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 391574 464294
rect 390954 428614 391574 464058
rect 390954 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 391574 428614
rect 390954 428294 391574 428378
rect 390954 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 391574 428294
rect 390954 392614 391574 428058
rect 390954 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 391574 392614
rect 390954 392294 391574 392378
rect 390954 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 391574 392294
rect 390954 356614 391574 392058
rect 390954 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 391574 356614
rect 390954 356294 391574 356378
rect 390954 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 391574 356294
rect 390954 320614 391574 356058
rect 390954 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 391574 320614
rect 390954 320294 391574 320378
rect 390954 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 391574 320294
rect 390954 284614 391574 320058
rect 390954 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 391574 284614
rect 390954 284294 391574 284378
rect 390954 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 391574 284294
rect 390954 248614 391574 284058
rect 390954 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 391574 248614
rect 390954 248294 391574 248378
rect 390954 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 391574 248294
rect 390954 212614 391574 248058
rect 390954 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 391574 212614
rect 390954 212294 391574 212378
rect 390954 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 391574 212294
rect 390954 176614 391574 212058
rect 390954 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 391574 176614
rect 390954 176294 391574 176378
rect 390954 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 391574 176294
rect 390954 140614 391574 176058
rect 390954 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 391574 140614
rect 390954 140294 391574 140378
rect 390954 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 391574 140294
rect 390954 104614 391574 140058
rect 390954 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 391574 104614
rect 390954 104294 391574 104378
rect 390954 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 391574 104294
rect 390954 68614 391574 104058
rect 390954 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 391574 68614
rect 390954 68294 391574 68378
rect 390954 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 391574 68294
rect 390954 32614 391574 68058
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 439174 402134 474618
rect 401514 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 402134 439174
rect 401514 438854 402134 438938
rect 401514 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 402134 438854
rect 401514 403174 402134 438618
rect 401514 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 402134 403174
rect 401514 402854 402134 402938
rect 401514 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 402134 402854
rect 401514 367174 402134 402618
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 331174 402134 366618
rect 401514 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 402134 331174
rect 401514 330854 402134 330938
rect 401514 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 402134 330854
rect 401514 295174 402134 330618
rect 401514 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 402134 295174
rect 401514 294854 402134 294938
rect 401514 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 402134 294854
rect 401514 259174 402134 294618
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 223174 402134 258618
rect 401514 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 402134 223174
rect 401514 222854 402134 222938
rect 401514 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 402134 222854
rect 401514 187174 402134 222618
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 151174 402134 186618
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 79174 402134 114618
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 442894 405854 478338
rect 405234 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 405854 442894
rect 405234 442574 405854 442658
rect 405234 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 405854 442574
rect 405234 406894 405854 442338
rect 405234 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 405854 406894
rect 405234 406574 405854 406658
rect 405234 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 405854 406574
rect 405234 370894 405854 406338
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 334894 405854 370338
rect 405234 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 405854 334894
rect 405234 334574 405854 334658
rect 405234 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 405854 334574
rect 405234 298894 405854 334338
rect 405234 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 405854 298894
rect 405234 298574 405854 298658
rect 405234 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 405854 298574
rect 405234 262894 405854 298338
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 226894 405854 262338
rect 405234 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 405854 226894
rect 405234 226574 405854 226658
rect 405234 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 405854 226574
rect 405234 190894 405854 226338
rect 405234 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 405854 190894
rect 405234 190574 405854 190658
rect 405234 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 405854 190574
rect 405234 154894 405854 190338
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 118894 405854 154338
rect 405234 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 405854 118894
rect 405234 118574 405854 118658
rect 405234 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 405854 118574
rect 405234 82894 405854 118338
rect 405234 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 405854 82894
rect 405234 82574 405854 82658
rect 405234 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 405854 82574
rect 405234 46894 405854 82338
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 446614 409574 482058
rect 408954 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 409574 446614
rect 408954 446294 409574 446378
rect 408954 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 409574 446294
rect 408954 410614 409574 446058
rect 408954 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 409574 410614
rect 408954 410294 409574 410378
rect 408954 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 409574 410294
rect 408954 374614 409574 410058
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 408954 338614 409574 374058
rect 408954 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 409574 338614
rect 408954 338294 409574 338378
rect 408954 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 409574 338294
rect 408954 302614 409574 338058
rect 408954 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 409574 302614
rect 408954 302294 409574 302378
rect 408954 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 409574 302294
rect 408954 266614 409574 302058
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 230614 409574 266058
rect 408954 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 409574 230614
rect 408954 230294 409574 230378
rect 408954 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 409574 230294
rect 408954 194614 409574 230058
rect 408954 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 409574 194614
rect 408954 194294 409574 194378
rect 408954 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 409574 194294
rect 408954 158614 409574 194058
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 122614 409574 158058
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 408954 86614 409574 122058
rect 408954 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 409574 86614
rect 408954 86294 409574 86378
rect 408954 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 409574 86294
rect 408954 50614 409574 86058
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 565174 420134 600618
rect 419514 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 420134 565174
rect 419514 564854 420134 564938
rect 419514 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 420134 564854
rect 419514 529174 420134 564618
rect 419514 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 420134 529174
rect 419514 528854 420134 528938
rect 419514 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 420134 528854
rect 419514 493174 420134 528618
rect 419514 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 420134 493174
rect 419514 492854 420134 492938
rect 419514 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 420134 492854
rect 419514 457174 420134 492618
rect 419514 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 420134 457174
rect 419514 456854 420134 456938
rect 419514 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 420134 456854
rect 419514 421174 420134 456618
rect 419514 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 420134 421174
rect 419514 420854 420134 420938
rect 419514 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 420134 420854
rect 419514 385174 420134 420618
rect 419514 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 420134 385174
rect 419514 384854 420134 384938
rect 419514 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 420134 384854
rect 419514 349174 420134 384618
rect 419514 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 420134 349174
rect 419514 348854 420134 348938
rect 419514 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 420134 348854
rect 419514 313174 420134 348618
rect 419514 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 420134 313174
rect 419514 312854 420134 312938
rect 419514 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 420134 312854
rect 419514 277174 420134 312618
rect 419514 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 420134 277174
rect 419514 276854 420134 276938
rect 419514 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 420134 276854
rect 419514 241174 420134 276618
rect 419514 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 420134 241174
rect 419514 240854 420134 240938
rect 419514 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 420134 240854
rect 419514 205174 420134 240618
rect 419514 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 420134 205174
rect 419514 204854 420134 204938
rect 419514 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 420134 204854
rect 419514 169174 420134 204618
rect 419514 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 420134 169174
rect 419514 168854 420134 168938
rect 419514 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 420134 168854
rect 419514 133174 420134 168618
rect 419514 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 420134 133174
rect 419514 132854 420134 132938
rect 419514 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 420134 132854
rect 419514 97174 420134 132618
rect 419514 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 420134 97174
rect 419514 96854 420134 96938
rect 419514 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 420134 96854
rect 419514 61174 420134 96618
rect 419514 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 420134 61174
rect 419514 60854 420134 60938
rect 419514 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 420134 60854
rect 419514 25174 420134 60618
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 568894 423854 604338
rect 423234 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 423854 568894
rect 423234 568574 423854 568658
rect 423234 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 423854 568574
rect 423234 532894 423854 568338
rect 423234 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 423854 532894
rect 423234 532574 423854 532658
rect 423234 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 423854 532574
rect 423234 496894 423854 532338
rect 423234 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 423854 496894
rect 423234 496574 423854 496658
rect 423234 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 423854 496574
rect 423234 460894 423854 496338
rect 423234 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 423854 460894
rect 423234 460574 423854 460658
rect 423234 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 423854 460574
rect 423234 424894 423854 460338
rect 423234 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 423854 424894
rect 423234 424574 423854 424658
rect 423234 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 423854 424574
rect 423234 388894 423854 424338
rect 423234 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 423854 388894
rect 423234 388574 423854 388658
rect 423234 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 423854 388574
rect 423234 352894 423854 388338
rect 423234 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 423854 352894
rect 423234 352574 423854 352658
rect 423234 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 423854 352574
rect 423234 316894 423854 352338
rect 423234 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 423854 316894
rect 423234 316574 423854 316658
rect 423234 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 423854 316574
rect 423234 280894 423854 316338
rect 423234 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 423854 280894
rect 423234 280574 423854 280658
rect 423234 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 423854 280574
rect 423234 244894 423854 280338
rect 423234 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 423854 244894
rect 423234 244574 423854 244658
rect 423234 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 423854 244574
rect 423234 208894 423854 244338
rect 423234 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 423854 208894
rect 423234 208574 423854 208658
rect 423234 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 423854 208574
rect 423234 172894 423854 208338
rect 423234 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 423854 172894
rect 423234 172574 423854 172658
rect 423234 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 423854 172574
rect 423234 136894 423854 172338
rect 423234 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 423854 136894
rect 423234 136574 423854 136658
rect 423234 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 423854 136574
rect 423234 100894 423854 136338
rect 423234 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 423854 100894
rect 423234 100574 423854 100658
rect 423234 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 423854 100574
rect 423234 64894 423854 100338
rect 423234 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 423854 64894
rect 423234 64574 423854 64658
rect 423234 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 423854 64574
rect 423234 28894 423854 64338
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 572614 427574 608058
rect 426954 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 427574 572614
rect 426954 572294 427574 572378
rect 426954 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 427574 572294
rect 426954 536614 427574 572058
rect 426954 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 427574 536614
rect 426954 536294 427574 536378
rect 426954 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 427574 536294
rect 426954 500614 427574 536058
rect 426954 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 427574 500614
rect 426954 500294 427574 500378
rect 426954 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 427574 500294
rect 426954 464614 427574 500058
rect 426954 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 427574 464614
rect 426954 464294 427574 464378
rect 426954 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 427574 464294
rect 426954 428614 427574 464058
rect 426954 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 427574 428614
rect 426954 428294 427574 428378
rect 426954 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 427574 428294
rect 426954 392614 427574 428058
rect 426954 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 427574 392614
rect 426954 392294 427574 392378
rect 426954 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 427574 392294
rect 426954 356614 427574 392058
rect 426954 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 427574 356614
rect 426954 356294 427574 356378
rect 426954 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 427574 356294
rect 426954 320614 427574 356058
rect 426954 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 427574 320614
rect 426954 320294 427574 320378
rect 426954 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 427574 320294
rect 426954 284614 427574 320058
rect 426954 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 427574 284614
rect 426954 284294 427574 284378
rect 426954 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 427574 284294
rect 426954 248614 427574 284058
rect 426954 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 427574 248614
rect 426954 248294 427574 248378
rect 426954 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 427574 248294
rect 426954 212614 427574 248058
rect 426954 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 427574 212614
rect 426954 212294 427574 212378
rect 426954 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 427574 212294
rect 426954 176614 427574 212058
rect 426954 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 427574 176614
rect 426954 176294 427574 176378
rect 426954 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 427574 176294
rect 426954 140614 427574 176058
rect 426954 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 427574 140614
rect 426954 140294 427574 140378
rect 426954 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 427574 140294
rect 426954 104614 427574 140058
rect 426954 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 427574 104614
rect 426954 104294 427574 104378
rect 426954 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 427574 104294
rect 426954 68614 427574 104058
rect 426954 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 427574 68614
rect 426954 68294 427574 68378
rect 426954 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 427574 68294
rect 426954 32614 427574 68058
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 439174 438134 474618
rect 437514 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 438134 439174
rect 437514 438854 438134 438938
rect 437514 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 438134 438854
rect 437514 403174 438134 438618
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 437514 367174 438134 402618
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 331174 438134 366618
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 295174 438134 330618
rect 437514 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 438134 295174
rect 437514 294854 438134 294938
rect 437514 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 438134 294854
rect 437514 259174 438134 294618
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 223174 438134 258618
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 187174 438134 222618
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 151174 438134 186618
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 437514 115174 438134 150618
rect 437514 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 438134 115174
rect 437514 114854 438134 114938
rect 437514 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 438134 114854
rect 437514 79174 438134 114618
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 442894 441854 478338
rect 441234 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 441854 442894
rect 441234 442574 441854 442658
rect 441234 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 441854 442574
rect 441234 406894 441854 442338
rect 441234 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 441854 406894
rect 441234 406574 441854 406658
rect 441234 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 441854 406574
rect 441234 370894 441854 406338
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 334894 441854 370338
rect 441234 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 441854 334894
rect 441234 334574 441854 334658
rect 441234 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 441854 334574
rect 441234 298894 441854 334338
rect 441234 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 441854 298894
rect 441234 298574 441854 298658
rect 441234 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 441854 298574
rect 441234 262894 441854 298338
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 226894 441854 262338
rect 441234 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 441854 226894
rect 441234 226574 441854 226658
rect 441234 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 441854 226574
rect 441234 190894 441854 226338
rect 441234 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 441854 190894
rect 441234 190574 441854 190658
rect 441234 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 441854 190574
rect 441234 154894 441854 190338
rect 441234 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 441854 154894
rect 441234 154574 441854 154658
rect 441234 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 441854 154574
rect 441234 118894 441854 154338
rect 441234 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 441854 118894
rect 441234 118574 441854 118658
rect 441234 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 441854 118574
rect 441234 82894 441854 118338
rect 441234 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 441854 82894
rect 441234 82574 441854 82658
rect 441234 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 441854 82574
rect 441234 46894 441854 82338
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 444954 410614 445574 446058
rect 444954 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 445574 410614
rect 444954 410294 445574 410378
rect 444954 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 445574 410294
rect 444954 374614 445574 410058
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 444954 338614 445574 374058
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 444954 302614 445574 338058
rect 444954 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 445574 302614
rect 444954 302294 445574 302378
rect 444954 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 445574 302294
rect 444954 266614 445574 302058
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 230614 445574 266058
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 444954 158614 445574 194058
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 444954 122614 445574 158058
rect 444954 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 445574 122614
rect 444954 122294 445574 122378
rect 444954 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 445574 122294
rect 444954 86614 445574 122058
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 444954 50614 445574 86058
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 529174 456134 564618
rect 455514 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 456134 529174
rect 455514 528854 456134 528938
rect 455514 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 456134 528854
rect 455514 493174 456134 528618
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 455514 457174 456134 492618
rect 455514 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 456134 457174
rect 455514 456854 456134 456938
rect 455514 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 456134 456854
rect 455514 421174 456134 456618
rect 455514 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 456134 421174
rect 455514 420854 456134 420938
rect 455514 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 456134 420854
rect 455514 385174 456134 420618
rect 455514 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 456134 385174
rect 455514 384854 456134 384938
rect 455514 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 456134 384854
rect 455514 349174 456134 384618
rect 455514 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 456134 349174
rect 455514 348854 456134 348938
rect 455514 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 456134 348854
rect 455514 313174 456134 348618
rect 455514 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 456134 313174
rect 455514 312854 456134 312938
rect 455514 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 456134 312854
rect 455514 277174 456134 312618
rect 455514 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 456134 277174
rect 455514 276854 456134 276938
rect 455514 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 456134 276854
rect 455514 241174 456134 276618
rect 455514 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 456134 241174
rect 455514 240854 456134 240938
rect 455514 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 456134 240854
rect 455514 205174 456134 240618
rect 455514 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 456134 205174
rect 455514 204854 456134 204938
rect 455514 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 456134 204854
rect 455514 169174 456134 204618
rect 455514 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 456134 169174
rect 455514 168854 456134 168938
rect 455514 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 456134 168854
rect 455514 133174 456134 168618
rect 455514 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 456134 133174
rect 455514 132854 456134 132938
rect 455514 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 456134 132854
rect 455514 97174 456134 132618
rect 455514 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 456134 97174
rect 455514 96854 456134 96938
rect 455514 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 456134 96854
rect 455514 61174 456134 96618
rect 455514 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 456134 61174
rect 455514 60854 456134 60938
rect 455514 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 456134 60854
rect 455514 25174 456134 60618
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 568894 459854 604338
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 532894 459854 568338
rect 459234 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 459854 532894
rect 459234 532574 459854 532658
rect 459234 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 459854 532574
rect 459234 496894 459854 532338
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 460894 459854 496338
rect 459234 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 459854 460894
rect 459234 460574 459854 460658
rect 459234 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 459854 460574
rect 459234 424894 459854 460338
rect 459234 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 459854 424894
rect 459234 424574 459854 424658
rect 459234 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 459854 424574
rect 459234 388894 459854 424338
rect 459234 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 459854 388894
rect 459234 388574 459854 388658
rect 459234 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 459854 388574
rect 459234 352894 459854 388338
rect 459234 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 459854 352894
rect 459234 352574 459854 352658
rect 459234 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 459854 352574
rect 459234 316894 459854 352338
rect 459234 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 459854 316894
rect 459234 316574 459854 316658
rect 459234 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 459854 316574
rect 459234 280894 459854 316338
rect 459234 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 459854 280894
rect 459234 280574 459854 280658
rect 459234 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 459854 280574
rect 459234 244894 459854 280338
rect 459234 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 459854 244894
rect 459234 244574 459854 244658
rect 459234 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 459854 244574
rect 459234 208894 459854 244338
rect 459234 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 459854 208894
rect 459234 208574 459854 208658
rect 459234 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 459854 208574
rect 459234 172894 459854 208338
rect 459234 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 459854 172894
rect 459234 172574 459854 172658
rect 459234 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 459854 172574
rect 459234 136894 459854 172338
rect 459234 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 459854 136894
rect 459234 136574 459854 136658
rect 459234 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 459854 136574
rect 459234 100894 459854 136338
rect 459234 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 459854 100894
rect 459234 100574 459854 100658
rect 459234 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 459854 100574
rect 459234 64894 459854 100338
rect 459234 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 459854 64894
rect 459234 64574 459854 64658
rect 459234 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 459854 64574
rect 459234 28894 459854 64338
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 572614 463574 608058
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 536614 463574 572058
rect 462954 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 463574 536614
rect 462954 536294 463574 536378
rect 462954 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 463574 536294
rect 462954 500614 463574 536058
rect 462954 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 463574 500614
rect 462954 500294 463574 500378
rect 462954 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 463574 500294
rect 462954 464614 463574 500058
rect 462954 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 463574 464614
rect 462954 464294 463574 464378
rect 462954 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 463574 464294
rect 462954 428614 463574 464058
rect 462954 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 463574 428614
rect 462954 428294 463574 428378
rect 462954 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 463574 428294
rect 462954 392614 463574 428058
rect 462954 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 463574 392614
rect 462954 392294 463574 392378
rect 462954 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 463574 392294
rect 462954 356614 463574 392058
rect 462954 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 463574 356614
rect 462954 356294 463574 356378
rect 462954 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 463574 356294
rect 462954 320614 463574 356058
rect 462954 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 463574 320614
rect 462954 320294 463574 320378
rect 462954 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 463574 320294
rect 462954 284614 463574 320058
rect 462954 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 463574 284614
rect 462954 284294 463574 284378
rect 462954 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 463574 284294
rect 462954 248614 463574 284058
rect 462954 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 463574 248614
rect 462954 248294 463574 248378
rect 462954 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 463574 248294
rect 462954 212614 463574 248058
rect 462954 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 463574 212614
rect 462954 212294 463574 212378
rect 462954 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 463574 212294
rect 462954 176614 463574 212058
rect 462954 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 463574 176614
rect 462954 176294 463574 176378
rect 462954 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 463574 176294
rect 462954 140614 463574 176058
rect 462954 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 463574 140614
rect 462954 140294 463574 140378
rect 462954 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 463574 140294
rect 462954 104614 463574 140058
rect 462954 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 463574 104614
rect 462954 104294 463574 104378
rect 462954 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 463574 104294
rect 462954 68614 463574 104058
rect 462954 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 463574 68614
rect 462954 68294 463574 68378
rect 462954 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 463574 68294
rect 462954 32614 463574 68058
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 439174 474134 474618
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 473514 403174 474134 438618
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 473514 367174 474134 402618
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 331174 474134 366618
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 473514 295174 474134 330618
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 473514 259174 474134 294618
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 223174 474134 258618
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 406894 477854 442338
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 477234 370894 477854 406338
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 334894 477854 370338
rect 477234 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 477854 334894
rect 477234 334574 477854 334658
rect 477234 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 477854 334574
rect 477234 298894 477854 334338
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 226894 477854 262338
rect 477234 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 477854 226894
rect 477234 226574 477854 226658
rect 477234 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 477854 226574
rect 477234 190894 477854 226338
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 446614 481574 482058
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 480954 410614 481574 446058
rect 480954 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 481574 410614
rect 480954 410294 481574 410378
rect 480954 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 481574 410294
rect 480954 374614 481574 410058
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 480954 338614 481574 374058
rect 480954 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 481574 338614
rect 480954 338294 481574 338378
rect 480954 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 481574 338294
rect 480954 302614 481574 338058
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 480954 266614 481574 302058
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 230614 481574 266058
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 480954 194614 481574 230058
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 601174 492134 636618
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 565174 492134 600618
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 491514 457174 492134 492618
rect 491514 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 492134 457174
rect 491514 456854 492134 456938
rect 491514 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 492134 456854
rect 491514 421174 492134 456618
rect 491514 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 492134 421174
rect 491514 420854 492134 420938
rect 491514 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 492134 420854
rect 491514 385174 492134 420618
rect 491514 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 492134 385174
rect 491514 384854 492134 384938
rect 491514 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 492134 384854
rect 491514 349174 492134 384618
rect 491514 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 492134 349174
rect 491514 348854 492134 348938
rect 491514 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 492134 348854
rect 491514 313174 492134 348618
rect 491514 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 492134 313174
rect 491514 312854 492134 312938
rect 491514 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 492134 312854
rect 491514 277174 492134 312618
rect 491514 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 492134 277174
rect 491514 276854 492134 276938
rect 491514 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 492134 276854
rect 491514 241174 492134 276618
rect 491514 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 492134 241174
rect 491514 240854 492134 240938
rect 491514 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 492134 240854
rect 491514 205174 492134 240618
rect 491514 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 492134 205174
rect 491514 204854 492134 204938
rect 491514 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 492134 204854
rect 491514 169174 492134 204618
rect 491514 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 492134 169174
rect 491514 168854 492134 168938
rect 491514 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 492134 168854
rect 491514 133174 492134 168618
rect 491514 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 492134 133174
rect 491514 132854 492134 132938
rect 491514 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 492134 132854
rect 491514 97174 492134 132618
rect 491514 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 492134 97174
rect 491514 96854 492134 96938
rect 491514 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 492134 96854
rect 491514 61174 492134 96618
rect 491514 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 492134 61174
rect 491514 60854 492134 60938
rect 491514 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 492134 60854
rect 491514 25174 492134 60618
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 604894 495854 640338
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 568894 495854 604338
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 532894 495854 568338
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 460894 495854 496338
rect 495234 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 495854 460894
rect 495234 460574 495854 460658
rect 495234 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 495854 460574
rect 495234 424894 495854 460338
rect 495234 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 495854 424894
rect 495234 424574 495854 424658
rect 495234 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 495854 424574
rect 495234 388894 495854 424338
rect 495234 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 495854 388894
rect 495234 388574 495854 388658
rect 495234 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 495854 388574
rect 495234 352894 495854 388338
rect 495234 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 495854 352894
rect 495234 352574 495854 352658
rect 495234 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 495854 352574
rect 495234 316894 495854 352338
rect 495234 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 495854 316894
rect 495234 316574 495854 316658
rect 495234 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 495854 316574
rect 495234 280894 495854 316338
rect 495234 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 495854 280894
rect 495234 280574 495854 280658
rect 495234 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 495854 280574
rect 495234 244894 495854 280338
rect 495234 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 495854 244894
rect 495234 244574 495854 244658
rect 495234 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 495854 244574
rect 495234 208894 495854 244338
rect 495234 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 495854 208894
rect 495234 208574 495854 208658
rect 495234 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 495854 208574
rect 495234 172894 495854 208338
rect 495234 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 495854 172894
rect 495234 172574 495854 172658
rect 495234 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 495854 172574
rect 495234 136894 495854 172338
rect 495234 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 495854 136894
rect 495234 136574 495854 136658
rect 495234 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 495854 136574
rect 495234 100894 495854 136338
rect 495234 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 495854 100894
rect 495234 100574 495854 100658
rect 495234 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 495854 100574
rect 495234 64894 495854 100338
rect 495234 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 495854 64894
rect 495234 64574 495854 64658
rect 495234 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 495854 64574
rect 495234 28894 495854 64338
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 608614 499574 644058
rect 498954 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 499574 608614
rect 498954 608294 499574 608378
rect 498954 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 499574 608294
rect 498954 572614 499574 608058
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 536614 499574 572058
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498954 464614 499574 500058
rect 498954 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 499574 464614
rect 498954 464294 499574 464378
rect 498954 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 499574 464294
rect 498954 428614 499574 464058
rect 498954 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 499574 428614
rect 498954 428294 499574 428378
rect 498954 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 499574 428294
rect 498954 392614 499574 428058
rect 498954 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 499574 392614
rect 498954 392294 499574 392378
rect 498954 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 499574 392294
rect 498954 356614 499574 392058
rect 498954 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 499574 356614
rect 498954 356294 499574 356378
rect 498954 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 499574 356294
rect 498954 320614 499574 356058
rect 498954 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 499574 320614
rect 498954 320294 499574 320378
rect 498954 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 499574 320294
rect 498954 284614 499574 320058
rect 498954 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 499574 284614
rect 498954 284294 499574 284378
rect 498954 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 499574 284294
rect 498954 248614 499574 284058
rect 498954 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 499574 248614
rect 498954 248294 499574 248378
rect 498954 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 499574 248294
rect 498954 212614 499574 248058
rect 498954 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 499574 212614
rect 498954 212294 499574 212378
rect 498954 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 499574 212294
rect 498954 176614 499574 212058
rect 498954 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 499574 176614
rect 498954 176294 499574 176378
rect 498954 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 499574 176294
rect 498954 140614 499574 176058
rect 498954 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 499574 140614
rect 498954 140294 499574 140378
rect 498954 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 499574 140294
rect 498954 104614 499574 140058
rect 498954 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 499574 104614
rect 498954 104294 499574 104378
rect 498954 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 499574 104294
rect 498954 68614 499574 104058
rect 498954 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 499574 68614
rect 498954 68294 499574 68378
rect 498954 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 499574 68294
rect 498954 32614 499574 68058
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509514 295174 510134 330618
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 513234 298894 513854 334338
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 513234 262894 513854 298338
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 516954 302614 517574 338058
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 516954 266614 517574 302058
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 59546 456938 59782 457174
rect 59866 456938 60102 457174
rect 59546 456618 59782 456854
rect 59866 456618 60102 456854
rect 59546 420938 59782 421174
rect 59866 420938 60102 421174
rect 59546 420618 59782 420854
rect 59866 420618 60102 420854
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 59546 384938 59782 385174
rect 59866 384938 60102 385174
rect 59546 384618 59782 384854
rect 59866 384618 60102 384854
rect 59546 348938 59782 349174
rect 59866 348938 60102 349174
rect 59546 348618 59782 348854
rect 59866 348618 60102 348854
rect 59546 312938 59782 313174
rect 59866 312938 60102 313174
rect 59546 312618 59782 312854
rect 59866 312618 60102 312854
rect 59546 276938 59782 277174
rect 59866 276938 60102 277174
rect 59546 276618 59782 276854
rect 59866 276618 60102 276854
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 63266 460658 63502 460894
rect 63586 460658 63822 460894
rect 63266 460338 63502 460574
rect 63586 460338 63822 460574
rect 66986 536378 67222 536614
rect 67306 536378 67542 536614
rect 66986 536058 67222 536294
rect 67306 536058 67542 536294
rect 66986 500378 67222 500614
rect 67306 500378 67542 500614
rect 66986 500058 67222 500294
rect 67306 500058 67542 500294
rect 73721 543218 73957 543454
rect 73721 542898 73957 543134
rect 66986 464378 67222 464614
rect 67306 464378 67542 464614
rect 66986 464058 67222 464294
rect 67306 464058 67542 464294
rect 63266 424658 63502 424894
rect 63586 424658 63822 424894
rect 63266 424338 63502 424574
rect 63586 424338 63822 424574
rect 63266 388658 63502 388894
rect 63586 388658 63822 388894
rect 63266 388338 63502 388574
rect 63586 388338 63822 388574
rect 63266 352658 63502 352894
rect 63586 352658 63822 352894
rect 63266 352338 63502 352574
rect 63586 352338 63822 352574
rect 66986 356378 67222 356614
rect 67306 356378 67542 356614
rect 66986 356058 67222 356294
rect 67306 356058 67542 356294
rect 63266 316658 63502 316894
rect 63586 316658 63822 316894
rect 63266 316338 63502 316574
rect 63586 316338 63822 316574
rect 63266 280658 63502 280894
rect 63586 280658 63822 280894
rect 63266 280338 63502 280574
rect 63586 280338 63822 280574
rect 59546 240938 59782 241174
rect 59866 240938 60102 241174
rect 59546 240618 59782 240854
rect 59866 240618 60102 240854
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 63266 244658 63502 244894
rect 63586 244658 63822 244894
rect 63266 244338 63502 244574
rect 63586 244338 63822 244574
rect 59546 204938 59782 205174
rect 59866 204938 60102 205174
rect 59546 204618 59782 204854
rect 59866 204618 60102 204854
rect 59546 168938 59782 169174
rect 59866 168938 60102 169174
rect 59546 168618 59782 168854
rect 59866 168618 60102 168854
rect 59546 132938 59782 133174
rect 59866 132938 60102 133174
rect 59546 132618 59782 132854
rect 59866 132618 60102 132854
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 66986 320378 67222 320614
rect 67306 320378 67542 320614
rect 66986 320058 67222 320294
rect 67306 320058 67542 320294
rect 63266 208658 63502 208894
rect 63586 208658 63822 208894
rect 63266 208338 63502 208574
rect 63586 208338 63822 208574
rect 63266 172658 63502 172894
rect 63586 172658 63822 172894
rect 63266 172338 63502 172574
rect 63586 172338 63822 172574
rect 63266 136658 63502 136894
rect 63586 136658 63822 136894
rect 63266 136338 63502 136574
rect 63586 136338 63822 136574
rect 59546 96938 59782 97174
rect 59866 96938 60102 97174
rect 59546 96618 59782 96854
rect 59866 96618 60102 96854
rect 59546 60938 59782 61174
rect 59866 60938 60102 61174
rect 59546 60618 59782 60854
rect 59866 60618 60102 60854
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 100658 63502 100894
rect 63586 100658 63822 100894
rect 63266 100338 63502 100574
rect 63586 100338 63822 100574
rect 66986 212378 67222 212614
rect 67306 212378 67542 212614
rect 66986 212058 67222 212294
rect 67306 212058 67542 212294
rect 66986 176378 67222 176614
rect 67306 176378 67542 176614
rect 66986 176058 67222 176294
rect 67306 176058 67542 176294
rect 66986 140378 67222 140614
rect 67306 140378 67542 140614
rect 66986 140058 67222 140294
rect 67306 140058 67542 140294
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73020 399218 73256 399454
rect 73020 398898 73256 399134
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 81266 586658 81502 586894
rect 81586 586658 81822 586894
rect 81266 586338 81502 586574
rect 81586 586338 81822 586574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 84986 590378 85222 590614
rect 85306 590378 85542 590614
rect 84986 590058 85222 590294
rect 85306 590058 85542 590294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 77686 561218 77922 561454
rect 77686 560898 77922 561134
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 77546 438938 77782 439174
rect 77866 438938 78102 439174
rect 77546 438618 77782 438854
rect 77866 438618 78102 438854
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 81651 543218 81887 543454
rect 81651 542898 81887 543134
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 81266 442658 81502 442894
rect 81586 442658 81822 442894
rect 81266 442338 81502 442574
rect 81586 442338 81822 442574
rect 85617 561218 85853 561454
rect 85617 560898 85853 561134
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 84986 446378 85222 446614
rect 85306 446378 85542 446614
rect 84986 446058 85222 446294
rect 85306 446058 85542 446294
rect 77546 366938 77782 367174
rect 77866 366938 78102 367174
rect 77546 366618 77782 366854
rect 77866 366618 78102 366854
rect 77546 330938 77782 331174
rect 77866 330938 78102 331174
rect 77546 330618 77782 330854
rect 77866 330618 78102 330854
rect 77546 294938 77782 295174
rect 77866 294938 78102 295174
rect 77546 294618 77782 294854
rect 77866 294618 78102 294854
rect 81266 370658 81502 370894
rect 81586 370658 81822 370894
rect 81266 370338 81502 370574
rect 81586 370338 81822 370574
rect 81266 334658 81502 334894
rect 81586 334658 81822 334894
rect 81266 334338 81502 334574
rect 81586 334338 81822 334574
rect 81266 298658 81502 298894
rect 81586 298658 81822 298894
rect 81266 298338 81502 298574
rect 81586 298338 81822 298574
rect 84986 374378 85222 374614
rect 85306 374378 85542 374614
rect 84986 374058 85222 374294
rect 85306 374058 85542 374294
rect 84986 338378 85222 338614
rect 85306 338378 85542 338614
rect 84986 338058 85222 338294
rect 85306 338058 85542 338294
rect 84986 302378 85222 302614
rect 85306 302378 85542 302614
rect 84986 302058 85222 302294
rect 85306 302058 85542 302294
rect 79019 273218 79255 273454
rect 79019 272898 79255 273134
rect 74387 255218 74623 255454
rect 74387 254898 74623 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 77546 222938 77782 223174
rect 77866 222938 78102 223174
rect 77546 222618 77782 222854
rect 77866 222618 78102 222854
rect 77546 186938 77782 187174
rect 77866 186938 78102 187174
rect 77546 186618 77782 186854
rect 77866 186618 78102 186854
rect 77546 150938 77782 151174
rect 77866 150938 78102 151174
rect 77546 150618 77782 150854
rect 77866 150618 78102 150854
rect 81266 226658 81502 226894
rect 81586 226658 81822 226894
rect 81266 226338 81502 226574
rect 81586 226338 81822 226574
rect 81266 190658 81502 190894
rect 81586 190658 81822 190894
rect 81266 190338 81502 190574
rect 81586 190338 81822 190574
rect 81266 154658 81502 154894
rect 81586 154658 81822 154894
rect 81266 154338 81502 154574
rect 81586 154338 81822 154574
rect 83651 255218 83887 255454
rect 83651 254898 83887 255134
rect 88380 417218 88616 417454
rect 88380 416898 88616 417134
rect 89582 543218 89818 543454
rect 89582 542898 89818 543134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 99266 568658 99502 568894
rect 99586 568658 99822 568894
rect 99266 568338 99502 568574
rect 99586 568338 99822 568574
rect 95546 528938 95782 529174
rect 95866 528938 96102 529174
rect 95546 528618 95782 528854
rect 95866 528618 96102 528854
rect 95546 492938 95782 493174
rect 95866 492938 96102 493174
rect 95546 492618 95782 492854
rect 95866 492618 96102 492854
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 95546 456938 95782 457174
rect 95866 456938 96102 457174
rect 95546 456618 95782 456854
rect 95866 456618 96102 456854
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 84986 230378 85222 230614
rect 85306 230378 85542 230614
rect 84986 230058 85222 230294
rect 85306 230058 85542 230294
rect 84986 194378 85222 194614
rect 85306 194378 85542 194614
rect 84986 194058 85222 194294
rect 85306 194058 85542 194294
rect 88283 273218 88519 273454
rect 88283 272898 88519 273134
rect 92915 255218 93151 255454
rect 92915 254898 93151 255134
rect 99266 532658 99502 532894
rect 99586 532658 99822 532894
rect 99266 532338 99502 532574
rect 99586 532338 99822 532574
rect 99266 496658 99502 496894
rect 99586 496658 99822 496894
rect 99266 496338 99502 496574
rect 99586 496338 99822 496574
rect 95546 384938 95782 385174
rect 95866 384938 96102 385174
rect 95546 384618 95782 384854
rect 95866 384618 96102 384854
rect 99266 460658 99502 460894
rect 99586 460658 99822 460894
rect 99266 460338 99502 460574
rect 99586 460338 99822 460574
rect 95546 348938 95782 349174
rect 95866 348938 96102 349174
rect 95546 348618 95782 348854
rect 95866 348618 96102 348854
rect 95546 312938 95782 313174
rect 95866 312938 96102 313174
rect 95546 312618 95782 312854
rect 95866 312618 96102 312854
rect 99266 352658 99502 352894
rect 99586 352658 99822 352894
rect 99266 352338 99502 352574
rect 99586 352338 99822 352574
rect 99266 316658 99502 316894
rect 99586 316658 99822 316894
rect 99266 316338 99502 316574
rect 99586 316338 99822 316574
rect 102986 572378 103222 572614
rect 103306 572378 103542 572614
rect 102986 572058 103222 572294
rect 103306 572058 103542 572294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 102986 536378 103222 536614
rect 103306 536378 103542 536614
rect 102986 536058 103222 536294
rect 103306 536058 103542 536294
rect 102986 500378 103222 500614
rect 103306 500378 103542 500614
rect 102986 500058 103222 500294
rect 103306 500058 103542 500294
rect 102986 464378 103222 464614
rect 103306 464378 103542 464614
rect 102986 464058 103222 464294
rect 103306 464058 103542 464294
rect 103740 399218 103976 399454
rect 103740 398898 103976 399134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 102986 356378 103222 356614
rect 103306 356378 103542 356614
rect 102986 356058 103222 356294
rect 103306 356058 103542 356294
rect 102986 320378 103222 320614
rect 103306 320378 103542 320614
rect 102986 320058 103222 320294
rect 103306 320058 103542 320294
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 102986 284378 103222 284614
rect 103306 284378 103542 284614
rect 102986 284058 103222 284294
rect 103306 284058 103542 284294
rect 84986 158378 85222 158614
rect 85306 158378 85542 158614
rect 84986 158058 85222 158294
rect 85306 158058 85542 158294
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 77686 129218 77922 129454
rect 77686 128898 77922 129134
rect 85617 129218 85853 129454
rect 85617 128898 85853 129134
rect 73721 111218 73957 111454
rect 73721 110898 73957 111134
rect 81651 111218 81887 111454
rect 81651 110898 81887 111134
rect 89582 111218 89818 111454
rect 89582 110898 89818 111134
rect 95546 204938 95782 205174
rect 95866 204938 96102 205174
rect 95546 204618 95782 204854
rect 95866 204618 96102 204854
rect 95546 168938 95782 169174
rect 95866 168938 96102 169174
rect 95546 168618 95782 168854
rect 95866 168618 96102 168854
rect 63266 64658 63502 64894
rect 63586 64658 63822 64894
rect 63266 64338 63502 64574
rect 63586 64338 63822 64574
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 66986 68378 67222 68614
rect 67306 68378 67542 68614
rect 66986 68058 67222 68294
rect 67306 68058 67542 68294
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 78938 77782 79174
rect 77866 78938 78102 79174
rect 77546 78618 77782 78854
rect 77866 78618 78102 78854
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 82658 81502 82894
rect 81586 82658 81822 82894
rect 81266 82338 81502 82574
rect 81586 82338 81822 82574
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 86378 85222 86614
rect 85306 86378 85542 86614
rect 84986 86058 85222 86294
rect 85306 86058 85542 86294
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 99266 208658 99502 208894
rect 99586 208658 99822 208894
rect 99266 208338 99502 208574
rect 99586 208338 99822 208574
rect 99266 172658 99502 172894
rect 99586 172658 99822 172894
rect 99266 172338 99502 172574
rect 99586 172338 99822 172574
rect 99266 136658 99502 136894
rect 99586 136658 99822 136894
rect 99266 136338 99502 136574
rect 99586 136338 99822 136574
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 102986 248378 103222 248614
rect 103306 248378 103542 248614
rect 102986 248058 103222 248294
rect 103306 248058 103542 248294
rect 102986 212378 103222 212614
rect 103306 212378 103542 212614
rect 102986 212058 103222 212294
rect 103306 212058 103542 212294
rect 102986 176378 103222 176614
rect 103306 176378 103542 176614
rect 102986 176058 103222 176294
rect 103306 176058 103542 176294
rect 102986 140378 103222 140614
rect 103306 140378 103542 140614
rect 102986 140058 103222 140294
rect 103306 140058 103542 140294
rect 99266 100658 99502 100894
rect 99586 100658 99822 100894
rect 99266 100338 99502 100574
rect 99586 100338 99822 100574
rect 95546 60938 95782 61174
rect 95866 60938 96102 61174
rect 95546 60618 95782 60854
rect 95866 60618 96102 60854
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 64658 99502 64894
rect 99586 64658 99822 64894
rect 99266 64338 99502 64574
rect 99586 64338 99822 64574
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 102986 104378 103222 104614
rect 103306 104378 103542 104614
rect 102986 104058 103222 104294
rect 103306 104058 103542 104294
rect 102986 68378 103222 68614
rect 103306 68378 103542 68614
rect 102986 68058 103222 68294
rect 103306 68058 103542 68294
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 113546 438938 113782 439174
rect 113866 438938 114102 439174
rect 113546 438618 113782 438854
rect 113866 438618 114102 438854
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 117266 442658 117502 442894
rect 117586 442658 117822 442894
rect 117266 442338 117502 442574
rect 117586 442338 117822 442574
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 120986 446378 121222 446614
rect 121306 446378 121542 446614
rect 120986 446058 121222 446294
rect 121306 446058 121542 446294
rect 117266 406658 117502 406894
rect 117586 406658 117822 406894
rect 117266 406338 117502 406574
rect 117586 406338 117822 406574
rect 113546 366938 113782 367174
rect 113866 366938 114102 367174
rect 113546 366618 113782 366854
rect 113866 366618 114102 366854
rect 113546 330938 113782 331174
rect 113866 330938 114102 331174
rect 113546 330618 113782 330854
rect 113866 330618 114102 330854
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 113546 294938 113782 295174
rect 113866 294938 114102 295174
rect 113546 294618 113782 294854
rect 113866 294618 114102 294854
rect 113546 258938 113782 259174
rect 113866 258938 114102 259174
rect 113546 258618 113782 258854
rect 113866 258618 114102 258854
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 113546 222938 113782 223174
rect 113866 222938 114102 223174
rect 113546 222618 113782 222854
rect 113866 222618 114102 222854
rect 113546 186938 113782 187174
rect 113866 186938 114102 187174
rect 113546 186618 113782 186854
rect 113866 186618 114102 186854
rect 113546 150938 113782 151174
rect 113866 150938 114102 151174
rect 113546 150618 113782 150854
rect 113866 150618 114102 150854
rect 113546 114938 113782 115174
rect 113866 114938 114102 115174
rect 113546 114618 113782 114854
rect 113866 114618 114102 114854
rect 113546 78938 113782 79174
rect 113866 78938 114102 79174
rect 113546 78618 113782 78854
rect 113866 78618 114102 78854
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 370658 117502 370894
rect 117586 370658 117822 370894
rect 117266 370338 117502 370574
rect 117586 370338 117822 370574
rect 117266 334658 117502 334894
rect 117586 334658 117822 334894
rect 117266 334338 117502 334574
rect 117586 334338 117822 334574
rect 120986 410378 121222 410614
rect 121306 410378 121542 410614
rect 120986 410058 121222 410294
rect 121306 410058 121542 410294
rect 120986 374378 121222 374614
rect 121306 374378 121542 374614
rect 120986 374058 121222 374294
rect 121306 374058 121542 374294
rect 120986 338378 121222 338614
rect 121306 338378 121542 338614
rect 120986 338058 121222 338294
rect 121306 338058 121542 338294
rect 117266 298658 117502 298894
rect 117586 298658 117822 298894
rect 117266 298338 117502 298574
rect 117586 298338 117822 298574
rect 117266 262658 117502 262894
rect 117586 262658 117822 262894
rect 117266 262338 117502 262574
rect 117586 262338 117822 262574
rect 117266 226658 117502 226894
rect 117586 226658 117822 226894
rect 117266 226338 117502 226574
rect 117586 226338 117822 226574
rect 117266 190658 117502 190894
rect 117586 190658 117822 190894
rect 117266 190338 117502 190574
rect 117586 190338 117822 190574
rect 117266 154658 117502 154894
rect 117586 154658 117822 154894
rect 117266 154338 117502 154574
rect 117586 154338 117822 154574
rect 117266 118658 117502 118894
rect 117586 118658 117822 118894
rect 117266 118338 117502 118574
rect 117586 118338 117822 118574
rect 117266 82658 117502 82894
rect 117586 82658 117822 82894
rect 117266 82338 117502 82574
rect 117586 82338 117822 82574
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 302378 121222 302614
rect 121306 302378 121542 302614
rect 120986 302058 121222 302294
rect 121306 302058 121542 302294
rect 120986 266378 121222 266614
rect 121306 266378 121542 266614
rect 120986 266058 121222 266294
rect 121306 266058 121542 266294
rect 120986 230378 121222 230614
rect 121306 230378 121542 230614
rect 120986 230058 121222 230294
rect 121306 230058 121542 230294
rect 120986 194378 121222 194614
rect 121306 194378 121542 194614
rect 120986 194058 121222 194294
rect 121306 194058 121542 194294
rect 120986 158378 121222 158614
rect 121306 158378 121542 158614
rect 120986 158058 121222 158294
rect 121306 158058 121542 158294
rect 120986 122378 121222 122614
rect 121306 122378 121542 122614
rect 120986 122058 121222 122294
rect 121306 122058 121542 122294
rect 120986 86378 121222 86614
rect 121306 86378 121542 86614
rect 120986 86058 121222 86294
rect 121306 86058 121542 86294
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 127826 165218 128062 165454
rect 128146 165218 128382 165454
rect 127826 164898 128062 165134
rect 128146 164898 128382 165134
rect 127826 129218 128062 129454
rect 128146 129218 128382 129454
rect 127826 128898 128062 129134
rect 128146 128898 128382 129134
rect 127826 93218 128062 93454
rect 128146 93218 128382 93454
rect 127826 92898 128062 93134
rect 128146 92898 128382 93134
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 131546 528938 131782 529174
rect 131866 528938 132102 529174
rect 131546 528618 131782 528854
rect 131866 528618 132102 528854
rect 131546 492938 131782 493174
rect 131866 492938 132102 493174
rect 131546 492618 131782 492854
rect 131866 492618 132102 492854
rect 131546 456938 131782 457174
rect 131866 456938 132102 457174
rect 131546 456618 131782 456854
rect 131866 456618 132102 456854
rect 131546 420938 131782 421174
rect 131866 420938 132102 421174
rect 131546 420618 131782 420854
rect 131866 420618 132102 420854
rect 131546 384938 131782 385174
rect 131866 384938 132102 385174
rect 131546 384618 131782 384854
rect 131866 384618 132102 384854
rect 131546 348938 131782 349174
rect 131866 348938 132102 349174
rect 131546 348618 131782 348854
rect 131866 348618 132102 348854
rect 131546 312938 131782 313174
rect 131866 312938 132102 313174
rect 131546 312618 131782 312854
rect 131866 312618 132102 312854
rect 131546 276938 131782 277174
rect 131866 276938 132102 277174
rect 131546 276618 131782 276854
rect 131866 276618 132102 276854
rect 131546 240938 131782 241174
rect 131866 240938 132102 241174
rect 131546 240618 131782 240854
rect 131866 240618 132102 240854
rect 131546 204938 131782 205174
rect 131866 204938 132102 205174
rect 131546 204618 131782 204854
rect 131866 204618 132102 204854
rect 131546 168938 131782 169174
rect 131866 168938 132102 169174
rect 131546 168618 131782 168854
rect 131866 168618 132102 168854
rect 131546 132938 131782 133174
rect 131866 132938 132102 133174
rect 131546 132618 131782 132854
rect 131866 132618 132102 132854
rect 131546 96938 131782 97174
rect 131866 96938 132102 97174
rect 131546 96618 131782 96854
rect 131866 96618 132102 96854
rect 131546 60938 131782 61174
rect 131866 60938 132102 61174
rect 131546 60618 131782 60854
rect 131866 60618 132102 60854
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 135266 532658 135502 532894
rect 135586 532658 135822 532894
rect 135266 532338 135502 532574
rect 135586 532338 135822 532574
rect 135266 496658 135502 496894
rect 135586 496658 135822 496894
rect 135266 496338 135502 496574
rect 135586 496338 135822 496574
rect 135266 460658 135502 460894
rect 135586 460658 135822 460894
rect 135266 460338 135502 460574
rect 135586 460338 135822 460574
rect 135266 424658 135502 424894
rect 135586 424658 135822 424894
rect 135266 424338 135502 424574
rect 135586 424338 135822 424574
rect 135266 388658 135502 388894
rect 135586 388658 135822 388894
rect 135266 388338 135502 388574
rect 135586 388338 135822 388574
rect 135266 352658 135502 352894
rect 135586 352658 135822 352894
rect 135266 352338 135502 352574
rect 135586 352338 135822 352574
rect 135266 316658 135502 316894
rect 135586 316658 135822 316894
rect 135266 316338 135502 316574
rect 135586 316338 135822 316574
rect 135266 280658 135502 280894
rect 135586 280658 135822 280894
rect 135266 280338 135502 280574
rect 135586 280338 135822 280574
rect 135266 244658 135502 244894
rect 135586 244658 135822 244894
rect 135266 244338 135502 244574
rect 135586 244338 135822 244574
rect 135266 208658 135502 208894
rect 135586 208658 135822 208894
rect 135266 208338 135502 208574
rect 135586 208338 135822 208574
rect 135266 172658 135502 172894
rect 135586 172658 135822 172894
rect 135266 172338 135502 172574
rect 135586 172338 135822 172574
rect 135266 136658 135502 136894
rect 135586 136658 135822 136894
rect 135266 136338 135502 136574
rect 135586 136338 135822 136574
rect 135266 100658 135502 100894
rect 135586 100658 135822 100894
rect 135266 100338 135502 100574
rect 135586 100338 135822 100574
rect 135266 64658 135502 64894
rect 135586 64658 135822 64894
rect 135266 64338 135502 64574
rect 135586 64338 135822 64574
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 138986 536378 139222 536614
rect 139306 536378 139542 536614
rect 138986 536058 139222 536294
rect 139306 536058 139542 536294
rect 138986 500378 139222 500614
rect 139306 500378 139542 500614
rect 138986 500058 139222 500294
rect 139306 500058 139542 500294
rect 138986 464378 139222 464614
rect 139306 464378 139542 464614
rect 138986 464058 139222 464294
rect 139306 464058 139542 464294
rect 138986 428378 139222 428614
rect 139306 428378 139542 428614
rect 138986 428058 139222 428294
rect 139306 428058 139542 428294
rect 138986 392378 139222 392614
rect 139306 392378 139542 392614
rect 138986 392058 139222 392294
rect 139306 392058 139542 392294
rect 138986 356378 139222 356614
rect 139306 356378 139542 356614
rect 138986 356058 139222 356294
rect 139306 356058 139542 356294
rect 138986 320378 139222 320614
rect 139306 320378 139542 320614
rect 138986 320058 139222 320294
rect 139306 320058 139542 320294
rect 138986 284378 139222 284614
rect 139306 284378 139542 284614
rect 138986 284058 139222 284294
rect 139306 284058 139542 284294
rect 138986 248378 139222 248614
rect 139306 248378 139542 248614
rect 138986 248058 139222 248294
rect 139306 248058 139542 248294
rect 138986 212378 139222 212614
rect 139306 212378 139542 212614
rect 138986 212058 139222 212294
rect 139306 212058 139542 212294
rect 138986 176378 139222 176614
rect 139306 176378 139542 176614
rect 138986 176058 139222 176294
rect 139306 176058 139542 176294
rect 138986 140378 139222 140614
rect 139306 140378 139542 140614
rect 138986 140058 139222 140294
rect 139306 140058 139542 140294
rect 138986 104378 139222 104614
rect 139306 104378 139542 104614
rect 138986 104058 139222 104294
rect 139306 104058 139542 104294
rect 138986 68378 139222 68614
rect 139306 68378 139542 68614
rect 138986 68058 139222 68294
rect 139306 68058 139542 68294
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 149546 438938 149782 439174
rect 149866 438938 150102 439174
rect 149546 438618 149782 438854
rect 149866 438618 150102 438854
rect 149546 402938 149782 403174
rect 149866 402938 150102 403174
rect 149546 402618 149782 402854
rect 149866 402618 150102 402854
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 149546 330938 149782 331174
rect 149866 330938 150102 331174
rect 149546 330618 149782 330854
rect 149866 330618 150102 330854
rect 149546 294938 149782 295174
rect 149866 294938 150102 295174
rect 149546 294618 149782 294854
rect 149866 294618 150102 294854
rect 149546 258938 149782 259174
rect 149866 258938 150102 259174
rect 149546 258618 149782 258854
rect 149866 258618 150102 258854
rect 149546 222938 149782 223174
rect 149866 222938 150102 223174
rect 149546 222618 149782 222854
rect 149866 222618 150102 222854
rect 149546 186938 149782 187174
rect 149866 186938 150102 187174
rect 149546 186618 149782 186854
rect 149866 186618 150102 186854
rect 149546 150938 149782 151174
rect 149866 150938 150102 151174
rect 149546 150618 149782 150854
rect 149866 150618 150102 150854
rect 149546 114938 149782 115174
rect 149866 114938 150102 115174
rect 149546 114618 149782 114854
rect 149866 114618 150102 114854
rect 149546 78938 149782 79174
rect 149866 78938 150102 79174
rect 149546 78618 149782 78854
rect 149866 78618 150102 78854
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 153266 514658 153502 514894
rect 153586 514658 153822 514894
rect 153266 514338 153502 514574
rect 153586 514338 153822 514574
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 153266 442658 153502 442894
rect 153586 442658 153822 442894
rect 153266 442338 153502 442574
rect 153586 442338 153822 442574
rect 153266 406658 153502 406894
rect 153586 406658 153822 406894
rect 153266 406338 153502 406574
rect 153586 406338 153822 406574
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 153266 334658 153502 334894
rect 153586 334658 153822 334894
rect 153266 334338 153502 334574
rect 153586 334338 153822 334574
rect 153266 298658 153502 298894
rect 153586 298658 153822 298894
rect 153266 298338 153502 298574
rect 153586 298338 153822 298574
rect 153266 262658 153502 262894
rect 153586 262658 153822 262894
rect 153266 262338 153502 262574
rect 153586 262338 153822 262574
rect 153266 226658 153502 226894
rect 153586 226658 153822 226894
rect 153266 226338 153502 226574
rect 153586 226338 153822 226574
rect 153266 190658 153502 190894
rect 153586 190658 153822 190894
rect 153266 190338 153502 190574
rect 153586 190338 153822 190574
rect 153266 154658 153502 154894
rect 153586 154658 153822 154894
rect 153266 154338 153502 154574
rect 153586 154338 153822 154574
rect 153266 118658 153502 118894
rect 153586 118658 153822 118894
rect 153266 118338 153502 118574
rect 153586 118338 153822 118574
rect 153266 82658 153502 82894
rect 153586 82658 153822 82894
rect 153266 82338 153502 82574
rect 153586 82338 153822 82574
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 156986 518378 157222 518614
rect 157306 518378 157542 518614
rect 156986 518058 157222 518294
rect 157306 518058 157542 518294
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 156986 446378 157222 446614
rect 157306 446378 157542 446614
rect 156986 446058 157222 446294
rect 157306 446058 157542 446294
rect 156986 410378 157222 410614
rect 157306 410378 157542 410614
rect 156986 410058 157222 410294
rect 157306 410058 157542 410294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 156986 374378 157222 374614
rect 157306 374378 157542 374614
rect 156986 374058 157222 374294
rect 157306 374058 157542 374294
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 156986 338378 157222 338614
rect 157306 338378 157542 338614
rect 156986 338058 157222 338294
rect 157306 338058 157542 338294
rect 156986 302378 157222 302614
rect 157306 302378 157542 302614
rect 156986 302058 157222 302294
rect 157306 302058 157542 302294
rect 156986 266378 157222 266614
rect 157306 266378 157542 266614
rect 156986 266058 157222 266294
rect 157306 266058 157542 266294
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 156986 230378 157222 230614
rect 157306 230378 157542 230614
rect 156986 230058 157222 230294
rect 157306 230058 157542 230294
rect 156986 194378 157222 194614
rect 157306 194378 157542 194614
rect 156986 194058 157222 194294
rect 157306 194058 157542 194294
rect 156986 158378 157222 158614
rect 157306 158378 157542 158614
rect 156986 158058 157222 158294
rect 157306 158058 157542 158294
rect 156986 122378 157222 122614
rect 157306 122378 157542 122614
rect 156986 122058 157222 122294
rect 157306 122058 157542 122294
rect 156986 86378 157222 86614
rect 157306 86378 157542 86614
rect 156986 86058 157222 86294
rect 157306 86058 157542 86294
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 163826 165218 164062 165454
rect 164146 165218 164382 165454
rect 163826 164898 164062 165134
rect 164146 164898 164382 165134
rect 163826 129218 164062 129454
rect 164146 129218 164382 129454
rect 163826 128898 164062 129134
rect 164146 128898 164382 129134
rect 163826 93218 164062 93454
rect 164146 93218 164382 93454
rect 163826 92898 164062 93134
rect 164146 92898 164382 93134
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 167546 528938 167782 529174
rect 167866 528938 168102 529174
rect 167546 528618 167782 528854
rect 167866 528618 168102 528854
rect 167546 492938 167782 493174
rect 167866 492938 168102 493174
rect 167546 492618 167782 492854
rect 167866 492618 168102 492854
rect 167546 456938 167782 457174
rect 167866 456938 168102 457174
rect 167546 456618 167782 456854
rect 167866 456618 168102 456854
rect 167546 420938 167782 421174
rect 167866 420938 168102 421174
rect 167546 420618 167782 420854
rect 167866 420618 168102 420854
rect 167546 384938 167782 385174
rect 167866 384938 168102 385174
rect 167546 384618 167782 384854
rect 167866 384618 168102 384854
rect 167546 348938 167782 349174
rect 167866 348938 168102 349174
rect 167546 348618 167782 348854
rect 167866 348618 168102 348854
rect 167546 312938 167782 313174
rect 167866 312938 168102 313174
rect 167546 312618 167782 312854
rect 167866 312618 168102 312854
rect 167546 276938 167782 277174
rect 167866 276938 168102 277174
rect 167546 276618 167782 276854
rect 167866 276618 168102 276854
rect 167546 240938 167782 241174
rect 167866 240938 168102 241174
rect 167546 240618 167782 240854
rect 167866 240618 168102 240854
rect 167546 204938 167782 205174
rect 167866 204938 168102 205174
rect 167546 204618 167782 204854
rect 167866 204618 168102 204854
rect 167546 168938 167782 169174
rect 167866 168938 168102 169174
rect 167546 168618 167782 168854
rect 167866 168618 168102 168854
rect 167546 132938 167782 133174
rect 167866 132938 168102 133174
rect 167546 132618 167782 132854
rect 167866 132618 168102 132854
rect 167546 96938 167782 97174
rect 167866 96938 168102 97174
rect 167546 96618 167782 96854
rect 167866 96618 168102 96854
rect 167546 60938 167782 61174
rect 167866 60938 168102 61174
rect 167546 60618 167782 60854
rect 167866 60618 168102 60854
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 171266 532658 171502 532894
rect 171586 532658 171822 532894
rect 171266 532338 171502 532574
rect 171586 532338 171822 532574
rect 171266 496658 171502 496894
rect 171586 496658 171822 496894
rect 171266 496338 171502 496574
rect 171586 496338 171822 496574
rect 171266 460658 171502 460894
rect 171586 460658 171822 460894
rect 171266 460338 171502 460574
rect 171586 460338 171822 460574
rect 171266 424658 171502 424894
rect 171586 424658 171822 424894
rect 171266 424338 171502 424574
rect 171586 424338 171822 424574
rect 171266 388658 171502 388894
rect 171586 388658 171822 388894
rect 171266 388338 171502 388574
rect 171586 388338 171822 388574
rect 171266 352658 171502 352894
rect 171586 352658 171822 352894
rect 171266 352338 171502 352574
rect 171586 352338 171822 352574
rect 171266 316658 171502 316894
rect 171586 316658 171822 316894
rect 171266 316338 171502 316574
rect 171586 316338 171822 316574
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 174986 536378 175222 536614
rect 175306 536378 175542 536614
rect 174986 536058 175222 536294
rect 175306 536058 175542 536294
rect 174986 500378 175222 500614
rect 175306 500378 175542 500614
rect 174986 500058 175222 500294
rect 175306 500058 175542 500294
rect 174986 464378 175222 464614
rect 175306 464378 175542 464614
rect 174986 464058 175222 464294
rect 175306 464058 175542 464294
rect 174986 428378 175222 428614
rect 175306 428378 175542 428614
rect 174986 428058 175222 428294
rect 175306 428058 175542 428294
rect 174986 392378 175222 392614
rect 175306 392378 175542 392614
rect 174986 392058 175222 392294
rect 175306 392058 175542 392294
rect 174986 356378 175222 356614
rect 175306 356378 175542 356614
rect 174986 356058 175222 356294
rect 175306 356058 175542 356294
rect 174986 320378 175222 320614
rect 175306 320378 175542 320614
rect 174986 320058 175222 320294
rect 175306 320058 175542 320294
rect 171266 280658 171502 280894
rect 171586 280658 171822 280894
rect 171266 280338 171502 280574
rect 171586 280338 171822 280574
rect 174986 284378 175222 284614
rect 175306 284378 175542 284614
rect 174986 284058 175222 284294
rect 175306 284058 175542 284294
rect 171266 244658 171502 244894
rect 171586 244658 171822 244894
rect 171266 244338 171502 244574
rect 171586 244338 171822 244574
rect 171266 208658 171502 208894
rect 171586 208658 171822 208894
rect 171266 208338 171502 208574
rect 171586 208338 171822 208574
rect 171266 172658 171502 172894
rect 171586 172658 171822 172894
rect 171266 172338 171502 172574
rect 171586 172338 171822 172574
rect 171266 136658 171502 136894
rect 171586 136658 171822 136894
rect 171266 136338 171502 136574
rect 171586 136338 171822 136574
rect 171266 100658 171502 100894
rect 171586 100658 171822 100894
rect 171266 100338 171502 100574
rect 171586 100338 171822 100574
rect 171266 64658 171502 64894
rect 171586 64658 171822 64894
rect 171266 64338 171502 64574
rect 171586 64338 171822 64574
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 185546 438938 185782 439174
rect 185866 438938 186102 439174
rect 185546 438618 185782 438854
rect 185866 438618 186102 438854
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 192986 518378 193222 518614
rect 193306 518378 193542 518614
rect 192986 518058 193222 518294
rect 193306 518058 193542 518294
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 189266 442658 189502 442894
rect 189586 442658 189822 442894
rect 189266 442338 189502 442574
rect 189586 442338 189822 442574
rect 185546 402938 185782 403174
rect 185866 402938 186102 403174
rect 185546 402618 185782 402854
rect 185866 402618 186102 402854
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 189266 406658 189502 406894
rect 189586 406658 189822 406894
rect 189266 406338 189502 406574
rect 189586 406338 189822 406574
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 185546 330938 185782 331174
rect 185866 330938 186102 331174
rect 185546 330618 185782 330854
rect 185866 330618 186102 330854
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 189266 334658 189502 334894
rect 189586 334658 189822 334894
rect 189266 334338 189502 334574
rect 189586 334338 189822 334574
rect 185546 294938 185782 295174
rect 185866 294938 186102 295174
rect 185546 294618 185782 294854
rect 185866 294618 186102 294854
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 174986 248378 175222 248614
rect 175306 248378 175542 248614
rect 174986 248058 175222 248294
rect 175306 248058 175542 248294
rect 174986 212378 175222 212614
rect 175306 212378 175542 212614
rect 174986 212058 175222 212294
rect 175306 212058 175542 212294
rect 174986 176378 175222 176614
rect 175306 176378 175542 176614
rect 174986 176058 175222 176294
rect 175306 176058 175542 176294
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 174986 140378 175222 140614
rect 175306 140378 175542 140614
rect 174986 140058 175222 140294
rect 175306 140058 175542 140294
rect 174986 104378 175222 104614
rect 175306 104378 175542 104614
rect 174986 104058 175222 104294
rect 175306 104058 175542 104294
rect 174986 68378 175222 68614
rect 175306 68378 175542 68614
rect 174986 68058 175222 68294
rect 175306 68058 175542 68294
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 185546 222938 185782 223174
rect 185866 222938 186102 223174
rect 185546 222618 185782 222854
rect 185866 222618 186102 222854
rect 192986 374378 193222 374614
rect 193306 374378 193542 374614
rect 192986 374058 193222 374294
rect 193306 374058 193542 374294
rect 192986 338378 193222 338614
rect 193306 338378 193542 338614
rect 192986 338058 193222 338294
rect 193306 338058 193542 338294
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 203546 528938 203782 529174
rect 203866 528938 204102 529174
rect 203546 528618 203782 528854
rect 203866 528618 204102 528854
rect 203546 492938 203782 493174
rect 203866 492938 204102 493174
rect 203546 492618 203782 492854
rect 203866 492618 204102 492854
rect 203546 456938 203782 457174
rect 203866 456938 204102 457174
rect 203546 456618 203782 456854
rect 203866 456618 204102 456854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 207266 532658 207502 532894
rect 207586 532658 207822 532894
rect 207266 532338 207502 532574
rect 207586 532338 207822 532574
rect 207266 496658 207502 496894
rect 207586 496658 207822 496894
rect 207266 496338 207502 496574
rect 207586 496338 207822 496574
rect 207266 460658 207502 460894
rect 207586 460658 207822 460894
rect 207266 460338 207502 460574
rect 207586 460338 207822 460574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 210986 536378 211222 536614
rect 211306 536378 211542 536614
rect 210986 536058 211222 536294
rect 211306 536058 211542 536294
rect 210986 500378 211222 500614
rect 211306 500378 211542 500614
rect 210986 500058 211222 500294
rect 211306 500058 211542 500294
rect 210986 464378 211222 464614
rect 211306 464378 211542 464614
rect 210986 464058 211222 464294
rect 211306 464058 211542 464294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 221546 510938 221782 511174
rect 221866 510938 222102 511174
rect 221546 510618 221782 510854
rect 221866 510618 222102 510854
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 225266 514658 225502 514894
rect 225586 514658 225822 514894
rect 225266 514338 225502 514574
rect 225586 514338 225822 514574
rect 225266 478658 225502 478894
rect 225586 478658 225822 478894
rect 225266 478338 225502 478574
rect 225586 478338 225822 478574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 228986 518378 229222 518614
rect 229306 518378 229542 518614
rect 228986 518058 229222 518294
rect 229306 518058 229542 518294
rect 228986 482378 229222 482614
rect 229306 482378 229542 482614
rect 228986 482058 229222 482294
rect 229306 482058 229542 482294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 239546 600938 239782 601174
rect 239866 600938 240102 601174
rect 239546 600618 239782 600854
rect 239866 600618 240102 600854
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 239546 528938 239782 529174
rect 239866 528938 240102 529174
rect 239546 528618 239782 528854
rect 239866 528618 240102 528854
rect 239546 492938 239782 493174
rect 239866 492938 240102 493174
rect 239546 492618 239782 492854
rect 239866 492618 240102 492854
rect 239546 456938 239782 457174
rect 239866 456938 240102 457174
rect 239546 456618 239782 456854
rect 239866 456618 240102 456854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 243266 604658 243502 604894
rect 243586 604658 243822 604894
rect 243266 604338 243502 604574
rect 243586 604338 243822 604574
rect 243266 568658 243502 568894
rect 243586 568658 243822 568894
rect 243266 568338 243502 568574
rect 243586 568338 243822 568574
rect 243266 532658 243502 532894
rect 243586 532658 243822 532894
rect 243266 532338 243502 532574
rect 243586 532338 243822 532574
rect 243266 496658 243502 496894
rect 243586 496658 243822 496894
rect 243266 496338 243502 496574
rect 243586 496338 243822 496574
rect 243266 460658 243502 460894
rect 243586 460658 243822 460894
rect 243266 460338 243502 460574
rect 243586 460338 243822 460574
rect 197818 435218 198054 435454
rect 197818 434898 198054 435134
rect 228538 435218 228774 435454
rect 228538 434898 228774 435134
rect 213178 417218 213414 417454
rect 213178 416898 213414 417134
rect 197818 399218 198054 399454
rect 197818 398898 198054 399134
rect 228538 399218 228774 399454
rect 228538 398898 228774 399134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 189266 298658 189502 298894
rect 189586 298658 189822 298894
rect 189266 298338 189502 298574
rect 189586 298338 189822 298574
rect 185546 186938 185782 187174
rect 185866 186938 186102 187174
rect 185546 186618 185782 186854
rect 185866 186618 186102 186854
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 185546 114938 185782 115174
rect 185866 114938 186102 115174
rect 185546 114618 185782 114854
rect 185866 114618 186102 114854
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 189266 262658 189502 262894
rect 189586 262658 189822 262894
rect 189266 262338 189502 262574
rect 189586 262338 189822 262574
rect 189266 226658 189502 226894
rect 189586 226658 189822 226894
rect 189266 226338 189502 226574
rect 189586 226338 189822 226574
rect 189266 190658 189502 190894
rect 189586 190658 189822 190894
rect 189266 190338 189502 190574
rect 189586 190338 189822 190574
rect 189266 154658 189502 154894
rect 189586 154658 189822 154894
rect 189266 154338 189502 154574
rect 189586 154338 189822 154574
rect 189266 118658 189502 118894
rect 189586 118658 189822 118894
rect 189266 118338 189502 118574
rect 189586 118338 189822 118574
rect 185546 78938 185782 79174
rect 185866 78938 186102 79174
rect 185546 78618 185782 78854
rect 185866 78618 186102 78854
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 197818 291218 198054 291454
rect 197818 290898 198054 291134
rect 192986 230378 193222 230614
rect 193306 230378 193542 230614
rect 192986 230058 193222 230294
rect 193306 230058 193542 230294
rect 192986 194378 193222 194614
rect 193306 194378 193542 194614
rect 192986 194058 193222 194294
rect 193306 194058 193542 194294
rect 192986 158378 193222 158614
rect 193306 158378 193542 158614
rect 192986 158058 193222 158294
rect 193306 158058 193542 158294
rect 197818 255218 198054 255454
rect 197818 254898 198054 255134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 203546 384938 203782 385174
rect 203866 384938 204102 385174
rect 203546 384618 203782 384854
rect 203866 384618 204102 384854
rect 203546 348938 203782 349174
rect 203866 348938 204102 349174
rect 203546 348618 203782 348854
rect 203866 348618 204102 348854
rect 203546 312938 203782 313174
rect 203866 312938 204102 313174
rect 203546 312618 203782 312854
rect 203866 312618 204102 312854
rect 207266 352658 207502 352894
rect 207586 352658 207822 352894
rect 207266 352338 207502 352574
rect 207586 352338 207822 352574
rect 207266 316658 207502 316894
rect 207586 316658 207822 316894
rect 207266 316338 207502 316574
rect 207586 316338 207822 316574
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 189266 82658 189502 82894
rect 189586 82658 189822 82894
rect 189266 82338 189502 82574
rect 189586 82338 189822 82574
rect 192986 86378 193222 86614
rect 193306 86378 193542 86614
rect 192986 86058 193222 86294
rect 193306 86058 193542 86294
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199430 111218 199666 111454
rect 199430 110898 199666 111134
rect 203546 204938 203782 205174
rect 203866 204938 204102 205174
rect 203546 204618 203782 204854
rect 203866 204618 204102 204854
rect 203546 168938 203782 169174
rect 203866 168938 204102 169174
rect 203546 168618 203782 168854
rect 203866 168618 204102 168854
rect 204306 129218 204542 129454
rect 204306 128898 204542 129134
rect 210986 356378 211222 356614
rect 211306 356378 211542 356614
rect 210986 356058 211222 356294
rect 211306 356058 211542 356294
rect 210986 320378 211222 320614
rect 211306 320378 211542 320614
rect 210986 320058 211222 320294
rect 211306 320058 211542 320294
rect 207266 208658 207502 208894
rect 207586 208658 207822 208894
rect 207266 208338 207502 208574
rect 207586 208338 207822 208574
rect 207266 172658 207502 172894
rect 207586 172658 207822 172894
rect 207266 172338 207502 172574
rect 207586 172338 207822 172574
rect 209182 111218 209418 111454
rect 209182 110898 209418 111134
rect 213178 273218 213414 273454
rect 213178 272898 213414 273134
rect 210986 212378 211222 212614
rect 211306 212378 211542 212614
rect 210986 212058 211222 212294
rect 211306 212058 211542 212294
rect 210986 176378 211222 176614
rect 211306 176378 211542 176614
rect 210986 176058 211222 176294
rect 211306 176058 211542 176294
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 60938 203782 61174
rect 203866 60938 204102 61174
rect 203546 60618 203782 60854
rect 203866 60618 204102 60854
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 221546 366938 221782 367174
rect 221866 366938 222102 367174
rect 221546 366618 221782 366854
rect 221866 366618 222102 366854
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 214058 129218 214294 129454
rect 214058 128898 214294 129134
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 218934 111218 219170 111454
rect 218934 110898 219170 111134
rect 221546 330938 221782 331174
rect 221866 330938 222102 331174
rect 221546 330618 221782 330854
rect 221866 330618 222102 330854
rect 225266 370658 225502 370894
rect 225586 370658 225822 370894
rect 225266 370338 225502 370574
rect 225586 370338 225822 370574
rect 225266 334658 225502 334894
rect 225586 334658 225822 334894
rect 225266 334338 225502 334574
rect 225586 334338 225822 334574
rect 221546 222938 221782 223174
rect 221866 222938 222102 223174
rect 221546 222618 221782 222854
rect 221866 222618 222102 222854
rect 221546 186938 221782 187174
rect 221866 186938 222102 187174
rect 221546 186618 221782 186854
rect 221866 186618 222102 186854
rect 221546 150938 221782 151174
rect 221866 150938 222102 151174
rect 221546 150618 221782 150854
rect 221866 150618 222102 150854
rect 228986 374378 229222 374614
rect 229306 374378 229542 374614
rect 228986 374058 229222 374294
rect 229306 374058 229542 374294
rect 228986 338378 229222 338614
rect 229306 338378 229542 338614
rect 228986 338058 229222 338294
rect 229306 338058 229542 338294
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 239546 384938 239782 385174
rect 239866 384938 240102 385174
rect 239546 384618 239782 384854
rect 239866 384618 240102 384854
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 225266 226658 225502 226894
rect 225586 226658 225822 226894
rect 225266 226338 225502 226574
rect 225586 226338 225822 226574
rect 225266 190658 225502 190894
rect 225586 190658 225822 190894
rect 225266 190338 225502 190574
rect 225586 190338 225822 190574
rect 228538 291218 228774 291454
rect 228538 290898 228774 291134
rect 228538 255218 228774 255454
rect 228538 254898 228774 255134
rect 228986 230378 229222 230614
rect 229306 230378 229542 230614
rect 228986 230058 229222 230294
rect 229306 230058 229542 230294
rect 228986 194378 229222 194614
rect 229306 194378 229542 194614
rect 228986 194058 229222 194294
rect 229306 194058 229542 194294
rect 225266 154658 225502 154894
rect 225586 154658 225822 154894
rect 225266 154338 225502 154574
rect 225586 154338 225822 154574
rect 228986 158378 229222 158614
rect 229306 158378 229542 158614
rect 228986 158058 229222 158294
rect 229306 158058 229542 158294
rect 228986 122378 229222 122614
rect 229306 122378 229542 122614
rect 228986 122058 229222 122294
rect 229306 122058 229542 122294
rect 207266 64658 207502 64894
rect 207586 64658 207822 64894
rect 207266 64338 207502 64574
rect 207586 64338 207822 64574
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 210986 68378 211222 68614
rect 211306 68378 211542 68614
rect 210986 68058 211222 68294
rect 211306 68058 211542 68294
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 78938 221782 79174
rect 221866 78938 222102 79174
rect 221546 78618 221782 78854
rect 221866 78618 222102 78854
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 82658 225502 82894
rect 225586 82658 225822 82894
rect 228986 86378 229222 86614
rect 229306 86378 229542 86614
rect 228986 86058 229222 86294
rect 229306 86058 229542 86294
rect 225266 82338 225502 82574
rect 225586 82338 225822 82574
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 239546 348938 239782 349174
rect 239866 348938 240102 349174
rect 239546 348618 239782 348854
rect 239866 348618 240102 348854
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 239546 312938 239782 313174
rect 239866 312938 240102 313174
rect 239546 312618 239782 312854
rect 239866 312618 240102 312854
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 246986 608378 247222 608614
rect 247306 608378 247542 608614
rect 246986 608058 247222 608294
rect 247306 608058 247542 608294
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 246986 536378 247222 536614
rect 247306 536378 247542 536614
rect 246986 536058 247222 536294
rect 247306 536058 247542 536294
rect 246986 500378 247222 500614
rect 247306 500378 247542 500614
rect 246986 500058 247222 500294
rect 247306 500058 247542 500294
rect 246986 464378 247222 464614
rect 247306 464378 247542 464614
rect 246986 464058 247222 464294
rect 247306 464058 247542 464294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 243898 417218 244134 417454
rect 243898 416898 244134 417134
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 243266 352658 243502 352894
rect 243586 352658 243822 352894
rect 243266 352338 243502 352574
rect 243586 352338 243822 352574
rect 243266 316658 243502 316894
rect 243586 316658 243822 316894
rect 243266 316338 243502 316574
rect 243586 316338 243822 316574
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 257546 510938 257782 511174
rect 257866 510938 258102 511174
rect 257546 510618 257782 510854
rect 257866 510618 258102 510854
rect 257546 474938 257782 475174
rect 257866 474938 258102 475174
rect 257546 474618 257782 474854
rect 257866 474618 258102 474854
rect 246986 356378 247222 356614
rect 247306 356378 247542 356614
rect 246986 356058 247222 356294
rect 247306 356058 247542 356294
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 246986 320378 247222 320614
rect 247306 320378 247542 320614
rect 246986 320058 247222 320294
rect 247306 320058 247542 320294
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 261266 514658 261502 514894
rect 261586 514658 261822 514894
rect 261266 514338 261502 514574
rect 261586 514338 261822 514574
rect 261266 478658 261502 478894
rect 261586 478658 261822 478894
rect 261266 478338 261502 478574
rect 261586 478338 261822 478574
rect 261266 442658 261502 442894
rect 261586 442658 261822 442894
rect 261266 442338 261502 442574
rect 261586 442338 261822 442574
rect 257546 438938 257782 439174
rect 257866 438938 258102 439174
rect 257546 438618 257782 438854
rect 257866 438618 258102 438854
rect 257546 402938 257782 403174
rect 257866 402938 258102 403174
rect 257546 402618 257782 402854
rect 257866 402618 258102 402854
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 264986 518378 265222 518614
rect 265306 518378 265542 518614
rect 264986 518058 265222 518294
rect 265306 518058 265542 518294
rect 264986 482378 265222 482614
rect 265306 482378 265542 482614
rect 264986 482058 265222 482294
rect 265306 482058 265542 482294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 264986 446378 265222 446614
rect 265306 446378 265542 446614
rect 264986 446058 265222 446294
rect 265306 446058 265542 446294
rect 261266 406658 261502 406894
rect 261586 406658 261822 406894
rect 261266 406338 261502 406574
rect 261586 406338 261822 406574
rect 257546 366938 257782 367174
rect 257866 366938 258102 367174
rect 257546 366618 257782 366854
rect 257866 366618 258102 366854
rect 257546 330938 257782 331174
rect 257866 330938 258102 331174
rect 257546 330618 257782 330854
rect 257866 330618 258102 330854
rect 239546 204938 239782 205174
rect 239866 204938 240102 205174
rect 239546 204618 239782 204854
rect 239866 204618 240102 204854
rect 243898 273218 244134 273454
rect 243898 272898 244134 273134
rect 243266 208658 243502 208894
rect 243586 208658 243822 208894
rect 243266 208338 243502 208574
rect 243586 208338 243822 208574
rect 239546 168938 239782 169174
rect 239866 168938 240102 169174
rect 239546 168618 239782 168854
rect 239866 168618 240102 168854
rect 239546 132938 239782 133174
rect 239866 132938 240102 133174
rect 239546 132618 239782 132854
rect 239866 132618 240102 132854
rect 239546 96938 239782 97174
rect 239866 96938 240102 97174
rect 239546 96618 239782 96854
rect 239866 96618 240102 96854
rect 239546 60938 239782 61174
rect 239866 60938 240102 61174
rect 239546 60618 239782 60854
rect 239866 60618 240102 60854
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 172658 243502 172894
rect 243586 172658 243822 172894
rect 243266 172338 243502 172574
rect 243586 172338 243822 172574
rect 243266 136658 243502 136894
rect 243586 136658 243822 136894
rect 243266 136338 243502 136574
rect 243586 136338 243822 136574
rect 243266 100658 243502 100894
rect 243586 100658 243822 100894
rect 243266 100338 243502 100574
rect 243586 100338 243822 100574
rect 243266 64658 243502 64894
rect 243586 64658 243822 64894
rect 243266 64338 243502 64574
rect 243586 64338 243822 64574
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 246986 212378 247222 212614
rect 247306 212378 247542 212614
rect 246986 212058 247222 212294
rect 247306 212058 247542 212294
rect 246986 176378 247222 176614
rect 247306 176378 247542 176614
rect 246986 176058 247222 176294
rect 247306 176058 247542 176294
rect 246986 140378 247222 140614
rect 247306 140378 247542 140614
rect 246986 140058 247222 140294
rect 247306 140058 247542 140294
rect 246986 104378 247222 104614
rect 247306 104378 247542 104614
rect 246986 104058 247222 104294
rect 247306 104058 247542 104294
rect 246986 68378 247222 68614
rect 247306 68378 247542 68614
rect 246986 68058 247222 68294
rect 247306 68058 247542 68294
rect 261266 370658 261502 370894
rect 261586 370658 261822 370894
rect 261266 370338 261502 370574
rect 261586 370338 261822 370574
rect 261266 334658 261502 334894
rect 261586 334658 261822 334894
rect 261266 334338 261502 334574
rect 261586 334338 261822 334574
rect 257546 294938 257782 295174
rect 257866 294938 258102 295174
rect 257546 294618 257782 294854
rect 257866 294618 258102 294854
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 257546 258938 257782 259174
rect 257866 258938 258102 259174
rect 257546 258618 257782 258854
rect 257866 258618 258102 258854
rect 257546 222938 257782 223174
rect 257866 222938 258102 223174
rect 257546 222618 257782 222854
rect 257866 222618 258102 222854
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 261266 298658 261502 298894
rect 261586 298658 261822 298894
rect 261266 298338 261502 298574
rect 261586 298338 261822 298574
rect 261266 262658 261502 262894
rect 261586 262658 261822 262894
rect 261266 262338 261502 262574
rect 261586 262338 261822 262574
rect 264986 410378 265222 410614
rect 265306 410378 265542 410614
rect 264986 410058 265222 410294
rect 265306 410058 265542 410294
rect 264986 374378 265222 374614
rect 265306 374378 265542 374614
rect 264986 374058 265222 374294
rect 265306 374058 265542 374294
rect 264986 338378 265222 338614
rect 265306 338378 265542 338614
rect 264986 338058 265222 338294
rect 265306 338058 265542 338294
rect 261266 226658 261502 226894
rect 261586 226658 261822 226894
rect 261266 226338 261502 226574
rect 261586 226338 261822 226574
rect 257546 186938 257782 187174
rect 257866 186938 258102 187174
rect 257546 186618 257782 186854
rect 257866 186618 258102 186854
rect 264986 302378 265222 302614
rect 265306 302378 265542 302614
rect 264986 302058 265222 302294
rect 265306 302058 265542 302294
rect 264986 266378 265222 266614
rect 265306 266378 265542 266614
rect 264986 266058 265222 266294
rect 265306 266058 265542 266294
rect 264986 230378 265222 230614
rect 265306 230378 265542 230614
rect 264986 230058 265222 230294
rect 265306 230058 265542 230294
rect 261266 190658 261502 190894
rect 261586 190658 261822 190894
rect 261266 190338 261502 190574
rect 261586 190338 261822 190574
rect 257546 150938 257782 151174
rect 257866 150938 258102 151174
rect 257546 150618 257782 150854
rect 257866 150618 258102 150854
rect 257546 114938 257782 115174
rect 257866 114938 258102 115174
rect 257546 114618 257782 114854
rect 257866 114618 258102 114854
rect 257546 78938 257782 79174
rect 257866 78938 258102 79174
rect 257546 78618 257782 78854
rect 257866 78618 258102 78854
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 154658 261502 154894
rect 261586 154658 261822 154894
rect 261266 154338 261502 154574
rect 261586 154338 261822 154574
rect 261266 118658 261502 118894
rect 261586 118658 261822 118894
rect 261266 118338 261502 118574
rect 261586 118338 261822 118574
rect 261266 82658 261502 82894
rect 261586 82658 261822 82894
rect 261266 82338 261502 82574
rect 261586 82338 261822 82574
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 275546 600938 275782 601174
rect 275866 600938 276102 601174
rect 275546 600618 275782 600854
rect 275866 600618 276102 600854
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 275546 528938 275782 529174
rect 275866 528938 276102 529174
rect 275546 528618 275782 528854
rect 275866 528618 276102 528854
rect 275546 492938 275782 493174
rect 275866 492938 276102 493174
rect 275546 492618 275782 492854
rect 275866 492618 276102 492854
rect 275546 456938 275782 457174
rect 275866 456938 276102 457174
rect 275546 456618 275782 456854
rect 275866 456618 276102 456854
rect 275546 420938 275782 421174
rect 275866 420938 276102 421174
rect 275546 420618 275782 420854
rect 275866 420618 276102 420854
rect 275546 384938 275782 385174
rect 275866 384938 276102 385174
rect 275546 384618 275782 384854
rect 275866 384618 276102 384854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 279266 604658 279502 604894
rect 279586 604658 279822 604894
rect 279266 604338 279502 604574
rect 279586 604338 279822 604574
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 279266 532658 279502 532894
rect 279586 532658 279822 532894
rect 279266 532338 279502 532574
rect 279586 532338 279822 532574
rect 279266 496658 279502 496894
rect 279586 496658 279822 496894
rect 279266 496338 279502 496574
rect 279586 496338 279822 496574
rect 279266 460658 279502 460894
rect 279586 460658 279822 460894
rect 279266 460338 279502 460574
rect 279586 460338 279822 460574
rect 279266 424658 279502 424894
rect 279586 424658 279822 424894
rect 279266 424338 279502 424574
rect 279586 424338 279822 424574
rect 279266 388658 279502 388894
rect 279586 388658 279822 388894
rect 279266 388338 279502 388574
rect 279586 388338 279822 388574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 282986 608378 283222 608614
rect 283306 608378 283542 608614
rect 282986 608058 283222 608294
rect 283306 608058 283542 608294
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 282986 536378 283222 536614
rect 283306 536378 283542 536614
rect 282986 536058 283222 536294
rect 283306 536058 283542 536294
rect 282986 500378 283222 500614
rect 283306 500378 283542 500614
rect 282986 500058 283222 500294
rect 283306 500058 283542 500294
rect 282986 464378 283222 464614
rect 283306 464378 283542 464614
rect 282986 464058 283222 464294
rect 283306 464058 283542 464294
rect 282986 428378 283222 428614
rect 283306 428378 283542 428614
rect 282986 428058 283222 428294
rect 283306 428058 283542 428294
rect 282986 392378 283222 392614
rect 283306 392378 283542 392614
rect 282986 392058 283222 392294
rect 283306 392058 283542 392294
rect 275546 348938 275782 349174
rect 275866 348938 276102 349174
rect 275546 348618 275782 348854
rect 275866 348618 276102 348854
rect 275546 312938 275782 313174
rect 275866 312938 276102 313174
rect 275546 312618 275782 312854
rect 275866 312618 276102 312854
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 264986 194378 265222 194614
rect 265306 194378 265542 194614
rect 264986 194058 265222 194294
rect 265306 194058 265542 194294
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 264986 158378 265222 158614
rect 265306 158378 265542 158614
rect 264986 158058 265222 158294
rect 265306 158058 265542 158294
rect 264986 122378 265222 122614
rect 265306 122378 265542 122614
rect 264986 122058 265222 122294
rect 265306 122058 265542 122294
rect 264986 86378 265222 86614
rect 265306 86378 265542 86614
rect 264986 86058 265222 86294
rect 265306 86058 265542 86294
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 275546 276938 275782 277174
rect 275866 276938 276102 277174
rect 275546 276618 275782 276854
rect 275866 276618 276102 276854
rect 279266 352658 279502 352894
rect 279586 352658 279822 352894
rect 279266 352338 279502 352574
rect 279586 352338 279822 352574
rect 279266 316658 279502 316894
rect 279586 316658 279822 316894
rect 279266 316338 279502 316574
rect 279586 316338 279822 316574
rect 275546 240938 275782 241174
rect 275866 240938 276102 241174
rect 275546 240618 275782 240854
rect 275866 240618 276102 240854
rect 279266 280658 279502 280894
rect 279586 280658 279822 280894
rect 279266 280338 279502 280574
rect 279586 280338 279822 280574
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 282986 356378 283222 356614
rect 283306 356378 283542 356614
rect 282986 356058 283222 356294
rect 283306 356058 283542 356294
rect 282986 320378 283222 320614
rect 283306 320378 283542 320614
rect 282986 320058 283222 320294
rect 283306 320058 283542 320294
rect 282986 284378 283222 284614
rect 283306 284378 283542 284614
rect 282986 284058 283222 284294
rect 283306 284058 283542 284294
rect 279266 244658 279502 244894
rect 279586 244658 279822 244894
rect 279266 244338 279502 244574
rect 279586 244338 279822 244574
rect 275546 204938 275782 205174
rect 275866 204938 276102 205174
rect 275546 204618 275782 204854
rect 275866 204618 276102 204854
rect 275546 168938 275782 169174
rect 275866 168938 276102 169174
rect 275546 168618 275782 168854
rect 275866 168618 276102 168854
rect 275546 132938 275782 133174
rect 275866 132938 276102 133174
rect 275546 132618 275782 132854
rect 275866 132618 276102 132854
rect 275546 96938 275782 97174
rect 275866 96938 276102 97174
rect 275546 96618 275782 96854
rect 275866 96618 276102 96854
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 60938 275782 61174
rect 275866 60938 276102 61174
rect 275546 60618 275782 60854
rect 275866 60618 276102 60854
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 208658 279502 208894
rect 279586 208658 279822 208894
rect 279266 208338 279502 208574
rect 279586 208338 279822 208574
rect 279266 172658 279502 172894
rect 279586 172658 279822 172894
rect 279266 172338 279502 172574
rect 279586 172338 279822 172574
rect 279266 136658 279502 136894
rect 279586 136658 279822 136894
rect 279266 136338 279502 136574
rect 279586 136338 279822 136574
rect 279266 100658 279502 100894
rect 279586 100658 279822 100894
rect 279266 100338 279502 100574
rect 279586 100338 279822 100574
rect 279266 64658 279502 64894
rect 279586 64658 279822 64894
rect 279266 64338 279502 64574
rect 279586 64338 279822 64574
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 282986 248378 283222 248614
rect 283306 248378 283542 248614
rect 282986 248058 283222 248294
rect 283306 248058 283542 248294
rect 282986 212378 283222 212614
rect 283306 212378 283542 212614
rect 282986 212058 283222 212294
rect 283306 212058 283542 212294
rect 282986 176378 283222 176614
rect 283306 176378 283542 176614
rect 282986 176058 283222 176294
rect 283306 176058 283542 176294
rect 282986 140378 283222 140614
rect 283306 140378 283542 140614
rect 282986 140058 283222 140294
rect 283306 140058 283542 140294
rect 282986 104378 283222 104614
rect 283306 104378 283542 104614
rect 282986 104058 283222 104294
rect 283306 104058 283542 104294
rect 282986 68378 283222 68614
rect 283306 68378 283542 68614
rect 282986 68058 283222 68294
rect 283306 68058 283542 68294
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 293546 510938 293782 511174
rect 293866 510938 294102 511174
rect 293546 510618 293782 510854
rect 293866 510618 294102 510854
rect 293546 474938 293782 475174
rect 293866 474938 294102 475174
rect 293546 474618 293782 474854
rect 293866 474618 294102 474854
rect 293546 438938 293782 439174
rect 293866 438938 294102 439174
rect 293546 438618 293782 438854
rect 293866 438618 294102 438854
rect 293546 402938 293782 403174
rect 293866 402938 294102 403174
rect 293546 402618 293782 402854
rect 293866 402618 294102 402854
rect 293546 366938 293782 367174
rect 293866 366938 294102 367174
rect 293546 366618 293782 366854
rect 293866 366618 294102 366854
rect 293546 330938 293782 331174
rect 293866 330938 294102 331174
rect 293546 330618 293782 330854
rect 293866 330618 294102 330854
rect 293546 294938 293782 295174
rect 293866 294938 294102 295174
rect 293546 294618 293782 294854
rect 293866 294618 294102 294854
rect 293546 258938 293782 259174
rect 293866 258938 294102 259174
rect 293546 258618 293782 258854
rect 293866 258618 294102 258854
rect 293546 222938 293782 223174
rect 293866 222938 294102 223174
rect 293546 222618 293782 222854
rect 293866 222618 294102 222854
rect 293546 186938 293782 187174
rect 293866 186938 294102 187174
rect 293546 186618 293782 186854
rect 293866 186618 294102 186854
rect 293546 150938 293782 151174
rect 293866 150938 294102 151174
rect 293546 150618 293782 150854
rect 293866 150618 294102 150854
rect 293546 114938 293782 115174
rect 293866 114938 294102 115174
rect 293546 114618 293782 114854
rect 293866 114618 294102 114854
rect 293546 78938 293782 79174
rect 293866 78938 294102 79174
rect 293546 78618 293782 78854
rect 293866 78618 294102 78854
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 297266 514658 297502 514894
rect 297586 514658 297822 514894
rect 297266 514338 297502 514574
rect 297586 514338 297822 514574
rect 297266 478658 297502 478894
rect 297586 478658 297822 478894
rect 297266 478338 297502 478574
rect 297586 478338 297822 478574
rect 297266 442658 297502 442894
rect 297586 442658 297822 442894
rect 297266 442338 297502 442574
rect 297586 442338 297822 442574
rect 297266 406658 297502 406894
rect 297586 406658 297822 406894
rect 297266 406338 297502 406574
rect 297586 406338 297822 406574
rect 297266 370658 297502 370894
rect 297586 370658 297822 370894
rect 297266 370338 297502 370574
rect 297586 370338 297822 370574
rect 297266 334658 297502 334894
rect 297586 334658 297822 334894
rect 297266 334338 297502 334574
rect 297586 334338 297822 334574
rect 297266 298658 297502 298894
rect 297586 298658 297822 298894
rect 297266 298338 297502 298574
rect 297586 298338 297822 298574
rect 297266 262658 297502 262894
rect 297586 262658 297822 262894
rect 297266 262338 297502 262574
rect 297586 262338 297822 262574
rect 297266 226658 297502 226894
rect 297586 226658 297822 226894
rect 297266 226338 297502 226574
rect 297586 226338 297822 226574
rect 297266 190658 297502 190894
rect 297586 190658 297822 190894
rect 297266 190338 297502 190574
rect 297586 190338 297822 190574
rect 297266 154658 297502 154894
rect 297586 154658 297822 154894
rect 297266 154338 297502 154574
rect 297586 154338 297822 154574
rect 297266 118658 297502 118894
rect 297586 118658 297822 118894
rect 297266 118338 297502 118574
rect 297586 118338 297822 118574
rect 297266 82658 297502 82894
rect 297586 82658 297822 82894
rect 297266 82338 297502 82574
rect 297586 82338 297822 82574
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 300986 518378 301222 518614
rect 301306 518378 301542 518614
rect 300986 518058 301222 518294
rect 301306 518058 301542 518294
rect 300986 482378 301222 482614
rect 301306 482378 301542 482614
rect 300986 482058 301222 482294
rect 301306 482058 301542 482294
rect 300986 446378 301222 446614
rect 301306 446378 301542 446614
rect 300986 446058 301222 446294
rect 301306 446058 301542 446294
rect 300986 410378 301222 410614
rect 301306 410378 301542 410614
rect 300986 410058 301222 410294
rect 301306 410058 301542 410294
rect 300986 374378 301222 374614
rect 301306 374378 301542 374614
rect 300986 374058 301222 374294
rect 301306 374058 301542 374294
rect 300986 338378 301222 338614
rect 301306 338378 301542 338614
rect 300986 338058 301222 338294
rect 301306 338058 301542 338294
rect 300986 302378 301222 302614
rect 301306 302378 301542 302614
rect 300986 302058 301222 302294
rect 301306 302058 301542 302294
rect 300986 266378 301222 266614
rect 301306 266378 301542 266614
rect 300986 266058 301222 266294
rect 301306 266058 301542 266294
rect 300986 230378 301222 230614
rect 301306 230378 301542 230614
rect 300986 230058 301222 230294
rect 301306 230058 301542 230294
rect 300986 194378 301222 194614
rect 301306 194378 301542 194614
rect 300986 194058 301222 194294
rect 301306 194058 301542 194294
rect 300986 158378 301222 158614
rect 301306 158378 301542 158614
rect 300986 158058 301222 158294
rect 301306 158058 301542 158294
rect 300986 122378 301222 122614
rect 301306 122378 301542 122614
rect 300986 122058 301222 122294
rect 301306 122058 301542 122294
rect 300986 86378 301222 86614
rect 301306 86378 301542 86614
rect 300986 86058 301222 86294
rect 301306 86058 301542 86294
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 311546 528938 311782 529174
rect 311866 528938 312102 529174
rect 311546 528618 311782 528854
rect 311866 528618 312102 528854
rect 311546 492938 311782 493174
rect 311866 492938 312102 493174
rect 311546 492618 311782 492854
rect 311866 492618 312102 492854
rect 311546 456938 311782 457174
rect 311866 456938 312102 457174
rect 311546 456618 311782 456854
rect 311866 456618 312102 456854
rect 311546 420938 311782 421174
rect 311866 420938 312102 421174
rect 311546 420618 311782 420854
rect 311866 420618 312102 420854
rect 311546 384938 311782 385174
rect 311866 384938 312102 385174
rect 311546 384618 311782 384854
rect 311866 384618 312102 384854
rect 311546 348938 311782 349174
rect 311866 348938 312102 349174
rect 311546 348618 311782 348854
rect 311866 348618 312102 348854
rect 311546 312938 311782 313174
rect 311866 312938 312102 313174
rect 311546 312618 311782 312854
rect 311866 312618 312102 312854
rect 311546 276938 311782 277174
rect 311866 276938 312102 277174
rect 311546 276618 311782 276854
rect 311866 276618 312102 276854
rect 311546 240938 311782 241174
rect 311866 240938 312102 241174
rect 311546 240618 311782 240854
rect 311866 240618 312102 240854
rect 311546 204938 311782 205174
rect 311866 204938 312102 205174
rect 311546 204618 311782 204854
rect 311866 204618 312102 204854
rect 311546 168938 311782 169174
rect 311866 168938 312102 169174
rect 311546 168618 311782 168854
rect 311866 168618 312102 168854
rect 311546 132938 311782 133174
rect 311866 132938 312102 133174
rect 311546 132618 311782 132854
rect 311866 132618 312102 132854
rect 311546 96938 311782 97174
rect 311866 96938 312102 97174
rect 311546 96618 311782 96854
rect 311866 96618 312102 96854
rect 311546 60938 311782 61174
rect 311866 60938 312102 61174
rect 311546 60618 311782 60854
rect 311866 60618 312102 60854
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 315266 532658 315502 532894
rect 315586 532658 315822 532894
rect 315266 532338 315502 532574
rect 315586 532338 315822 532574
rect 315266 496658 315502 496894
rect 315586 496658 315822 496894
rect 315266 496338 315502 496574
rect 315586 496338 315822 496574
rect 315266 460658 315502 460894
rect 315586 460658 315822 460894
rect 315266 460338 315502 460574
rect 315586 460338 315822 460574
rect 315266 424658 315502 424894
rect 315586 424658 315822 424894
rect 315266 424338 315502 424574
rect 315586 424338 315822 424574
rect 315266 388658 315502 388894
rect 315586 388658 315822 388894
rect 315266 388338 315502 388574
rect 315586 388338 315822 388574
rect 315266 352658 315502 352894
rect 315586 352658 315822 352894
rect 315266 352338 315502 352574
rect 315586 352338 315822 352574
rect 315266 316658 315502 316894
rect 315586 316658 315822 316894
rect 315266 316338 315502 316574
rect 315586 316338 315822 316574
rect 315266 280658 315502 280894
rect 315586 280658 315822 280894
rect 315266 280338 315502 280574
rect 315586 280338 315822 280574
rect 315266 244658 315502 244894
rect 315586 244658 315822 244894
rect 315266 244338 315502 244574
rect 315586 244338 315822 244574
rect 315266 208658 315502 208894
rect 315586 208658 315822 208894
rect 315266 208338 315502 208574
rect 315586 208338 315822 208574
rect 315266 172658 315502 172894
rect 315586 172658 315822 172894
rect 315266 172338 315502 172574
rect 315586 172338 315822 172574
rect 315266 136658 315502 136894
rect 315586 136658 315822 136894
rect 315266 136338 315502 136574
rect 315586 136338 315822 136574
rect 315266 100658 315502 100894
rect 315586 100658 315822 100894
rect 315266 100338 315502 100574
rect 315586 100338 315822 100574
rect 315266 64658 315502 64894
rect 315586 64658 315822 64894
rect 315266 64338 315502 64574
rect 315586 64338 315822 64574
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 318986 536378 319222 536614
rect 319306 536378 319542 536614
rect 318986 536058 319222 536294
rect 319306 536058 319542 536294
rect 318986 500378 319222 500614
rect 319306 500378 319542 500614
rect 318986 500058 319222 500294
rect 319306 500058 319542 500294
rect 318986 464378 319222 464614
rect 319306 464378 319542 464614
rect 318986 464058 319222 464294
rect 319306 464058 319542 464294
rect 318986 428378 319222 428614
rect 319306 428378 319542 428614
rect 318986 428058 319222 428294
rect 319306 428058 319542 428294
rect 318986 392378 319222 392614
rect 319306 392378 319542 392614
rect 318986 392058 319222 392294
rect 319306 392058 319542 392294
rect 318986 356378 319222 356614
rect 319306 356378 319542 356614
rect 318986 356058 319222 356294
rect 319306 356058 319542 356294
rect 318986 320378 319222 320614
rect 319306 320378 319542 320614
rect 318986 320058 319222 320294
rect 319306 320058 319542 320294
rect 318986 284378 319222 284614
rect 319306 284378 319542 284614
rect 318986 284058 319222 284294
rect 319306 284058 319542 284294
rect 318986 248378 319222 248614
rect 319306 248378 319542 248614
rect 318986 248058 319222 248294
rect 319306 248058 319542 248294
rect 318986 212378 319222 212614
rect 319306 212378 319542 212614
rect 318986 212058 319222 212294
rect 319306 212058 319542 212294
rect 318986 176378 319222 176614
rect 319306 176378 319542 176614
rect 318986 176058 319222 176294
rect 319306 176058 319542 176294
rect 318986 140378 319222 140614
rect 319306 140378 319542 140614
rect 318986 140058 319222 140294
rect 319306 140058 319542 140294
rect 318986 104378 319222 104614
rect 319306 104378 319542 104614
rect 318986 104058 319222 104294
rect 319306 104058 319542 104294
rect 318986 68378 319222 68614
rect 319306 68378 319542 68614
rect 318986 68058 319222 68294
rect 319306 68058 319542 68294
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 329546 546938 329782 547174
rect 329866 546938 330102 547174
rect 329546 546618 329782 546854
rect 329866 546618 330102 546854
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 329546 474938 329782 475174
rect 329866 474938 330102 475174
rect 329546 474618 329782 474854
rect 329866 474618 330102 474854
rect 329546 438938 329782 439174
rect 329866 438938 330102 439174
rect 329546 438618 329782 438854
rect 329866 438618 330102 438854
rect 329546 402938 329782 403174
rect 329866 402938 330102 403174
rect 329546 402618 329782 402854
rect 329866 402618 330102 402854
rect 329546 366938 329782 367174
rect 329866 366938 330102 367174
rect 329546 366618 329782 366854
rect 329866 366618 330102 366854
rect 329546 330938 329782 331174
rect 329866 330938 330102 331174
rect 329546 330618 329782 330854
rect 329866 330618 330102 330854
rect 329546 294938 329782 295174
rect 329866 294938 330102 295174
rect 329546 294618 329782 294854
rect 329866 294618 330102 294854
rect 329546 258938 329782 259174
rect 329866 258938 330102 259174
rect 329546 258618 329782 258854
rect 329866 258618 330102 258854
rect 329546 222938 329782 223174
rect 329866 222938 330102 223174
rect 329546 222618 329782 222854
rect 329866 222618 330102 222854
rect 329546 186938 329782 187174
rect 329866 186938 330102 187174
rect 329546 186618 329782 186854
rect 329866 186618 330102 186854
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 329546 114938 329782 115174
rect 329866 114938 330102 115174
rect 329546 114618 329782 114854
rect 329866 114618 330102 114854
rect 329546 78938 329782 79174
rect 329866 78938 330102 79174
rect 329546 78618 329782 78854
rect 329866 78618 330102 78854
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 333266 550658 333502 550894
rect 333586 550658 333822 550894
rect 333266 550338 333502 550574
rect 333586 550338 333822 550574
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 333266 478658 333502 478894
rect 333586 478658 333822 478894
rect 333266 478338 333502 478574
rect 333586 478338 333822 478574
rect 333266 442658 333502 442894
rect 333586 442658 333822 442894
rect 333266 442338 333502 442574
rect 333586 442338 333822 442574
rect 333266 406658 333502 406894
rect 333586 406658 333822 406894
rect 333266 406338 333502 406574
rect 333586 406338 333822 406574
rect 333266 370658 333502 370894
rect 333586 370658 333822 370894
rect 333266 370338 333502 370574
rect 333586 370338 333822 370574
rect 333266 334658 333502 334894
rect 333586 334658 333822 334894
rect 333266 334338 333502 334574
rect 333586 334338 333822 334574
rect 333266 298658 333502 298894
rect 333586 298658 333822 298894
rect 333266 298338 333502 298574
rect 333586 298338 333822 298574
rect 333266 262658 333502 262894
rect 333586 262658 333822 262894
rect 333266 262338 333502 262574
rect 333586 262338 333822 262574
rect 333266 226658 333502 226894
rect 333586 226658 333822 226894
rect 333266 226338 333502 226574
rect 333586 226338 333822 226574
rect 333266 190658 333502 190894
rect 333586 190658 333822 190894
rect 333266 190338 333502 190574
rect 333586 190338 333822 190574
rect 333266 154658 333502 154894
rect 333586 154658 333822 154894
rect 333266 154338 333502 154574
rect 333586 154338 333822 154574
rect 333266 118658 333502 118894
rect 333586 118658 333822 118894
rect 333266 118338 333502 118574
rect 333586 118338 333822 118574
rect 333266 82658 333502 82894
rect 333586 82658 333822 82894
rect 333266 82338 333502 82574
rect 333586 82338 333822 82574
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 336986 518378 337222 518614
rect 337306 518378 337542 518614
rect 336986 518058 337222 518294
rect 337306 518058 337542 518294
rect 336986 482378 337222 482614
rect 337306 482378 337542 482614
rect 336986 482058 337222 482294
rect 337306 482058 337542 482294
rect 336986 446378 337222 446614
rect 337306 446378 337542 446614
rect 336986 446058 337222 446294
rect 337306 446058 337542 446294
rect 336986 410378 337222 410614
rect 337306 410378 337542 410614
rect 336986 410058 337222 410294
rect 337306 410058 337542 410294
rect 336986 374378 337222 374614
rect 337306 374378 337542 374614
rect 336986 374058 337222 374294
rect 337306 374058 337542 374294
rect 336986 338378 337222 338614
rect 337306 338378 337542 338614
rect 336986 338058 337222 338294
rect 337306 338058 337542 338294
rect 336986 302378 337222 302614
rect 337306 302378 337542 302614
rect 336986 302058 337222 302294
rect 337306 302058 337542 302294
rect 336986 266378 337222 266614
rect 337306 266378 337542 266614
rect 336986 266058 337222 266294
rect 337306 266058 337542 266294
rect 336986 230378 337222 230614
rect 337306 230378 337542 230614
rect 336986 230058 337222 230294
rect 337306 230058 337542 230294
rect 336986 194378 337222 194614
rect 337306 194378 337542 194614
rect 336986 194058 337222 194294
rect 337306 194058 337542 194294
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 336986 122378 337222 122614
rect 337306 122378 337542 122614
rect 336986 122058 337222 122294
rect 337306 122058 337542 122294
rect 336986 86378 337222 86614
rect 337306 86378 337542 86614
rect 336986 86058 337222 86294
rect 337306 86058 337542 86294
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 347546 564938 347782 565174
rect 347866 564938 348102 565174
rect 347546 564618 347782 564854
rect 347866 564618 348102 564854
rect 347546 528938 347782 529174
rect 347866 528938 348102 529174
rect 347546 528618 347782 528854
rect 347866 528618 348102 528854
rect 347546 492938 347782 493174
rect 347866 492938 348102 493174
rect 347546 492618 347782 492854
rect 347866 492618 348102 492854
rect 347546 456938 347782 457174
rect 347866 456938 348102 457174
rect 347546 456618 347782 456854
rect 347866 456618 348102 456854
rect 347546 420938 347782 421174
rect 347866 420938 348102 421174
rect 347546 420618 347782 420854
rect 347866 420618 348102 420854
rect 347546 384938 347782 385174
rect 347866 384938 348102 385174
rect 347546 384618 347782 384854
rect 347866 384618 348102 384854
rect 347546 348938 347782 349174
rect 347866 348938 348102 349174
rect 347546 348618 347782 348854
rect 347866 348618 348102 348854
rect 347546 312938 347782 313174
rect 347866 312938 348102 313174
rect 347546 312618 347782 312854
rect 347866 312618 348102 312854
rect 347546 276938 347782 277174
rect 347866 276938 348102 277174
rect 347546 276618 347782 276854
rect 347866 276618 348102 276854
rect 347546 240938 347782 241174
rect 347866 240938 348102 241174
rect 347546 240618 347782 240854
rect 347866 240618 348102 240854
rect 347546 204938 347782 205174
rect 347866 204938 348102 205174
rect 347546 204618 347782 204854
rect 347866 204618 348102 204854
rect 347546 168938 347782 169174
rect 347866 168938 348102 169174
rect 347546 168618 347782 168854
rect 347866 168618 348102 168854
rect 347546 132938 347782 133174
rect 347866 132938 348102 133174
rect 347546 132618 347782 132854
rect 347866 132618 348102 132854
rect 347546 96938 347782 97174
rect 347866 96938 348102 97174
rect 347546 96618 347782 96854
rect 347866 96618 348102 96854
rect 347546 60938 347782 61174
rect 347866 60938 348102 61174
rect 347546 60618 347782 60854
rect 347866 60618 348102 60854
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 351266 568658 351502 568894
rect 351586 568658 351822 568894
rect 351266 568338 351502 568574
rect 351586 568338 351822 568574
rect 351266 532658 351502 532894
rect 351586 532658 351822 532894
rect 351266 532338 351502 532574
rect 351586 532338 351822 532574
rect 351266 496658 351502 496894
rect 351586 496658 351822 496894
rect 351266 496338 351502 496574
rect 351586 496338 351822 496574
rect 351266 460658 351502 460894
rect 351586 460658 351822 460894
rect 351266 460338 351502 460574
rect 351586 460338 351822 460574
rect 351266 424658 351502 424894
rect 351586 424658 351822 424894
rect 351266 424338 351502 424574
rect 351586 424338 351822 424574
rect 351266 388658 351502 388894
rect 351586 388658 351822 388894
rect 351266 388338 351502 388574
rect 351586 388338 351822 388574
rect 351266 352658 351502 352894
rect 351586 352658 351822 352894
rect 351266 352338 351502 352574
rect 351586 352338 351822 352574
rect 351266 316658 351502 316894
rect 351586 316658 351822 316894
rect 351266 316338 351502 316574
rect 351586 316338 351822 316574
rect 351266 280658 351502 280894
rect 351586 280658 351822 280894
rect 351266 280338 351502 280574
rect 351586 280338 351822 280574
rect 351266 244658 351502 244894
rect 351586 244658 351822 244894
rect 351266 244338 351502 244574
rect 351586 244338 351822 244574
rect 351266 208658 351502 208894
rect 351586 208658 351822 208894
rect 351266 208338 351502 208574
rect 351586 208338 351822 208574
rect 351266 172658 351502 172894
rect 351586 172658 351822 172894
rect 351266 172338 351502 172574
rect 351586 172338 351822 172574
rect 351266 136658 351502 136894
rect 351586 136658 351822 136894
rect 351266 136338 351502 136574
rect 351586 136338 351822 136574
rect 351266 100658 351502 100894
rect 351586 100658 351822 100894
rect 351266 100338 351502 100574
rect 351586 100338 351822 100574
rect 351266 64658 351502 64894
rect 351586 64658 351822 64894
rect 351266 64338 351502 64574
rect 351586 64338 351822 64574
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 354986 536378 355222 536614
rect 355306 536378 355542 536614
rect 354986 536058 355222 536294
rect 355306 536058 355542 536294
rect 354986 500378 355222 500614
rect 355306 500378 355542 500614
rect 354986 500058 355222 500294
rect 355306 500058 355542 500294
rect 354986 464378 355222 464614
rect 355306 464378 355542 464614
rect 354986 464058 355222 464294
rect 355306 464058 355542 464294
rect 354986 428378 355222 428614
rect 355306 428378 355542 428614
rect 354986 428058 355222 428294
rect 355306 428058 355542 428294
rect 354986 392378 355222 392614
rect 355306 392378 355542 392614
rect 354986 392058 355222 392294
rect 355306 392058 355542 392294
rect 354986 356378 355222 356614
rect 355306 356378 355542 356614
rect 354986 356058 355222 356294
rect 355306 356058 355542 356294
rect 354986 320378 355222 320614
rect 355306 320378 355542 320614
rect 354986 320058 355222 320294
rect 355306 320058 355542 320294
rect 354986 284378 355222 284614
rect 355306 284378 355542 284614
rect 354986 284058 355222 284294
rect 355306 284058 355542 284294
rect 354986 248378 355222 248614
rect 355306 248378 355542 248614
rect 354986 248058 355222 248294
rect 355306 248058 355542 248294
rect 354986 212378 355222 212614
rect 355306 212378 355542 212614
rect 354986 212058 355222 212294
rect 355306 212058 355542 212294
rect 354986 176378 355222 176614
rect 355306 176378 355542 176614
rect 354986 176058 355222 176294
rect 355306 176058 355542 176294
rect 354986 140378 355222 140614
rect 355306 140378 355542 140614
rect 354986 140058 355222 140294
rect 355306 140058 355542 140294
rect 354986 104378 355222 104614
rect 355306 104378 355542 104614
rect 354986 104058 355222 104294
rect 355306 104058 355542 104294
rect 354986 68378 355222 68614
rect 355306 68378 355542 68614
rect 354986 68058 355222 68294
rect 355306 68058 355542 68294
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 365546 366938 365782 367174
rect 365866 366938 366102 367174
rect 365546 366618 365782 366854
rect 365866 366618 366102 366854
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 365546 294938 365782 295174
rect 365866 294938 366102 295174
rect 365546 294618 365782 294854
rect 365866 294618 366102 294854
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 369266 298658 369502 298894
rect 369586 298658 369822 298894
rect 369266 298338 369502 298574
rect 369586 298338 369822 298574
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 369266 226658 369502 226894
rect 369586 226658 369822 226894
rect 369266 226338 369502 226574
rect 369586 226338 369822 226574
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 383546 564938 383782 565174
rect 383866 564938 384102 565174
rect 383546 564618 383782 564854
rect 383866 564618 384102 564854
rect 383546 528938 383782 529174
rect 383866 528938 384102 529174
rect 383546 528618 383782 528854
rect 383866 528618 384102 528854
rect 383546 492938 383782 493174
rect 383866 492938 384102 493174
rect 383546 492618 383782 492854
rect 383866 492618 384102 492854
rect 383546 456938 383782 457174
rect 383866 456938 384102 457174
rect 383546 456618 383782 456854
rect 383866 456618 384102 456854
rect 383546 420938 383782 421174
rect 383866 420938 384102 421174
rect 383546 420618 383782 420854
rect 383866 420618 384102 420854
rect 383546 384938 383782 385174
rect 383866 384938 384102 385174
rect 383546 384618 383782 384854
rect 383866 384618 384102 384854
rect 383546 348938 383782 349174
rect 383866 348938 384102 349174
rect 383546 348618 383782 348854
rect 383866 348618 384102 348854
rect 383546 312938 383782 313174
rect 383866 312938 384102 313174
rect 383546 312618 383782 312854
rect 383866 312618 384102 312854
rect 383546 276938 383782 277174
rect 383866 276938 384102 277174
rect 383546 276618 383782 276854
rect 383866 276618 384102 276854
rect 383546 240938 383782 241174
rect 383866 240938 384102 241174
rect 383546 240618 383782 240854
rect 383866 240618 384102 240854
rect 383546 204938 383782 205174
rect 383866 204938 384102 205174
rect 383546 204618 383782 204854
rect 383866 204618 384102 204854
rect 383546 168938 383782 169174
rect 383866 168938 384102 169174
rect 383546 168618 383782 168854
rect 383866 168618 384102 168854
rect 383546 132938 383782 133174
rect 383866 132938 384102 133174
rect 383546 132618 383782 132854
rect 383866 132618 384102 132854
rect 383546 96938 383782 97174
rect 383866 96938 384102 97174
rect 383546 96618 383782 96854
rect 383866 96618 384102 96854
rect 383546 60938 383782 61174
rect 383866 60938 384102 61174
rect 383546 60618 383782 60854
rect 383866 60618 384102 60854
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 387266 568658 387502 568894
rect 387586 568658 387822 568894
rect 387266 568338 387502 568574
rect 387586 568338 387822 568574
rect 387266 532658 387502 532894
rect 387586 532658 387822 532894
rect 387266 532338 387502 532574
rect 387586 532338 387822 532574
rect 387266 496658 387502 496894
rect 387586 496658 387822 496894
rect 387266 496338 387502 496574
rect 387586 496338 387822 496574
rect 387266 460658 387502 460894
rect 387586 460658 387822 460894
rect 387266 460338 387502 460574
rect 387586 460338 387822 460574
rect 387266 424658 387502 424894
rect 387586 424658 387822 424894
rect 387266 424338 387502 424574
rect 387586 424338 387822 424574
rect 387266 388658 387502 388894
rect 387586 388658 387822 388894
rect 387266 388338 387502 388574
rect 387586 388338 387822 388574
rect 387266 352658 387502 352894
rect 387586 352658 387822 352894
rect 387266 352338 387502 352574
rect 387586 352338 387822 352574
rect 387266 316658 387502 316894
rect 387586 316658 387822 316894
rect 387266 316338 387502 316574
rect 387586 316338 387822 316574
rect 387266 280658 387502 280894
rect 387586 280658 387822 280894
rect 387266 280338 387502 280574
rect 387586 280338 387822 280574
rect 387266 244658 387502 244894
rect 387586 244658 387822 244894
rect 387266 244338 387502 244574
rect 387586 244338 387822 244574
rect 387266 208658 387502 208894
rect 387586 208658 387822 208894
rect 387266 208338 387502 208574
rect 387586 208338 387822 208574
rect 387266 172658 387502 172894
rect 387586 172658 387822 172894
rect 387266 172338 387502 172574
rect 387586 172338 387822 172574
rect 387266 136658 387502 136894
rect 387586 136658 387822 136894
rect 387266 136338 387502 136574
rect 387586 136338 387822 136574
rect 387266 100658 387502 100894
rect 387586 100658 387822 100894
rect 387266 100338 387502 100574
rect 387586 100338 387822 100574
rect 387266 64658 387502 64894
rect 387586 64658 387822 64894
rect 387266 64338 387502 64574
rect 387586 64338 387822 64574
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 390986 536378 391222 536614
rect 391306 536378 391542 536614
rect 390986 536058 391222 536294
rect 391306 536058 391542 536294
rect 390986 500378 391222 500614
rect 391306 500378 391542 500614
rect 390986 500058 391222 500294
rect 391306 500058 391542 500294
rect 390986 464378 391222 464614
rect 391306 464378 391542 464614
rect 390986 464058 391222 464294
rect 391306 464058 391542 464294
rect 390986 428378 391222 428614
rect 391306 428378 391542 428614
rect 390986 428058 391222 428294
rect 391306 428058 391542 428294
rect 390986 392378 391222 392614
rect 391306 392378 391542 392614
rect 390986 392058 391222 392294
rect 391306 392058 391542 392294
rect 390986 356378 391222 356614
rect 391306 356378 391542 356614
rect 390986 356058 391222 356294
rect 391306 356058 391542 356294
rect 390986 320378 391222 320614
rect 391306 320378 391542 320614
rect 390986 320058 391222 320294
rect 391306 320058 391542 320294
rect 390986 284378 391222 284614
rect 391306 284378 391542 284614
rect 390986 284058 391222 284294
rect 391306 284058 391542 284294
rect 390986 248378 391222 248614
rect 391306 248378 391542 248614
rect 390986 248058 391222 248294
rect 391306 248058 391542 248294
rect 390986 212378 391222 212614
rect 391306 212378 391542 212614
rect 390986 212058 391222 212294
rect 391306 212058 391542 212294
rect 390986 176378 391222 176614
rect 391306 176378 391542 176614
rect 390986 176058 391222 176294
rect 391306 176058 391542 176294
rect 390986 140378 391222 140614
rect 391306 140378 391542 140614
rect 390986 140058 391222 140294
rect 391306 140058 391542 140294
rect 390986 104378 391222 104614
rect 391306 104378 391542 104614
rect 390986 104058 391222 104294
rect 391306 104058 391542 104294
rect 390986 68378 391222 68614
rect 391306 68378 391542 68614
rect 390986 68058 391222 68294
rect 391306 68058 391542 68294
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 401546 438938 401782 439174
rect 401866 438938 402102 439174
rect 401546 438618 401782 438854
rect 401866 438618 402102 438854
rect 401546 402938 401782 403174
rect 401866 402938 402102 403174
rect 401546 402618 401782 402854
rect 401866 402618 402102 402854
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 401546 330938 401782 331174
rect 401866 330938 402102 331174
rect 401546 330618 401782 330854
rect 401866 330618 402102 330854
rect 401546 294938 401782 295174
rect 401866 294938 402102 295174
rect 401546 294618 401782 294854
rect 401866 294618 402102 294854
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 401546 222938 401782 223174
rect 401866 222938 402102 223174
rect 401546 222618 401782 222854
rect 401866 222618 402102 222854
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 405266 442658 405502 442894
rect 405586 442658 405822 442894
rect 405266 442338 405502 442574
rect 405586 442338 405822 442574
rect 405266 406658 405502 406894
rect 405586 406658 405822 406894
rect 405266 406338 405502 406574
rect 405586 406338 405822 406574
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 405266 334658 405502 334894
rect 405586 334658 405822 334894
rect 405266 334338 405502 334574
rect 405586 334338 405822 334574
rect 405266 298658 405502 298894
rect 405586 298658 405822 298894
rect 405266 298338 405502 298574
rect 405586 298338 405822 298574
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 405266 226658 405502 226894
rect 405586 226658 405822 226894
rect 405266 226338 405502 226574
rect 405586 226338 405822 226574
rect 405266 190658 405502 190894
rect 405586 190658 405822 190894
rect 405266 190338 405502 190574
rect 405586 190338 405822 190574
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 405266 118658 405502 118894
rect 405586 118658 405822 118894
rect 405266 118338 405502 118574
rect 405586 118338 405822 118574
rect 405266 82658 405502 82894
rect 405586 82658 405822 82894
rect 405266 82338 405502 82574
rect 405586 82338 405822 82574
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 408986 446378 409222 446614
rect 409306 446378 409542 446614
rect 408986 446058 409222 446294
rect 409306 446058 409542 446294
rect 408986 410378 409222 410614
rect 409306 410378 409542 410614
rect 408986 410058 409222 410294
rect 409306 410058 409542 410294
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 408986 338378 409222 338614
rect 409306 338378 409542 338614
rect 408986 338058 409222 338294
rect 409306 338058 409542 338294
rect 408986 302378 409222 302614
rect 409306 302378 409542 302614
rect 408986 302058 409222 302294
rect 409306 302058 409542 302294
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 408986 230378 409222 230614
rect 409306 230378 409542 230614
rect 408986 230058 409222 230294
rect 409306 230058 409542 230294
rect 408986 194378 409222 194614
rect 409306 194378 409542 194614
rect 408986 194058 409222 194294
rect 409306 194058 409542 194294
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 408986 86378 409222 86614
rect 409306 86378 409542 86614
rect 408986 86058 409222 86294
rect 409306 86058 409542 86294
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 419546 564938 419782 565174
rect 419866 564938 420102 565174
rect 419546 564618 419782 564854
rect 419866 564618 420102 564854
rect 419546 528938 419782 529174
rect 419866 528938 420102 529174
rect 419546 528618 419782 528854
rect 419866 528618 420102 528854
rect 419546 492938 419782 493174
rect 419866 492938 420102 493174
rect 419546 492618 419782 492854
rect 419866 492618 420102 492854
rect 419546 456938 419782 457174
rect 419866 456938 420102 457174
rect 419546 456618 419782 456854
rect 419866 456618 420102 456854
rect 419546 420938 419782 421174
rect 419866 420938 420102 421174
rect 419546 420618 419782 420854
rect 419866 420618 420102 420854
rect 419546 384938 419782 385174
rect 419866 384938 420102 385174
rect 419546 384618 419782 384854
rect 419866 384618 420102 384854
rect 419546 348938 419782 349174
rect 419866 348938 420102 349174
rect 419546 348618 419782 348854
rect 419866 348618 420102 348854
rect 419546 312938 419782 313174
rect 419866 312938 420102 313174
rect 419546 312618 419782 312854
rect 419866 312618 420102 312854
rect 419546 276938 419782 277174
rect 419866 276938 420102 277174
rect 419546 276618 419782 276854
rect 419866 276618 420102 276854
rect 419546 240938 419782 241174
rect 419866 240938 420102 241174
rect 419546 240618 419782 240854
rect 419866 240618 420102 240854
rect 419546 204938 419782 205174
rect 419866 204938 420102 205174
rect 419546 204618 419782 204854
rect 419866 204618 420102 204854
rect 419546 168938 419782 169174
rect 419866 168938 420102 169174
rect 419546 168618 419782 168854
rect 419866 168618 420102 168854
rect 419546 132938 419782 133174
rect 419866 132938 420102 133174
rect 419546 132618 419782 132854
rect 419866 132618 420102 132854
rect 419546 96938 419782 97174
rect 419866 96938 420102 97174
rect 419546 96618 419782 96854
rect 419866 96618 420102 96854
rect 419546 60938 419782 61174
rect 419866 60938 420102 61174
rect 419546 60618 419782 60854
rect 419866 60618 420102 60854
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 423266 568658 423502 568894
rect 423586 568658 423822 568894
rect 423266 568338 423502 568574
rect 423586 568338 423822 568574
rect 423266 532658 423502 532894
rect 423586 532658 423822 532894
rect 423266 532338 423502 532574
rect 423586 532338 423822 532574
rect 423266 496658 423502 496894
rect 423586 496658 423822 496894
rect 423266 496338 423502 496574
rect 423586 496338 423822 496574
rect 423266 460658 423502 460894
rect 423586 460658 423822 460894
rect 423266 460338 423502 460574
rect 423586 460338 423822 460574
rect 423266 424658 423502 424894
rect 423586 424658 423822 424894
rect 423266 424338 423502 424574
rect 423586 424338 423822 424574
rect 423266 388658 423502 388894
rect 423586 388658 423822 388894
rect 423266 388338 423502 388574
rect 423586 388338 423822 388574
rect 423266 352658 423502 352894
rect 423586 352658 423822 352894
rect 423266 352338 423502 352574
rect 423586 352338 423822 352574
rect 423266 316658 423502 316894
rect 423586 316658 423822 316894
rect 423266 316338 423502 316574
rect 423586 316338 423822 316574
rect 423266 280658 423502 280894
rect 423586 280658 423822 280894
rect 423266 280338 423502 280574
rect 423586 280338 423822 280574
rect 423266 244658 423502 244894
rect 423586 244658 423822 244894
rect 423266 244338 423502 244574
rect 423586 244338 423822 244574
rect 423266 208658 423502 208894
rect 423586 208658 423822 208894
rect 423266 208338 423502 208574
rect 423586 208338 423822 208574
rect 423266 172658 423502 172894
rect 423586 172658 423822 172894
rect 423266 172338 423502 172574
rect 423586 172338 423822 172574
rect 423266 136658 423502 136894
rect 423586 136658 423822 136894
rect 423266 136338 423502 136574
rect 423586 136338 423822 136574
rect 423266 100658 423502 100894
rect 423586 100658 423822 100894
rect 423266 100338 423502 100574
rect 423586 100338 423822 100574
rect 423266 64658 423502 64894
rect 423586 64658 423822 64894
rect 423266 64338 423502 64574
rect 423586 64338 423822 64574
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 426986 572378 427222 572614
rect 427306 572378 427542 572614
rect 426986 572058 427222 572294
rect 427306 572058 427542 572294
rect 426986 536378 427222 536614
rect 427306 536378 427542 536614
rect 426986 536058 427222 536294
rect 427306 536058 427542 536294
rect 426986 500378 427222 500614
rect 427306 500378 427542 500614
rect 426986 500058 427222 500294
rect 427306 500058 427542 500294
rect 426986 464378 427222 464614
rect 427306 464378 427542 464614
rect 426986 464058 427222 464294
rect 427306 464058 427542 464294
rect 426986 428378 427222 428614
rect 427306 428378 427542 428614
rect 426986 428058 427222 428294
rect 427306 428058 427542 428294
rect 426986 392378 427222 392614
rect 427306 392378 427542 392614
rect 426986 392058 427222 392294
rect 427306 392058 427542 392294
rect 426986 356378 427222 356614
rect 427306 356378 427542 356614
rect 426986 356058 427222 356294
rect 427306 356058 427542 356294
rect 426986 320378 427222 320614
rect 427306 320378 427542 320614
rect 426986 320058 427222 320294
rect 427306 320058 427542 320294
rect 426986 284378 427222 284614
rect 427306 284378 427542 284614
rect 426986 284058 427222 284294
rect 427306 284058 427542 284294
rect 426986 248378 427222 248614
rect 427306 248378 427542 248614
rect 426986 248058 427222 248294
rect 427306 248058 427542 248294
rect 426986 212378 427222 212614
rect 427306 212378 427542 212614
rect 426986 212058 427222 212294
rect 427306 212058 427542 212294
rect 426986 176378 427222 176614
rect 427306 176378 427542 176614
rect 426986 176058 427222 176294
rect 427306 176058 427542 176294
rect 426986 140378 427222 140614
rect 427306 140378 427542 140614
rect 426986 140058 427222 140294
rect 427306 140058 427542 140294
rect 426986 104378 427222 104614
rect 427306 104378 427542 104614
rect 426986 104058 427222 104294
rect 427306 104058 427542 104294
rect 426986 68378 427222 68614
rect 427306 68378 427542 68614
rect 426986 68058 427222 68294
rect 427306 68058 427542 68294
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 437546 438938 437782 439174
rect 437866 438938 438102 439174
rect 437546 438618 437782 438854
rect 437866 438618 438102 438854
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 437546 294938 437782 295174
rect 437866 294938 438102 295174
rect 437546 294618 437782 294854
rect 437866 294618 438102 294854
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 437546 114938 437782 115174
rect 437866 114938 438102 115174
rect 437546 114618 437782 114854
rect 437866 114618 438102 114854
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 441266 442658 441502 442894
rect 441586 442658 441822 442894
rect 441266 442338 441502 442574
rect 441586 442338 441822 442574
rect 441266 406658 441502 406894
rect 441586 406658 441822 406894
rect 441266 406338 441502 406574
rect 441586 406338 441822 406574
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 441266 334658 441502 334894
rect 441586 334658 441822 334894
rect 441266 334338 441502 334574
rect 441586 334338 441822 334574
rect 441266 298658 441502 298894
rect 441586 298658 441822 298894
rect 441266 298338 441502 298574
rect 441586 298338 441822 298574
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 441266 226658 441502 226894
rect 441586 226658 441822 226894
rect 441266 226338 441502 226574
rect 441586 226338 441822 226574
rect 441266 190658 441502 190894
rect 441586 190658 441822 190894
rect 441266 190338 441502 190574
rect 441586 190338 441822 190574
rect 441266 154658 441502 154894
rect 441586 154658 441822 154894
rect 441266 154338 441502 154574
rect 441586 154338 441822 154574
rect 441266 118658 441502 118894
rect 441586 118658 441822 118894
rect 441266 118338 441502 118574
rect 441586 118338 441822 118574
rect 441266 82658 441502 82894
rect 441586 82658 441822 82894
rect 441266 82338 441502 82574
rect 441586 82338 441822 82574
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 444986 410378 445222 410614
rect 445306 410378 445542 410614
rect 444986 410058 445222 410294
rect 445306 410058 445542 410294
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 444986 302378 445222 302614
rect 445306 302378 445542 302614
rect 444986 302058 445222 302294
rect 445306 302058 445542 302294
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 444986 122378 445222 122614
rect 445306 122378 445542 122614
rect 444986 122058 445222 122294
rect 445306 122058 445542 122294
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 455546 528938 455782 529174
rect 455866 528938 456102 529174
rect 455546 528618 455782 528854
rect 455866 528618 456102 528854
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 455546 456938 455782 457174
rect 455866 456938 456102 457174
rect 455546 456618 455782 456854
rect 455866 456618 456102 456854
rect 455546 420938 455782 421174
rect 455866 420938 456102 421174
rect 455546 420618 455782 420854
rect 455866 420618 456102 420854
rect 455546 384938 455782 385174
rect 455866 384938 456102 385174
rect 455546 384618 455782 384854
rect 455866 384618 456102 384854
rect 455546 348938 455782 349174
rect 455866 348938 456102 349174
rect 455546 348618 455782 348854
rect 455866 348618 456102 348854
rect 455546 312938 455782 313174
rect 455866 312938 456102 313174
rect 455546 312618 455782 312854
rect 455866 312618 456102 312854
rect 455546 276938 455782 277174
rect 455866 276938 456102 277174
rect 455546 276618 455782 276854
rect 455866 276618 456102 276854
rect 455546 240938 455782 241174
rect 455866 240938 456102 241174
rect 455546 240618 455782 240854
rect 455866 240618 456102 240854
rect 455546 204938 455782 205174
rect 455866 204938 456102 205174
rect 455546 204618 455782 204854
rect 455866 204618 456102 204854
rect 455546 168938 455782 169174
rect 455866 168938 456102 169174
rect 455546 168618 455782 168854
rect 455866 168618 456102 168854
rect 455546 132938 455782 133174
rect 455866 132938 456102 133174
rect 455546 132618 455782 132854
rect 455866 132618 456102 132854
rect 455546 96938 455782 97174
rect 455866 96938 456102 97174
rect 455546 96618 455782 96854
rect 455866 96618 456102 96854
rect 455546 60938 455782 61174
rect 455866 60938 456102 61174
rect 455546 60618 455782 60854
rect 455866 60618 456102 60854
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 459266 532658 459502 532894
rect 459586 532658 459822 532894
rect 459266 532338 459502 532574
rect 459586 532338 459822 532574
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 459266 460658 459502 460894
rect 459586 460658 459822 460894
rect 459266 460338 459502 460574
rect 459586 460338 459822 460574
rect 459266 424658 459502 424894
rect 459586 424658 459822 424894
rect 459266 424338 459502 424574
rect 459586 424338 459822 424574
rect 459266 388658 459502 388894
rect 459586 388658 459822 388894
rect 459266 388338 459502 388574
rect 459586 388338 459822 388574
rect 459266 352658 459502 352894
rect 459586 352658 459822 352894
rect 459266 352338 459502 352574
rect 459586 352338 459822 352574
rect 459266 316658 459502 316894
rect 459586 316658 459822 316894
rect 459266 316338 459502 316574
rect 459586 316338 459822 316574
rect 459266 280658 459502 280894
rect 459586 280658 459822 280894
rect 459266 280338 459502 280574
rect 459586 280338 459822 280574
rect 459266 244658 459502 244894
rect 459586 244658 459822 244894
rect 459266 244338 459502 244574
rect 459586 244338 459822 244574
rect 459266 208658 459502 208894
rect 459586 208658 459822 208894
rect 459266 208338 459502 208574
rect 459586 208338 459822 208574
rect 459266 172658 459502 172894
rect 459586 172658 459822 172894
rect 459266 172338 459502 172574
rect 459586 172338 459822 172574
rect 459266 136658 459502 136894
rect 459586 136658 459822 136894
rect 459266 136338 459502 136574
rect 459586 136338 459822 136574
rect 459266 100658 459502 100894
rect 459586 100658 459822 100894
rect 459266 100338 459502 100574
rect 459586 100338 459822 100574
rect 459266 64658 459502 64894
rect 459586 64658 459822 64894
rect 459266 64338 459502 64574
rect 459586 64338 459822 64574
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 462986 536378 463222 536614
rect 463306 536378 463542 536614
rect 462986 536058 463222 536294
rect 463306 536058 463542 536294
rect 462986 500378 463222 500614
rect 463306 500378 463542 500614
rect 462986 500058 463222 500294
rect 463306 500058 463542 500294
rect 462986 464378 463222 464614
rect 463306 464378 463542 464614
rect 462986 464058 463222 464294
rect 463306 464058 463542 464294
rect 462986 428378 463222 428614
rect 463306 428378 463542 428614
rect 462986 428058 463222 428294
rect 463306 428058 463542 428294
rect 462986 392378 463222 392614
rect 463306 392378 463542 392614
rect 462986 392058 463222 392294
rect 463306 392058 463542 392294
rect 462986 356378 463222 356614
rect 463306 356378 463542 356614
rect 462986 356058 463222 356294
rect 463306 356058 463542 356294
rect 462986 320378 463222 320614
rect 463306 320378 463542 320614
rect 462986 320058 463222 320294
rect 463306 320058 463542 320294
rect 462986 284378 463222 284614
rect 463306 284378 463542 284614
rect 462986 284058 463222 284294
rect 463306 284058 463542 284294
rect 462986 248378 463222 248614
rect 463306 248378 463542 248614
rect 462986 248058 463222 248294
rect 463306 248058 463542 248294
rect 462986 212378 463222 212614
rect 463306 212378 463542 212614
rect 462986 212058 463222 212294
rect 463306 212058 463542 212294
rect 462986 176378 463222 176614
rect 463306 176378 463542 176614
rect 462986 176058 463222 176294
rect 463306 176058 463542 176294
rect 462986 140378 463222 140614
rect 463306 140378 463542 140614
rect 462986 140058 463222 140294
rect 463306 140058 463542 140294
rect 462986 104378 463222 104614
rect 463306 104378 463542 104614
rect 462986 104058 463222 104294
rect 463306 104058 463542 104294
rect 462986 68378 463222 68614
rect 463306 68378 463542 68614
rect 462986 68058 463222 68294
rect 463306 68058 463542 68294
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 477266 334658 477502 334894
rect 477586 334658 477822 334894
rect 477266 334338 477502 334574
rect 477586 334338 477822 334574
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 477266 226658 477502 226894
rect 477586 226658 477822 226894
rect 477266 226338 477502 226574
rect 477586 226338 477822 226574
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 480986 410378 481222 410614
rect 481306 410378 481542 410614
rect 480986 410058 481222 410294
rect 481306 410058 481542 410294
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 480986 338378 481222 338614
rect 481306 338378 481542 338614
rect 480986 338058 481222 338294
rect 481306 338058 481542 338294
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 491546 456938 491782 457174
rect 491866 456938 492102 457174
rect 491546 456618 491782 456854
rect 491866 456618 492102 456854
rect 491546 420938 491782 421174
rect 491866 420938 492102 421174
rect 491546 420618 491782 420854
rect 491866 420618 492102 420854
rect 491546 384938 491782 385174
rect 491866 384938 492102 385174
rect 491546 384618 491782 384854
rect 491866 384618 492102 384854
rect 491546 348938 491782 349174
rect 491866 348938 492102 349174
rect 491546 348618 491782 348854
rect 491866 348618 492102 348854
rect 491546 312938 491782 313174
rect 491866 312938 492102 313174
rect 491546 312618 491782 312854
rect 491866 312618 492102 312854
rect 491546 276938 491782 277174
rect 491866 276938 492102 277174
rect 491546 276618 491782 276854
rect 491866 276618 492102 276854
rect 491546 240938 491782 241174
rect 491866 240938 492102 241174
rect 491546 240618 491782 240854
rect 491866 240618 492102 240854
rect 491546 204938 491782 205174
rect 491866 204938 492102 205174
rect 491546 204618 491782 204854
rect 491866 204618 492102 204854
rect 491546 168938 491782 169174
rect 491866 168938 492102 169174
rect 491546 168618 491782 168854
rect 491866 168618 492102 168854
rect 491546 132938 491782 133174
rect 491866 132938 492102 133174
rect 491546 132618 491782 132854
rect 491866 132618 492102 132854
rect 491546 96938 491782 97174
rect 491866 96938 492102 97174
rect 491546 96618 491782 96854
rect 491866 96618 492102 96854
rect 491546 60938 491782 61174
rect 491866 60938 492102 61174
rect 491546 60618 491782 60854
rect 491866 60618 492102 60854
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 495266 460658 495502 460894
rect 495586 460658 495822 460894
rect 495266 460338 495502 460574
rect 495586 460338 495822 460574
rect 495266 424658 495502 424894
rect 495586 424658 495822 424894
rect 495266 424338 495502 424574
rect 495586 424338 495822 424574
rect 495266 388658 495502 388894
rect 495586 388658 495822 388894
rect 495266 388338 495502 388574
rect 495586 388338 495822 388574
rect 495266 352658 495502 352894
rect 495586 352658 495822 352894
rect 495266 352338 495502 352574
rect 495586 352338 495822 352574
rect 495266 316658 495502 316894
rect 495586 316658 495822 316894
rect 495266 316338 495502 316574
rect 495586 316338 495822 316574
rect 495266 280658 495502 280894
rect 495586 280658 495822 280894
rect 495266 280338 495502 280574
rect 495586 280338 495822 280574
rect 495266 244658 495502 244894
rect 495586 244658 495822 244894
rect 495266 244338 495502 244574
rect 495586 244338 495822 244574
rect 495266 208658 495502 208894
rect 495586 208658 495822 208894
rect 495266 208338 495502 208574
rect 495586 208338 495822 208574
rect 495266 172658 495502 172894
rect 495586 172658 495822 172894
rect 495266 172338 495502 172574
rect 495586 172338 495822 172574
rect 495266 136658 495502 136894
rect 495586 136658 495822 136894
rect 495266 136338 495502 136574
rect 495586 136338 495822 136574
rect 495266 100658 495502 100894
rect 495586 100658 495822 100894
rect 495266 100338 495502 100574
rect 495586 100338 495822 100574
rect 495266 64658 495502 64894
rect 495586 64658 495822 64894
rect 495266 64338 495502 64574
rect 495586 64338 495822 64574
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 498986 608378 499222 608614
rect 499306 608378 499542 608614
rect 498986 608058 499222 608294
rect 499306 608058 499542 608294
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 498986 464378 499222 464614
rect 499306 464378 499542 464614
rect 498986 464058 499222 464294
rect 499306 464058 499542 464294
rect 498986 428378 499222 428614
rect 499306 428378 499542 428614
rect 498986 428058 499222 428294
rect 499306 428058 499542 428294
rect 498986 392378 499222 392614
rect 499306 392378 499542 392614
rect 498986 392058 499222 392294
rect 499306 392058 499542 392294
rect 498986 356378 499222 356614
rect 499306 356378 499542 356614
rect 498986 356058 499222 356294
rect 499306 356058 499542 356294
rect 498986 320378 499222 320614
rect 499306 320378 499542 320614
rect 498986 320058 499222 320294
rect 499306 320058 499542 320294
rect 498986 284378 499222 284614
rect 499306 284378 499542 284614
rect 498986 284058 499222 284294
rect 499306 284058 499542 284294
rect 498986 248378 499222 248614
rect 499306 248378 499542 248614
rect 498986 248058 499222 248294
rect 499306 248058 499542 248294
rect 498986 212378 499222 212614
rect 499306 212378 499542 212614
rect 498986 212058 499222 212294
rect 499306 212058 499542 212294
rect 498986 176378 499222 176614
rect 499306 176378 499542 176614
rect 498986 176058 499222 176294
rect 499306 176058 499542 176294
rect 498986 140378 499222 140614
rect 499306 140378 499542 140614
rect 498986 140058 499222 140294
rect 499306 140058 499542 140294
rect 498986 104378 499222 104614
rect 499306 104378 499542 104614
rect 498986 104058 499222 104294
rect 499306 104058 499542 104294
rect 498986 68378 499222 68614
rect 499306 68378 499542 68614
rect 498986 68058 499222 68294
rect 499306 68058 499542 68294
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 77686 561454
rect 77922 561218 85617 561454
rect 85853 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 77686 561134
rect 77922 560898 85617 561134
rect 85853 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73721 543454
rect 73957 543218 81651 543454
rect 81887 543218 89582 543454
rect 89818 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73721 543134
rect 73957 542898 81651 543134
rect 81887 542898 89582 543134
rect 89818 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 197818 435454
rect 198054 435218 228538 435454
rect 228774 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 197818 435134
rect 198054 434898 228538 435134
rect 228774 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 88380 417454
rect 88616 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 213178 417454
rect 213414 417218 243898 417454
rect 244134 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 88380 417134
rect 88616 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 213178 417134
rect 213414 416898 243898 417134
rect 244134 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73020 399454
rect 73256 399218 103740 399454
rect 103976 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 197818 399454
rect 198054 399218 228538 399454
rect 228774 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73020 399134
rect 73256 398898 103740 399134
rect 103976 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 197818 399134
rect 198054 398898 228538 399134
rect 228774 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 197818 291454
rect 198054 291218 228538 291454
rect 228774 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 197818 291134
rect 198054 290898 228538 291134
rect 228774 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 79019 273454
rect 79255 273218 88283 273454
rect 88519 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 213178 273454
rect 213414 273218 243898 273454
rect 244134 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 79019 273134
rect 79255 272898 88283 273134
rect 88519 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 213178 273134
rect 213414 272898 243898 273134
rect 244134 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 74387 255454
rect 74623 255218 83651 255454
rect 83887 255218 92915 255454
rect 93151 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 197818 255454
rect 198054 255218 228538 255454
rect 228774 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 74387 255134
rect 74623 254898 83651 255134
rect 83887 254898 92915 255134
rect 93151 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 197818 255134
rect 198054 254898 228538 255134
rect 228774 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 102986 176614
rect 103222 176378 103306 176614
rect 103542 176378 138986 176614
rect 139222 176378 139306 176614
rect 139542 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 102986 176294
rect 103222 176058 103306 176294
rect 103542 176058 138986 176294
rect 139222 176058 139306 176294
rect 139542 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 99266 172894
rect 99502 172658 99586 172894
rect 99822 172658 135266 172894
rect 135502 172658 135586 172894
rect 135822 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 279266 172894
rect 279502 172658 279586 172894
rect 279822 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 99266 172574
rect 99502 172338 99586 172574
rect 99822 172338 135266 172574
rect 135502 172338 135586 172574
rect 135822 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 279266 172574
rect 279502 172338 279586 172574
rect 279822 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 95546 169174
rect 95782 168938 95866 169174
rect 96102 168938 131546 169174
rect 131782 168938 131866 169174
rect 132102 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 275546 169174
rect 275782 168938 275866 169174
rect 276102 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 95546 168854
rect 95782 168618 95866 168854
rect 96102 168618 131546 168854
rect 131782 168618 131866 168854
rect 132102 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 275546 168854
rect 275782 168618 275866 168854
rect 276102 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 102986 140614
rect 103222 140378 103306 140614
rect 103542 140378 138986 140614
rect 139222 140378 139306 140614
rect 139542 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 102986 140294
rect 103222 140058 103306 140294
rect 103542 140058 138986 140294
rect 139222 140058 139306 140294
rect 139542 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 99266 136894
rect 99502 136658 99586 136894
rect 99822 136658 135266 136894
rect 135502 136658 135586 136894
rect 135822 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 279266 136894
rect 279502 136658 279586 136894
rect 279822 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 99266 136574
rect 99502 136338 99586 136574
rect 99822 136338 135266 136574
rect 135502 136338 135586 136574
rect 135822 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 279266 136574
rect 279502 136338 279586 136574
rect 279822 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 131546 133174
rect 131782 132938 131866 133174
rect 132102 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 131546 132854
rect 131782 132618 131866 132854
rect 132102 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 77686 129454
rect 77922 129218 85617 129454
rect 85853 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 204306 129454
rect 204542 129218 214058 129454
rect 214294 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 77686 129134
rect 77922 128898 85617 129134
rect 85853 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 204306 129134
rect 204542 128898 214058 129134
rect 214294 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73721 111454
rect 73957 111218 81651 111454
rect 81887 111218 89582 111454
rect 89818 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 199430 111454
rect 199666 111218 209182 111454
rect 209418 111218 218934 111454
rect 219170 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73721 111134
rect 73957 110898 81651 111134
rect 81887 110898 89582 111134
rect 89818 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 199430 111134
rect 199666 110898 209182 111134
rect 209418 110898 218934 111134
rect 219170 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 102986 104614
rect 103222 104378 103306 104614
rect 103542 104378 138986 104614
rect 139222 104378 139306 104614
rect 139542 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 102986 104294
rect 103222 104058 103306 104294
rect 103542 104058 138986 104294
rect 139222 104058 139306 104294
rect 139542 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 99266 100894
rect 99502 100658 99586 100894
rect 99822 100658 135266 100894
rect 135502 100658 135586 100894
rect 135822 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 279266 100894
rect 279502 100658 279586 100894
rect 279822 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 99266 100574
rect 99502 100338 99586 100574
rect 99822 100338 135266 100574
rect 135502 100338 135586 100574
rect 135822 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 279266 100574
rect 279502 100338 279586 100574
rect 279822 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 131546 97174
rect 131782 96938 131866 97174
rect 132102 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 131546 96854
rect 131782 96618 131866 96854
rect 132102 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use zube_wrapped_project  zube_wrapped_project_5
timestamp 1635332755
transform 1 0 193568 0 1 241592
box 0 0 60000 60000
use wrapped_ws2812  wrapped_ws2812_4
timestamp 1635332755
transform 1 0 193568 0 1 92782
box 0 0 31475 48253
use wrapped_vga_clock  wrapped_vga_clock_2
timestamp 1635332755
transform 1 0 68770 0 1 390356
box 0 0 44000 44000
use wrapped_tpm2137  wrapped_tpm2137_3
timestamp 1635332755
transform 1 0 68770 0 1 539166
box 0 0 26000 42000
use wrapped_rgb_mixer  wrapped_rgb_mixer_0
timestamp 1635332755
transform 1 0 68770 0 1 92782
box 0 0 26000 42000
use wrapped_hack_soc  wrapped_hack_soc_6
timestamp 1635332755
transform 1 0 193568 0 1 390356
box 0 0 60000 60000
use wrapped_frequency_counter  wrapped_frequency_counter_1
timestamp 1635332755
transform 1 0 68770 0 1 241592
box 0 0 30000 42000
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 90782 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 90782 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 136782 74414 239592 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 143035 218414 239592 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 239592 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 285592 74414 388356 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 388356 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 303592 218414 388356 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 303592 254414 388356 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 436356 74414 537166 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 583166 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 436356 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 452356 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 452356 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 90782 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 90782 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 136782 78134 239592 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 143035 222134 239592 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 285592 78134 388356 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 388356 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 303592 222134 388356 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 436356 78134 537166 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 583166 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 436356 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 452356 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 90782 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 90782 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 136782 81854 239592 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 143035 225854 239592 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 285592 81854 388356 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 303592 225854 388356 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 436356 81854 537166 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 583166 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 452356 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 90782 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 90782 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 136782 85574 239592 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 143035 193574 239592 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 239592 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 285592 85574 388356 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 303592 193574 388356 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 303592 229574 388356 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 436356 85574 537166 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 583166 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 452356 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 452356 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 90782 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 239592 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 143035 207854 239592 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 239592 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 285592 99854 388356 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 303592 207854 388356 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 303592 243854 388356 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 436356 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 452356 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 452356 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 90782 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 90782 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 136782 67574 239592 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 143035 211574 239592 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 239592 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 285592 67574 388356 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 388356 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 303592 211574 388356 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 303592 247574 388356 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 436356 67574 537166 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 583166 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 436356 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 452356 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 452356 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 90782 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 90782 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 136782 92414 239592 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 143035 200414 239592 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 239592 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 285592 92414 388356 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 303592 200414 388356 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 303592 236414 388356 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 436356 92414 537166 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 583166 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 452356 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 452356 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 90782 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 90782 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 136782 96134 239592 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 143035 204134 239592 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 239592 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 285592 96134 388356 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 303592 204134 388356 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 303592 240134 388356 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 436356 96134 537166 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 583166 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 452356 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 452356 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
