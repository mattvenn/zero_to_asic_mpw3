magic
tech sky130A
magscale 1 2
timestamp 1635266113
<< metal1 >>
rect 264238 703332 264244 703384
rect 264296 703372 264302 703384
rect 332502 703372 332508 703384
rect 264296 703344 332508 703372
rect 264296 703332 264302 703344
rect 332502 703332 332508 703344
rect 332560 703332 332566 703384
rect 70302 703264 70308 703316
rect 70360 703304 70366 703316
rect 154114 703304 154120 703316
rect 70360 703276 154120 703304
rect 70360 703264 70366 703276
rect 154114 703264 154120 703276
rect 154172 703264 154178 703316
rect 282178 703264 282184 703316
rect 282236 703304 282242 703316
rect 397454 703304 397460 703316
rect 282236 703276 397460 703304
rect 282236 703264 282242 703276
rect 397454 703264 397460 703276
rect 397512 703264 397518 703316
rect 90358 703196 90364 703248
rect 90416 703236 90422 703248
rect 235166 703236 235172 703248
rect 90416 703208 235172 703236
rect 90416 703196 90422 703208
rect 235166 703196 235172 703208
rect 235224 703196 235230 703248
rect 273898 703196 273904 703248
rect 273956 703236 273962 703248
rect 413646 703236 413652 703248
rect 273956 703208 413652 703236
rect 273956 703196 273962 703208
rect 413646 703196 413652 703208
rect 413704 703196 413710 703248
rect 119338 703128 119344 703180
rect 119396 703168 119402 703180
rect 218974 703168 218980 703180
rect 119396 703140 218980 703168
rect 119396 703128 119402 703140
rect 218974 703128 218980 703140
rect 219032 703128 219038 703180
rect 280798 703128 280804 703180
rect 280856 703168 280862 703180
rect 462314 703168 462320 703180
rect 280856 703140 462320 703168
rect 280856 703128 280862 703140
rect 462314 703128 462320 703140
rect 462372 703128 462378 703180
rect 102042 703060 102048 703112
rect 102100 703100 102106 703112
rect 300118 703100 300124 703112
rect 102100 703072 300124 703100
rect 102100 703060 102106 703072
rect 300118 703060 300124 703072
rect 300176 703060 300182 703112
rect 67634 702992 67640 703044
rect 67692 703032 67698 703044
rect 170306 703032 170312 703044
rect 67692 703004 170312 703032
rect 67692 702992 67698 703004
rect 170306 702992 170312 703004
rect 170364 702992 170370 703044
rect 287698 702992 287704 703044
rect 287756 703032 287762 703044
rect 580166 703032 580172 703044
rect 287756 703004 580172 703032
rect 287756 702992 287762 703004
rect 580166 702992 580172 703004
rect 580224 702992 580230 703044
rect 71774 702924 71780 702976
rect 71832 702964 71838 702976
rect 72970 702964 72976 702976
rect 71832 702936 72976 702964
rect 71832 702924 71838 702936
rect 72970 702924 72976 702936
rect 73028 702924 73034 702976
rect 84102 702924 84108 702976
rect 84160 702964 84166 702976
rect 202782 702964 202788 702976
rect 84160 702936 202788 702964
rect 84160 702924 84166 702936
rect 202782 702924 202788 702936
rect 202840 702924 202846 702976
rect 286318 702924 286324 702976
rect 286376 702964 286382 702976
rect 543458 702964 543464 702976
rect 286376 702936 543464 702964
rect 286376 702924 286382 702936
rect 543458 702924 543464 702936
rect 543516 702924 543522 702976
rect 61930 702856 61936 702908
rect 61988 702896 61994 702908
rect 364978 702896 364984 702908
rect 61988 702868 364984 702896
rect 61988 702856 61994 702868
rect 364978 702856 364984 702868
rect 365036 702856 365042 702908
rect 97258 702788 97264 702840
rect 97316 702828 97322 702840
rect 478506 702828 478512 702840
rect 97316 702800 478512 702828
rect 97316 702788 97322 702800
rect 478506 702788 478512 702800
rect 478564 702788 478570 702840
rect 24302 702720 24308 702772
rect 24360 702760 24366 702772
rect 86218 702760 86224 702772
rect 24360 702732 86224 702760
rect 24360 702720 24366 702732
rect 86218 702720 86224 702732
rect 86276 702720 86282 702772
rect 116578 702720 116584 702772
rect 116636 702760 116642 702772
rect 429838 702760 429844 702772
rect 116636 702732 429844 702760
rect 116636 702720 116642 702732
rect 429838 702720 429844 702732
rect 429896 702720 429902 702772
rect 77202 702652 77208 702704
rect 77260 702692 77266 702704
rect 494790 702692 494796 702704
rect 77260 702664 494796 702692
rect 77260 702652 77266 702664
rect 494790 702652 494796 702664
rect 494848 702652 494854 702704
rect 8110 702584 8116 702636
rect 8168 702624 8174 702636
rect 94682 702624 94688 702636
rect 8168 702596 94688 702624
rect 8168 702584 8174 702596
rect 94682 702584 94688 702596
rect 94740 702584 94746 702636
rect 105630 702584 105636 702636
rect 105688 702624 105694 702636
rect 527174 702624 527180 702636
rect 105688 702596 527180 702624
rect 105688 702584 105694 702596
rect 527174 702584 527180 702596
rect 527232 702584 527238 702636
rect 57790 702516 57796 702568
rect 57848 702556 57854 702568
rect 582374 702556 582380 702568
rect 57848 702528 582380 702556
rect 57848 702516 57854 702528
rect 582374 702516 582380 702528
rect 582432 702516 582438 702568
rect 66070 702448 66076 702500
rect 66128 702488 66134 702500
rect 559650 702488 559656 702500
rect 66128 702460 559656 702488
rect 66128 702448 66134 702460
rect 559650 702448 559656 702460
rect 559708 702448 559714 702500
rect 71682 700272 71688 700324
rect 71740 700312 71746 700324
rect 105446 700312 105452 700324
rect 71740 700284 105452 700312
rect 71740 700272 71746 700284
rect 105446 700272 105452 700284
rect 105504 700272 105510 700324
rect 277302 700272 277308 700324
rect 277360 700312 277366 700324
rect 283834 700312 283840 700324
rect 277360 700284 283840 700312
rect 277360 700272 277366 700284
rect 283834 700272 283840 700284
rect 283892 700272 283898 700324
rect 87598 699660 87604 699712
rect 87656 699700 87662 699712
rect 89162 699700 89168 699712
rect 87656 699672 89168 699700
rect 87656 699660 87662 699672
rect 89162 699660 89168 699672
rect 89220 699660 89226 699712
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 17218 670732 17224 670744
rect 3568 670704 17224 670732
rect 3568 670692 3574 670704
rect 17218 670692 17224 670704
rect 17276 670692 17282 670744
rect 3510 656888 3516 656940
rect 3568 656928 3574 656940
rect 15838 656928 15844 656940
rect 3568 656900 15844 656928
rect 3568 656888 3574 656900
rect 15838 656888 15844 656900
rect 15896 656888 15902 656940
rect 3510 632068 3516 632120
rect 3568 632108 3574 632120
rect 21358 632108 21364 632120
rect 3568 632080 21364 632108
rect 3568 632068 3574 632080
rect 21358 632068 21364 632080
rect 21416 632068 21422 632120
rect 3510 618264 3516 618316
rect 3568 618304 3574 618316
rect 43438 618304 43444 618316
rect 3568 618276 43444 618304
rect 3568 618264 3574 618276
rect 43438 618264 43444 618276
rect 43496 618264 43502 618316
rect 2774 605888 2780 605940
rect 2832 605928 2838 605940
rect 4798 605928 4804 605940
rect 2832 605900 4804 605928
rect 2832 605888 2838 605900
rect 4798 605888 4804 605900
rect 4856 605888 4862 605940
rect 67542 589908 67548 589960
rect 67600 589948 67606 589960
rect 71682 589948 71688 589960
rect 67600 589920 71688 589948
rect 67600 589908 67606 589920
rect 71682 589908 71688 589920
rect 71740 589948 71746 589960
rect 124214 589948 124220 589960
rect 71740 589920 124220 589948
rect 71740 589908 71746 589920
rect 124214 589908 124220 589920
rect 124272 589908 124278 589960
rect 40034 588548 40040 588600
rect 40092 588588 40098 588600
rect 95326 588588 95332 588600
rect 40092 588560 95332 588588
rect 40092 588548 40098 588560
rect 95326 588548 95332 588560
rect 95384 588548 95390 588600
rect 84102 587868 84108 587920
rect 84160 587908 84166 587920
rect 101398 587908 101404 587920
rect 84160 587880 101404 587908
rect 84160 587868 84166 587880
rect 101398 587868 101404 587880
rect 101456 587868 101462 587920
rect 4798 587120 4804 587172
rect 4856 587160 4862 587172
rect 96614 587160 96620 587172
rect 4856 587132 96620 587160
rect 4856 587120 4862 587132
rect 96614 587120 96620 587132
rect 96672 587120 96678 587172
rect 86494 586508 86500 586560
rect 86552 586548 86558 586560
rect 140774 586548 140780 586560
rect 86552 586520 140780 586548
rect 86552 586508 86558 586520
rect 140774 586508 140780 586520
rect 140832 586508 140838 586560
rect 78582 585760 78588 585812
rect 78640 585800 78646 585812
rect 87598 585800 87604 585812
rect 78640 585772 87604 585800
rect 78640 585760 78646 585772
rect 87598 585760 87604 585772
rect 87656 585760 87662 585812
rect 121730 585760 121736 585812
rect 121788 585800 121794 585812
rect 582650 585800 582656 585812
rect 121788 585772 582656 585800
rect 121788 585760 121794 585772
rect 582650 585760 582656 585772
rect 582708 585760 582714 585812
rect 82722 585216 82728 585268
rect 82780 585256 82786 585268
rect 98638 585256 98644 585268
rect 82780 585228 98644 585256
rect 82780 585216 82786 585228
rect 98638 585216 98644 585228
rect 98696 585216 98702 585268
rect 55122 585148 55128 585200
rect 55180 585188 55186 585200
rect 77938 585188 77944 585200
rect 55180 585160 77944 585188
rect 55180 585148 55186 585160
rect 77938 585148 77944 585160
rect 77996 585188 78002 585200
rect 78582 585188 78588 585200
rect 77996 585160 78588 585188
rect 77996 585148 78002 585160
rect 78582 585148 78588 585160
rect 78640 585148 78646 585200
rect 87506 585148 87512 585200
rect 87564 585188 87570 585200
rect 121454 585188 121460 585200
rect 87564 585160 121460 585188
rect 87564 585148 87570 585160
rect 121454 585148 121460 585160
rect 121512 585188 121518 585200
rect 121730 585188 121736 585200
rect 121512 585160 121736 585188
rect 121512 585148 121518 585160
rect 121730 585148 121736 585160
rect 121788 585148 121794 585200
rect 92106 583788 92112 583840
rect 92164 583828 92170 583840
rect 92164 583800 122834 583828
rect 92164 583788 92170 583800
rect 122806 583772 122834 583800
rect 73522 583720 73528 583772
rect 73580 583760 73586 583772
rect 111058 583760 111064 583772
rect 73580 583732 111064 583760
rect 73580 583720 73586 583732
rect 111058 583720 111064 583732
rect 111116 583720 111122 583772
rect 122806 583732 122840 583772
rect 122834 583720 122840 583732
rect 122892 583760 122898 583772
rect 582834 583760 582840 583772
rect 122892 583732 582840 583760
rect 122892 583720 122898 583732
rect 582834 583720 582840 583732
rect 582892 583720 582898 583772
rect 81802 582564 81808 582616
rect 81860 582604 81866 582616
rect 84102 582604 84108 582616
rect 81860 582576 84108 582604
rect 81860 582564 81866 582576
rect 84102 582564 84108 582576
rect 84160 582564 84166 582616
rect 62022 582428 62028 582480
rect 62080 582468 62086 582480
rect 73798 582468 73804 582480
rect 62080 582440 73804 582468
rect 62080 582428 62086 582440
rect 73798 582428 73804 582440
rect 73856 582428 73862 582480
rect 93762 582428 93768 582480
rect 93820 582468 93826 582480
rect 105538 582468 105544 582480
rect 93820 582440 105544 582468
rect 93820 582428 93826 582440
rect 105538 582428 105544 582440
rect 105596 582428 105602 582480
rect 52362 582360 52368 582412
rect 52420 582400 52426 582412
rect 69934 582400 69940 582412
rect 52420 582372 69940 582400
rect 52420 582360 52426 582372
rect 69934 582360 69940 582372
rect 69992 582360 69998 582412
rect 76282 582360 76288 582412
rect 76340 582400 76346 582412
rect 87874 582400 87880 582412
rect 76340 582372 87880 582400
rect 76340 582360 76346 582372
rect 87874 582360 87880 582372
rect 87932 582360 87938 582412
rect 90266 582360 90272 582412
rect 90324 582400 90330 582412
rect 103514 582400 103520 582412
rect 90324 582372 103520 582400
rect 90324 582360 90330 582372
rect 103514 582360 103520 582372
rect 103572 582360 103578 582412
rect 87874 581612 87880 581664
rect 87932 581652 87938 581664
rect 108298 581652 108304 581664
rect 87932 581624 108304 581652
rect 87932 581612 87938 581624
rect 108298 581612 108304 581624
rect 108356 581612 108362 581664
rect 69658 581068 69664 581120
rect 69716 581108 69722 581120
rect 80238 581108 80244 581120
rect 69716 581080 80244 581108
rect 69716 581068 69722 581080
rect 80238 581068 80244 581080
rect 80296 581068 80302 581120
rect 50982 581000 50988 581052
rect 51040 581040 51046 581052
rect 90542 581040 90548 581052
rect 51040 581012 90548 581040
rect 51040 581000 51046 581012
rect 90542 581000 90548 581012
rect 90600 581000 90606 581052
rect 69658 580700 69664 580712
rect 64846 580672 69664 580700
rect 57882 580252 57888 580304
rect 57940 580292 57946 580304
rect 64846 580292 64874 580672
rect 69658 580660 69664 580672
rect 69716 580660 69722 580712
rect 85482 580660 85488 580712
rect 85540 580700 85546 580712
rect 85540 580672 93854 580700
rect 85540 580660 85546 580672
rect 57940 580264 64874 580292
rect 57940 580252 57946 580264
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 57882 579680 57888 579692
rect 3384 579652 57888 579680
rect 3384 579640 3390 579652
rect 57882 579640 57888 579652
rect 57940 579640 57946 579692
rect 64782 579640 64788 579692
rect 64840 579680 64846 579692
rect 66806 579680 66812 579692
rect 64840 579652 66812 579680
rect 64840 579640 64846 579652
rect 66806 579640 66812 579652
rect 66864 579640 66870 579692
rect 93826 579680 93854 580672
rect 94682 580456 94688 580508
rect 94740 580456 94746 580508
rect 94700 580304 94728 580456
rect 94682 580252 94688 580304
rect 94740 580252 94746 580304
rect 113450 579680 113456 579692
rect 93826 579652 113456 579680
rect 113450 579640 113456 579652
rect 113508 579640 113514 579692
rect 96890 578212 96896 578264
rect 96948 578252 96954 578264
rect 130378 578252 130384 578264
rect 96948 578224 130384 578252
rect 96948 578212 96954 578224
rect 130378 578212 130384 578224
rect 130436 578212 130442 578264
rect 102042 576920 102048 576972
rect 102100 576960 102106 576972
rect 118694 576960 118700 576972
rect 102100 576932 118700 576960
rect 102100 576920 102106 576932
rect 118694 576920 118700 576932
rect 118752 576920 118758 576972
rect 97074 576852 97080 576904
rect 97132 576892 97138 576904
rect 128354 576892 128360 576904
rect 97132 576864 128360 576892
rect 97132 576852 97138 576864
rect 128354 576852 128360 576864
rect 128412 576852 128418 576904
rect 97902 576716 97908 576768
rect 97960 576756 97966 576768
rect 102042 576756 102048 576768
rect 97960 576728 102048 576756
rect 97960 576716 97966 576728
rect 102042 576716 102048 576728
rect 102100 576716 102106 576768
rect 21358 576104 21364 576156
rect 21416 576144 21422 576156
rect 31754 576144 31760 576156
rect 21416 576116 31760 576144
rect 21416 576104 21422 576116
rect 31754 576104 31760 576116
rect 31812 576104 31818 576156
rect 31754 575492 31760 575544
rect 31812 575532 31818 575544
rect 33042 575532 33048 575544
rect 31812 575504 33048 575532
rect 31812 575492 31818 575504
rect 33042 575492 33048 575504
rect 33100 575532 33106 575544
rect 66530 575532 66536 575544
rect 33100 575504 66536 575532
rect 33100 575492 33106 575504
rect 66530 575492 66536 575504
rect 66588 575492 66594 575544
rect 94774 574744 94780 574796
rect 94832 574784 94838 574796
rect 120074 574784 120080 574796
rect 94832 574756 120080 574784
rect 94832 574744 94838 574756
rect 120074 574744 120080 574756
rect 120132 574744 120138 574796
rect 96246 574064 96252 574116
rect 96304 574104 96310 574116
rect 105630 574104 105636 574116
rect 96304 574076 105636 574104
rect 96304 574064 96310 574076
rect 105630 574064 105636 574076
rect 105688 574064 105694 574116
rect 56502 571956 56508 572008
rect 56560 571996 56566 572008
rect 66438 571996 66444 572008
rect 56560 571968 66444 571996
rect 56560 571956 56566 571968
rect 66438 571956 66444 571968
rect 66496 571956 66502 572008
rect 64690 571344 64696 571396
rect 64748 571384 64754 571396
rect 66714 571384 66720 571396
rect 64748 571356 66720 571384
rect 64748 571344 64754 571356
rect 66714 571344 66720 571356
rect 66772 571344 66778 571396
rect 107562 570596 107568 570648
rect 107620 570636 107626 570648
rect 582742 570636 582748 570648
rect 107620 570608 582748 570636
rect 107620 570596 107626 570608
rect 582742 570596 582748 570608
rect 582800 570596 582806 570648
rect 97902 569916 97908 569968
rect 97960 569956 97966 569968
rect 107562 569956 107568 569968
rect 97960 569928 107568 569956
rect 97960 569916 97966 569928
rect 107562 569916 107568 569928
rect 107620 569916 107626 569968
rect 97902 569168 97908 569220
rect 97960 569208 97966 569220
rect 133874 569208 133880 569220
rect 97960 569180 133880 569208
rect 97960 569168 97966 569180
rect 133874 569168 133880 569180
rect 133932 569168 133938 569220
rect 3418 568488 3424 568540
rect 3476 568528 3482 568540
rect 4798 568528 4804 568540
rect 3476 568500 4804 568528
rect 3476 568488 3482 568500
rect 4798 568488 4804 568500
rect 4856 568488 4862 568540
rect 60642 567196 60648 567248
rect 60700 567236 60706 567248
rect 66990 567236 66996 567248
rect 60700 567208 66996 567236
rect 60700 567196 60706 567208
rect 66990 567196 66996 567208
rect 67048 567196 67054 567248
rect 52270 565836 52276 565888
rect 52328 565876 52334 565888
rect 67634 565876 67640 565888
rect 52328 565848 67640 565876
rect 52328 565836 52334 565848
rect 67634 565836 67640 565848
rect 67692 565836 67698 565888
rect 41322 564408 41328 564460
rect 41380 564448 41386 564460
rect 66714 564448 66720 564460
rect 41380 564420 66720 564448
rect 41380 564408 41386 564420
rect 66714 564408 66720 564420
rect 66772 564408 66778 564460
rect 57790 564340 57796 564392
rect 57848 564380 57854 564392
rect 66438 564380 66444 564392
rect 57848 564352 66444 564380
rect 57848 564340 57854 564352
rect 66438 564340 66444 564352
rect 66496 564340 66502 564392
rect 48130 563660 48136 563712
rect 48188 563700 48194 563712
rect 57790 563700 57796 563712
rect 48188 563672 57796 563700
rect 48188 563660 48194 563672
rect 57790 563660 57796 563672
rect 57848 563660 57854 563712
rect 50890 560260 50896 560312
rect 50948 560300 50954 560312
rect 66990 560300 66996 560312
rect 50948 560272 66996 560300
rect 50948 560260 50954 560272
rect 66990 560260 66996 560272
rect 67048 560260 67054 560312
rect 59170 558900 59176 558952
rect 59228 558940 59234 558952
rect 66990 558940 66996 558952
rect 59228 558912 66996 558940
rect 59228 558900 59234 558912
rect 66990 558900 66996 558912
rect 67048 558900 67054 558952
rect 97258 558152 97264 558204
rect 97316 558192 97322 558204
rect 115198 558192 115204 558204
rect 97316 558164 115204 558192
rect 97316 558152 97322 558164
rect 115198 558152 115204 558164
rect 115256 558152 115262 558204
rect 53742 557540 53748 557592
rect 53800 557580 53806 557592
rect 66990 557580 66996 557592
rect 53800 557552 66996 557580
rect 53800 557540 53806 557552
rect 66990 557540 66996 557552
rect 67048 557540 67054 557592
rect 97350 555432 97356 555484
rect 97408 555472 97414 555484
rect 121546 555472 121552 555484
rect 97408 555444 121552 555472
rect 97408 555432 97414 555444
rect 121546 555432 121552 555444
rect 121604 555432 121610 555484
rect 63310 554752 63316 554804
rect 63368 554792 63374 554804
rect 66990 554792 66996 554804
rect 63368 554764 66996 554792
rect 63368 554752 63374 554764
rect 66990 554752 66996 554764
rect 67048 554752 67054 554804
rect 3510 553800 3516 553852
rect 3568 553840 3574 553852
rect 7558 553840 7564 553852
rect 3568 553812 7564 553840
rect 3568 553800 3574 553812
rect 7558 553800 7564 553812
rect 7616 553800 7622 553852
rect 57790 553392 57796 553444
rect 57848 553432 57854 553444
rect 66990 553432 66996 553444
rect 57848 553404 66996 553432
rect 57848 553392 57854 553404
rect 66990 553392 66996 553404
rect 67048 553392 67054 553444
rect 96982 552032 96988 552084
rect 97040 552072 97046 552084
rect 109678 552072 109684 552084
rect 97040 552044 109684 552072
rect 97040 552032 97046 552044
rect 109678 552032 109684 552044
rect 109736 552032 109742 552084
rect 96798 551896 96804 551948
rect 96856 551896 96862 551948
rect 96816 551744 96844 551896
rect 96798 551692 96804 551744
rect 96856 551692 96862 551744
rect 97902 550604 97908 550656
rect 97960 550644 97966 550656
rect 115934 550644 115940 550656
rect 97960 550616 115940 550644
rect 97960 550604 97966 550616
rect 115934 550604 115940 550616
rect 115992 550604 115998 550656
rect 48038 549244 48044 549296
rect 48096 549284 48102 549296
rect 66530 549284 66536 549296
rect 48096 549256 66536 549284
rect 48096 549244 48102 549256
rect 66530 549244 66536 549256
rect 66588 549244 66594 549296
rect 53466 546456 53472 546508
rect 53524 546496 53530 546508
rect 66990 546496 66996 546508
rect 53524 546468 66996 546496
rect 53524 546456 53530 546468
rect 66990 546456 66996 546468
rect 67048 546456 67054 546508
rect 95142 546456 95148 546508
rect 95200 546496 95206 546508
rect 96706 546496 96712 546508
rect 95200 546468 96712 546496
rect 95200 546456 95206 546468
rect 96706 546456 96712 546468
rect 96764 546456 96770 546508
rect 54938 544348 54944 544400
rect 54996 544388 55002 544400
rect 61930 544388 61936 544400
rect 54996 544360 61936 544388
rect 54996 544348 55002 544360
rect 61930 544348 61936 544360
rect 61988 544388 61994 544400
rect 66714 544388 66720 544400
rect 61988 544360 66720 544388
rect 61988 544348 61994 544360
rect 66714 544348 66720 544360
rect 66772 544348 66778 544400
rect 97534 543736 97540 543788
rect 97592 543776 97598 543788
rect 108390 543776 108396 543788
rect 97592 543748 108396 543776
rect 97592 543736 97598 543748
rect 108390 543736 108396 543748
rect 108448 543736 108454 543788
rect 3418 540200 3424 540252
rect 3476 540240 3482 540252
rect 34514 540240 34520 540252
rect 3476 540212 34520 540240
rect 3476 540200 3482 540212
rect 34514 540200 34520 540212
rect 34572 540200 34578 540252
rect 67726 539792 67732 539844
rect 67784 539832 67790 539844
rect 71774 539832 71780 539844
rect 67784 539804 71780 539832
rect 67784 539792 67790 539804
rect 71774 539792 71780 539804
rect 71832 539792 71838 539844
rect 93210 539792 93216 539844
rect 93268 539832 93274 539844
rect 94682 539832 94688 539844
rect 93268 539804 94688 539832
rect 93268 539792 93274 539804
rect 94682 539792 94688 539804
rect 94740 539792 94746 539844
rect 70302 539656 70308 539708
rect 70360 539696 70366 539708
rect 72326 539696 72332 539708
rect 70360 539668 72332 539696
rect 70360 539656 70366 539668
rect 72326 539656 72332 539668
rect 72384 539656 72390 539708
rect 34514 539588 34520 539640
rect 34572 539628 34578 539640
rect 35710 539628 35716 539640
rect 34572 539600 35716 539628
rect 34572 539588 34578 539600
rect 35710 539588 35716 539600
rect 35768 539628 35774 539640
rect 61286 539628 61292 539640
rect 35768 539600 61292 539628
rect 35768 539588 35774 539600
rect 61286 539588 61292 539600
rect 61344 539588 61350 539640
rect 67818 539520 67824 539572
rect 67876 539560 67882 539572
rect 68922 539560 68928 539572
rect 67876 539532 68928 539560
rect 67876 539520 67882 539532
rect 68922 539520 68928 539532
rect 68980 539520 68986 539572
rect 68922 538840 68928 538892
rect 68980 538880 68986 538892
rect 82906 538880 82912 538892
rect 68980 538852 82912 538880
rect 68980 538840 68986 538852
rect 82906 538840 82912 538852
rect 82964 538840 82970 538892
rect 88242 538296 88248 538348
rect 88300 538336 88306 538348
rect 95418 538336 95424 538348
rect 88300 538308 95424 538336
rect 88300 538296 88306 538308
rect 95418 538296 95424 538308
rect 95476 538296 95482 538348
rect 15838 538228 15844 538280
rect 15896 538268 15902 538280
rect 93946 538268 93952 538280
rect 15896 538240 93952 538268
rect 15896 538228 15902 538240
rect 93946 538228 93952 538240
rect 94004 538228 94010 538280
rect 7558 538160 7564 538212
rect 7616 538200 7622 538212
rect 70670 538200 70676 538212
rect 7616 538172 70676 538200
rect 7616 538160 7622 538172
rect 70670 538160 70676 538172
rect 70728 538160 70734 538212
rect 90358 538160 90364 538212
rect 90416 538200 90422 538212
rect 136634 538200 136640 538212
rect 90416 538172 136640 538200
rect 90416 538160 90422 538172
rect 136634 538160 136640 538172
rect 136692 538160 136698 538212
rect 61838 537480 61844 537532
rect 61896 537520 61902 537532
rect 96890 537520 96896 537532
rect 61896 537492 96896 537520
rect 61896 537480 61902 537492
rect 96890 537480 96896 537492
rect 96948 537480 96954 537532
rect 70670 536800 70676 536852
rect 70728 536840 70734 536852
rect 71130 536840 71136 536852
rect 70728 536812 71136 536840
rect 70728 536800 70734 536812
rect 71130 536800 71136 536812
rect 71188 536800 71194 536852
rect 43438 536732 43444 536784
rect 43496 536772 43502 536784
rect 73430 536772 73436 536784
rect 43496 536744 73436 536772
rect 43496 536732 43502 536744
rect 73430 536732 73436 536744
rect 73488 536732 73494 536784
rect 86862 536732 86868 536784
rect 86920 536772 86926 536784
rect 119338 536772 119344 536784
rect 86920 536744 119344 536772
rect 86920 536732 86926 536744
rect 119338 536732 119344 536744
rect 119396 536732 119402 536784
rect 61286 536664 61292 536716
rect 61344 536704 61350 536716
rect 69382 536704 69388 536716
rect 61344 536676 69388 536704
rect 61344 536664 61350 536676
rect 69382 536664 69388 536676
rect 69440 536664 69446 536716
rect 73430 535712 73436 535764
rect 73488 535752 73494 535764
rect 76558 535752 76564 535764
rect 73488 535724 76564 535752
rect 73488 535712 73494 535724
rect 76558 535712 76564 535724
rect 76616 535712 76622 535764
rect 72786 535440 72792 535492
rect 72844 535480 72850 535492
rect 73798 535480 73804 535492
rect 72844 535452 73804 535480
rect 72844 535440 72850 535452
rect 73798 535440 73804 535452
rect 73856 535440 73862 535492
rect 91002 535440 91008 535492
rect 91060 535480 91066 535492
rect 92750 535480 92756 535492
rect 91060 535452 92756 535480
rect 91060 535440 91066 535452
rect 92750 535440 92756 535452
rect 92808 535440 92814 535492
rect 3418 534692 3424 534744
rect 3476 534732 3482 534744
rect 94498 534732 94504 534744
rect 3476 534704 94504 534732
rect 3476 534692 3482 534704
rect 94498 534692 94504 534704
rect 94556 534692 94562 534744
rect 49510 533400 49516 533452
rect 49568 533440 49574 533452
rect 84286 533440 84292 533452
rect 49568 533412 84292 533440
rect 49568 533400 49574 533412
rect 84286 533400 84292 533412
rect 84344 533400 84350 533452
rect 88334 533400 88340 533452
rect 88392 533440 88398 533452
rect 88886 533440 88892 533452
rect 88392 533412 88892 533440
rect 88392 533400 88398 533412
rect 88886 533400 88892 533412
rect 88944 533400 88950 533452
rect 80054 533332 80060 533384
rect 80112 533372 80118 533384
rect 80606 533372 80612 533384
rect 80112 533344 80612 533372
rect 80112 533332 80118 533344
rect 80606 533332 80612 533344
rect 80664 533332 80670 533384
rect 84010 533332 84016 533384
rect 84068 533372 84074 533384
rect 136634 533372 136640 533384
rect 84068 533344 136640 533372
rect 84068 533332 84074 533344
rect 136634 533332 136640 533344
rect 136692 533332 136698 533384
rect 59998 531972 60004 532024
rect 60056 532012 60062 532024
rect 98086 532012 98092 532024
rect 60056 531984 98092 532012
rect 60056 531972 60062 531984
rect 98086 531972 98092 531984
rect 98144 531972 98150 532024
rect 65978 529184 65984 529236
rect 66036 529224 66042 529236
rect 117314 529224 117320 529236
rect 66036 529196 117320 529224
rect 66036 529184 66042 529196
rect 117314 529184 117320 529196
rect 117372 529184 117378 529236
rect 3510 527824 3516 527876
rect 3568 527864 3574 527876
rect 128354 527864 128360 527876
rect 3568 527836 128360 527864
rect 3568 527824 3574 527836
rect 128354 527824 128360 527836
rect 128412 527824 128418 527876
rect 75178 526396 75184 526448
rect 75236 526436 75242 526448
rect 96798 526436 96804 526448
rect 75236 526408 96804 526436
rect 75236 526396 75242 526408
rect 96798 526396 96804 526408
rect 96856 526396 96862 526448
rect 109678 521568 109684 521620
rect 109736 521608 109742 521620
rect 111794 521608 111800 521620
rect 109736 521580 111800 521608
rect 109736 521568 109742 521580
rect 111794 521568 111800 521580
rect 111852 521568 111858 521620
rect 71038 520888 71044 520940
rect 71096 520928 71102 520940
rect 91186 520928 91192 520940
rect 71096 520900 91192 520928
rect 71096 520888 71102 520900
rect 91186 520888 91192 520900
rect 91244 520888 91250 520940
rect 55030 518168 55036 518220
rect 55088 518208 55094 518220
rect 97994 518208 98000 518220
rect 55088 518180 98000 518208
rect 55088 518168 55094 518180
rect 97994 518168 98000 518180
rect 98052 518168 98058 518220
rect 3510 514768 3516 514820
rect 3568 514808 3574 514820
rect 40678 514808 40684 514820
rect 3568 514780 40684 514808
rect 3568 514768 3574 514780
rect 40678 514768 40684 514780
rect 40736 514768 40742 514820
rect 50890 511232 50896 511284
rect 50948 511272 50954 511284
rect 580166 511272 580172 511284
rect 50948 511244 580172 511272
rect 50948 511232 50954 511244
rect 580166 511232 580172 511244
rect 580224 511232 580230 511284
rect 63310 490560 63316 490612
rect 63368 490600 63374 490612
rect 128446 490600 128452 490612
rect 63368 490572 128452 490600
rect 63368 490560 63374 490572
rect 128446 490560 128452 490572
rect 128504 490560 128510 490612
rect 80146 487772 80152 487824
rect 80204 487812 80210 487824
rect 129734 487812 129740 487824
rect 80204 487784 129740 487812
rect 80204 487772 80210 487784
rect 129734 487772 129740 487784
rect 129792 487772 129798 487824
rect 71130 485052 71136 485104
rect 71188 485092 71194 485104
rect 122926 485092 122932 485104
rect 71188 485064 122932 485092
rect 71188 485052 71194 485064
rect 122926 485052 122932 485064
rect 122984 485052 122990 485104
rect 66070 482264 66076 482316
rect 66128 482304 66134 482316
rect 118786 482304 118792 482316
rect 66128 482276 118792 482304
rect 66128 482264 66134 482276
rect 118786 482264 118792 482276
rect 118844 482264 118850 482316
rect 3418 478116 3424 478168
rect 3476 478156 3482 478168
rect 15838 478156 15844 478168
rect 3476 478128 15844 478156
rect 3476 478116 3482 478128
rect 15838 478116 15844 478128
rect 15896 478116 15902 478168
rect 67726 478116 67732 478168
rect 67784 478156 67790 478168
rect 98730 478156 98736 478168
rect 67784 478128 98736 478156
rect 67784 478116 67790 478128
rect 98730 478116 98736 478128
rect 98788 478116 98794 478168
rect 85482 475124 85488 475176
rect 85540 475164 85546 475176
rect 93210 475164 93216 475176
rect 85540 475136 93216 475164
rect 85540 475124 85546 475136
rect 93210 475124 93216 475136
rect 93268 475124 93274 475176
rect 77202 473288 77208 473340
rect 77260 473328 77266 473340
rect 77938 473328 77944 473340
rect 77260 473300 77944 473328
rect 77260 473288 77266 473300
rect 77938 473288 77944 473300
rect 77996 473288 78002 473340
rect 73798 472608 73804 472660
rect 73856 472648 73862 472660
rect 116118 472648 116124 472660
rect 73856 472620 116124 472648
rect 73856 472608 73862 472620
rect 116118 472608 116124 472620
rect 116176 472608 116182 472660
rect 82814 467100 82820 467152
rect 82872 467140 82878 467152
rect 109034 467140 109040 467152
rect 82872 467112 109040 467140
rect 82872 467100 82878 467112
rect 109034 467100 109040 467112
rect 109092 467100 109098 467152
rect 65978 466420 65984 466472
rect 66036 466460 66042 466472
rect 70486 466460 70492 466472
rect 66036 466432 70492 466460
rect 66036 466420 66042 466432
rect 70486 466420 70492 466432
rect 70544 466420 70550 466472
rect 86310 464312 86316 464364
rect 86368 464352 86374 464364
rect 95234 464352 95240 464364
rect 86368 464324 95240 464352
rect 86368 464312 86374 464324
rect 95234 464312 95240 464324
rect 95292 464312 95298 464364
rect 85574 462952 85580 463004
rect 85632 462992 85638 463004
rect 120166 462992 120172 463004
rect 85632 462964 120172 462992
rect 85632 462952 85638 462964
rect 120166 462952 120172 462964
rect 120224 462952 120230 463004
rect 3510 462340 3516 462392
rect 3568 462380 3574 462392
rect 14458 462380 14464 462392
rect 3568 462352 14464 462380
rect 3568 462340 3574 462352
rect 14458 462340 14464 462352
rect 14516 462340 14522 462392
rect 67726 460164 67732 460216
rect 67784 460204 67790 460216
rect 96706 460204 96712 460216
rect 67784 460176 96712 460204
rect 67784 460164 67790 460176
rect 96706 460164 96712 460176
rect 96764 460164 96770 460216
rect 64782 458804 64788 458856
rect 64840 458844 64846 458856
rect 92566 458844 92572 458856
rect 64840 458816 92572 458844
rect 64840 458804 64846 458816
rect 92566 458804 92572 458816
rect 92624 458804 92630 458856
rect 86862 457512 86868 457564
rect 86920 457552 86926 457564
rect 104342 457552 104348 457564
rect 86920 457524 104348 457552
rect 86920 457512 86926 457524
rect 104342 457512 104348 457524
rect 104400 457512 104406 457564
rect 64598 457444 64604 457496
rect 64656 457484 64662 457496
rect 86954 457484 86960 457496
rect 64656 457456 86960 457484
rect 64656 457444 64662 457456
rect 86954 457444 86960 457456
rect 87012 457444 87018 457496
rect 64690 454656 64696 454708
rect 64748 454696 64754 454708
rect 106918 454696 106924 454708
rect 64748 454668 106924 454696
rect 64748 454656 64754 454668
rect 106918 454656 106924 454668
rect 106976 454656 106982 454708
rect 60642 453296 60648 453348
rect 60700 453336 60706 453348
rect 123110 453336 123116 453348
rect 60700 453308 123116 453336
rect 60700 453296 60706 453308
rect 123110 453296 123116 453308
rect 123168 453296 123174 453348
rect 79318 451868 79324 451920
rect 79376 451908 79382 451920
rect 90358 451908 90364 451920
rect 79376 451880 90364 451908
rect 79376 451868 79382 451880
rect 90358 451868 90364 451880
rect 90416 451868 90422 451920
rect 68922 449896 68928 449948
rect 68980 449936 68986 449948
rect 80054 449936 80060 449948
rect 68980 449908 80060 449936
rect 68980 449896 68986 449908
rect 80054 449896 80060 449908
rect 80112 449896 80118 449948
rect 78674 449216 78680 449268
rect 78732 449256 78738 449268
rect 101490 449256 101496 449268
rect 78732 449228 101496 449256
rect 78732 449216 78738 449228
rect 101490 449216 101496 449228
rect 101548 449216 101554 449268
rect 53742 449148 53748 449200
rect 53800 449188 53806 449200
rect 85666 449188 85672 449200
rect 53800 449160 85672 449188
rect 53800 449148 53806 449160
rect 85666 449148 85672 449160
rect 85724 449148 85730 449200
rect 101398 449148 101404 449200
rect 101456 449188 101462 449200
rect 117498 449188 117504 449200
rect 101456 449160 117504 449188
rect 101456 449148 101462 449160
rect 117498 449148 117504 449160
rect 117556 449148 117562 449200
rect 3142 448536 3148 448588
rect 3200 448576 3206 448588
rect 36538 448576 36544 448588
rect 3200 448548 36544 448576
rect 3200 448536 3206 448548
rect 36538 448536 36544 448548
rect 36596 448536 36602 448588
rect 78030 447856 78036 447908
rect 78088 447896 78094 447908
rect 91094 447896 91100 447908
rect 78088 447868 91100 447896
rect 78088 447856 78094 447868
rect 91094 447856 91100 447868
rect 91152 447856 91158 447908
rect 88334 447788 88340 447840
rect 88392 447828 88398 447840
rect 113266 447828 113272 447840
rect 88392 447800 113272 447828
rect 88392 447788 88398 447800
rect 113266 447788 113272 447800
rect 113324 447788 113330 447840
rect 91002 446428 91008 446480
rect 91060 446468 91066 446480
rect 118878 446468 118884 446480
rect 91060 446440 118884 446468
rect 91060 446428 91066 446440
rect 118878 446428 118884 446440
rect 118936 446428 118942 446480
rect 52362 446360 52368 446412
rect 52420 446400 52426 446412
rect 95970 446400 95976 446412
rect 52420 446372 95976 446400
rect 52420 446360 52426 446372
rect 95970 446360 95976 446372
rect 96028 446360 96034 446412
rect 95878 444388 95884 444440
rect 95936 444428 95942 444440
rect 96522 444428 96528 444440
rect 95936 444400 96528 444428
rect 95936 444388 95942 444400
rect 96522 444388 96528 444400
rect 96580 444428 96586 444440
rect 116026 444428 116032 444440
rect 96580 444400 116032 444428
rect 96580 444388 96586 444400
rect 116026 444388 116032 444400
rect 116084 444388 116090 444440
rect 81434 443708 81440 443760
rect 81492 443748 81498 443760
rect 96522 443748 96528 443760
rect 81492 443720 96528 443748
rect 81492 443708 81498 443720
rect 96522 443708 96528 443720
rect 96580 443708 96586 443760
rect 48130 443640 48136 443692
rect 48188 443680 48194 443692
rect 88426 443680 88432 443692
rect 48188 443652 88432 443680
rect 48188 443640 48194 443652
rect 88426 443640 88432 443652
rect 88484 443640 88490 443692
rect 100018 443640 100024 443692
rect 100076 443680 100082 443692
rect 115290 443680 115296 443692
rect 100076 443652 115296 443680
rect 100076 443640 100082 443652
rect 115290 443640 115296 443652
rect 115348 443640 115354 443692
rect 93854 442960 93860 443012
rect 93912 443000 93918 443012
rect 95142 443000 95148 443012
rect 93912 442972 95148 443000
rect 93912 442960 93918 442972
rect 95142 442960 95148 442972
rect 95200 443000 95206 443012
rect 124306 443000 124312 443012
rect 95200 442972 124312 443000
rect 95200 442960 95206 442972
rect 124306 442960 124312 442972
rect 124364 442960 124370 443012
rect 40678 442892 40684 442944
rect 40736 442932 40742 442944
rect 103514 442932 103520 442944
rect 40736 442904 103520 442932
rect 40736 442892 40742 442904
rect 103514 442892 103520 442904
rect 103572 442892 103578 442944
rect 115198 442892 115204 442944
rect 115256 442932 115262 442944
rect 120258 442932 120264 442944
rect 115256 442904 120264 442932
rect 115256 442892 115262 442904
rect 120258 442892 120264 442904
rect 120316 442892 120322 442944
rect 106274 442280 106280 442332
rect 106332 442320 106338 442332
rect 106918 442320 106924 442332
rect 106332 442292 106924 442320
rect 106332 442280 106338 442292
rect 106918 442280 106924 442292
rect 106976 442280 106982 442332
rect 77294 442212 77300 442264
rect 77352 442252 77358 442264
rect 113358 442252 113364 442264
rect 77352 442224 113364 442252
rect 77352 442212 77358 442224
rect 113358 442212 113364 442224
rect 113416 442212 113422 442264
rect 106274 441600 106280 441652
rect 106332 441640 106338 441652
rect 131114 441640 131120 441652
rect 106332 441612 131120 441640
rect 106332 441600 106338 441612
rect 131114 441600 131120 441612
rect 131172 441600 131178 441652
rect 54938 440920 54944 440972
rect 54996 440960 55002 440972
rect 78398 440960 78404 440972
rect 54996 440932 78404 440960
rect 54996 440920 55002 440932
rect 78398 440920 78404 440932
rect 78456 440920 78462 440972
rect 67634 440852 67640 440904
rect 67692 440892 67698 440904
rect 114554 440892 114560 440904
rect 67692 440864 114560 440892
rect 67692 440852 67698 440864
rect 114554 440852 114560 440864
rect 114612 440852 114618 440904
rect 102594 438948 102600 439000
rect 102652 438988 102658 439000
rect 102778 438988 102784 439000
rect 102652 438960 102784 438988
rect 102652 438948 102658 438960
rect 102778 438948 102784 438960
rect 102836 438988 102842 439000
rect 127066 438988 127072 439000
rect 102836 438960 127072 438988
rect 102836 438948 102842 438960
rect 127066 438948 127072 438960
rect 127124 438948 127130 439000
rect 108114 438880 108120 438932
rect 108172 438920 108178 438932
rect 108390 438920 108396 438932
rect 108172 438892 108396 438920
rect 108172 438880 108178 438892
rect 108390 438880 108396 438892
rect 108448 438920 108454 438932
rect 137278 438920 137284 438932
rect 108448 438892 137284 438920
rect 108448 438880 108454 438892
rect 137278 438880 137284 438892
rect 137336 438880 137342 438932
rect 50890 438132 50896 438184
rect 50948 438172 50954 438184
rect 74718 438172 74724 438184
rect 50948 438144 74724 438172
rect 50948 438132 50954 438144
rect 74718 438132 74724 438144
rect 74776 438132 74782 438184
rect 122190 438132 122196 438184
rect 122248 438172 122254 438184
rect 583110 438172 583116 438184
rect 122248 438144 583116 438172
rect 122248 438132 122254 438144
rect 583110 438132 583116 438144
rect 583168 438132 583174 438184
rect 108298 437520 108304 437572
rect 108356 437560 108362 437572
rect 125594 437560 125600 437572
rect 108356 437532 125600 437560
rect 108356 437520 108362 437532
rect 125594 437520 125600 437532
rect 125652 437520 125658 437572
rect 95970 437452 95976 437504
rect 96028 437492 96034 437504
rect 122190 437492 122196 437504
rect 96028 437464 122196 437492
rect 96028 437452 96034 437464
rect 122190 437452 122196 437464
rect 122248 437452 122254 437504
rect 71130 437384 71136 437436
rect 71188 437424 71194 437436
rect 75178 437424 75184 437436
rect 71188 437396 75184 437424
rect 71188 437384 71194 437396
rect 75178 437384 75184 437396
rect 75236 437384 75242 437436
rect 57698 436160 57704 436212
rect 57756 436200 57762 436212
rect 73982 436200 73988 436212
rect 57756 436172 73988 436200
rect 57756 436160 57762 436172
rect 73982 436160 73988 436172
rect 74040 436160 74046 436212
rect 77938 436160 77944 436212
rect 77996 436200 78002 436212
rect 82906 436200 82912 436212
rect 77996 436172 82912 436200
rect 77996 436160 78002 436172
rect 82906 436160 82912 436172
rect 82964 436160 82970 436212
rect 123018 436200 123024 436212
rect 109006 436172 123024 436200
rect 33778 436092 33784 436144
rect 33836 436132 33842 436144
rect 71130 436132 71136 436144
rect 33836 436104 71136 436132
rect 33836 436092 33842 436104
rect 71130 436092 71136 436104
rect 71188 436092 71194 436144
rect 76834 436092 76840 436144
rect 76892 436132 76898 436144
rect 79318 436132 79324 436144
rect 76892 436104 79324 436132
rect 76892 436092 76898 436104
rect 79318 436092 79324 436104
rect 79376 436092 79382 436144
rect 98730 436092 98736 436144
rect 98788 436132 98794 436144
rect 99926 436132 99932 436144
rect 98788 436104 99932 436132
rect 98788 436092 98794 436104
rect 99926 436092 99932 436104
rect 99984 436092 99990 436144
rect 101490 436092 101496 436144
rect 101548 436132 101554 436144
rect 103698 436132 103704 436144
rect 101548 436104 103704 436132
rect 101548 436092 101554 436104
rect 103698 436092 103704 436104
rect 103756 436132 103762 436144
rect 109006 436132 109034 436172
rect 123018 436160 123024 436172
rect 123076 436160 123082 436212
rect 103756 436104 109034 436132
rect 103756 436092 103762 436104
rect 111058 436092 111064 436144
rect 111116 436132 111122 436144
rect 140866 436132 140872 436144
rect 111116 436104 140872 436132
rect 111116 436092 111122 436104
rect 140866 436092 140872 436104
rect 140924 436092 140930 436144
rect 68462 435344 68468 435396
rect 68520 435384 68526 435396
rect 71774 435384 71780 435396
rect 68520 435356 71780 435384
rect 68520 435344 68526 435356
rect 71774 435344 71780 435356
rect 71832 435384 71838 435396
rect 72694 435384 72700 435396
rect 71832 435356 72700 435384
rect 71832 435344 71838 435356
rect 72694 435344 72700 435356
rect 72752 435344 72758 435396
rect 72602 434800 72608 434852
rect 72660 434840 72666 434852
rect 132494 434840 132500 434852
rect 72660 434812 132500 434840
rect 72660 434800 72666 434812
rect 132494 434800 132500 434812
rect 132552 434800 132558 434852
rect 4798 434732 4804 434784
rect 4856 434772 4862 434784
rect 111794 434772 111800 434784
rect 4856 434744 111800 434772
rect 4856 434732 4862 434744
rect 111794 434732 111800 434744
rect 111852 434772 111858 434784
rect 112438 434772 112444 434784
rect 111852 434744 112444 434772
rect 111852 434732 111858 434744
rect 112438 434732 112444 434744
rect 112496 434772 112502 434784
rect 117406 434772 117412 434784
rect 112496 434744 117412 434772
rect 112496 434732 112502 434744
rect 117406 434732 117412 434744
rect 117464 434732 117470 434784
rect 67358 433984 67364 434036
rect 67416 434024 67422 434036
rect 74534 434024 74540 434036
rect 67416 433996 74540 434024
rect 67416 433984 67422 433996
rect 74534 433984 74540 433996
rect 74592 433984 74598 434036
rect 105906 433984 105912 434036
rect 105964 434024 105970 434036
rect 118970 434024 118976 434036
rect 105964 433996 118976 434024
rect 105964 433984 105970 433996
rect 118970 433984 118976 433996
rect 119028 433984 119034 434036
rect 68370 433712 68376 433764
rect 68428 433752 68434 433764
rect 71222 433752 71228 433764
rect 68428 433724 71228 433752
rect 68428 433712 68434 433724
rect 71222 433712 71228 433724
rect 71280 433712 71286 433764
rect 68646 433644 68652 433696
rect 68704 433684 68710 433696
rect 69198 433684 69204 433696
rect 68704 433656 69204 433684
rect 68704 433644 68710 433656
rect 69198 433644 69204 433656
rect 69256 433644 69262 433696
rect 110874 433644 110880 433696
rect 110932 433644 110938 433696
rect 61746 433304 61752 433356
rect 61804 433344 61810 433356
rect 63402 433344 63408 433356
rect 61804 433316 63408 433344
rect 61804 433304 61810 433316
rect 63402 433304 63408 433316
rect 63460 433344 63466 433356
rect 66254 433344 66260 433356
rect 63460 433316 66260 433344
rect 63460 433304 63466 433316
rect 66254 433304 66260 433316
rect 66312 433304 66318 433356
rect 110892 433276 110920 433644
rect 112714 433276 112720 433288
rect 110892 433248 112720 433276
rect 112714 433236 112720 433248
rect 112772 433236 112778 433288
rect 112714 432012 112720 432064
rect 112772 432052 112778 432064
rect 117590 432052 117596 432064
rect 112772 432024 117596 432052
rect 112772 432012 112778 432024
rect 117590 432012 117596 432024
rect 117648 432012 117654 432064
rect 59078 431944 59084 431996
rect 59136 431984 59142 431996
rect 66438 431984 66444 431996
rect 59136 431956 66444 431984
rect 59136 431944 59142 431956
rect 66438 431944 66444 431956
rect 66496 431944 66502 431996
rect 115566 431944 115572 431996
rect 115624 431984 115630 431996
rect 133966 431984 133972 431996
rect 115624 431956 133972 431984
rect 115624 431944 115630 431956
rect 133966 431944 133972 431956
rect 134024 431944 134030 431996
rect 60550 430584 60556 430636
rect 60608 430624 60614 430636
rect 66714 430624 66720 430636
rect 60608 430596 66720 430624
rect 60608 430584 60614 430596
rect 66714 430584 66720 430596
rect 66772 430584 66778 430636
rect 115842 430584 115848 430636
rect 115900 430624 115906 430636
rect 135898 430624 135904 430636
rect 115900 430596 135904 430624
rect 115900 430584 115906 430596
rect 135898 430584 135904 430596
rect 135956 430584 135962 430636
rect 115750 430516 115756 430568
rect 115808 430556 115814 430568
rect 136634 430556 136640 430568
rect 115808 430528 136640 430556
rect 115808 430516 115814 430528
rect 136634 430516 136640 430528
rect 136692 430556 136698 430568
rect 142798 430556 142804 430568
rect 136692 430528 142804 430556
rect 136692 430516 136698 430528
rect 142798 430516 142804 430528
rect 142856 430516 142862 430568
rect 52362 429224 52368 429276
rect 52420 429264 52426 429276
rect 66714 429264 66720 429276
rect 52420 429236 66720 429264
rect 52420 429224 52426 429236
rect 66714 429224 66720 429236
rect 66772 429224 66778 429276
rect 115842 429088 115848 429140
rect 115900 429128 115906 429140
rect 118786 429128 118792 429140
rect 115900 429100 118792 429128
rect 115900 429088 115906 429100
rect 118786 429088 118792 429100
rect 118844 429128 118850 429140
rect 124858 429128 124864 429140
rect 118844 429100 124864 429128
rect 118844 429088 118850 429100
rect 124858 429088 124864 429100
rect 124916 429088 124922 429140
rect 60642 427796 60648 427848
rect 60700 427836 60706 427848
rect 66714 427836 66720 427848
rect 60700 427808 66720 427836
rect 60700 427796 60706 427808
rect 66714 427796 66720 427808
rect 66772 427796 66778 427848
rect 53742 426436 53748 426488
rect 53800 426476 53806 426488
rect 66714 426476 66720 426488
rect 53800 426448 66720 426476
rect 53800 426436 53806 426448
rect 66714 426436 66720 426448
rect 66772 426436 66778 426488
rect 118786 426368 118792 426420
rect 118844 426408 118850 426420
rect 122834 426408 122840 426420
rect 118844 426380 122840 426408
rect 118844 426368 118850 426380
rect 122834 426368 122840 426380
rect 122892 426368 122898 426420
rect 50890 425688 50896 425740
rect 50948 425728 50954 425740
rect 65978 425728 65984 425740
rect 50948 425700 65984 425728
rect 50948 425688 50954 425700
rect 65978 425688 65984 425700
rect 66036 425728 66042 425740
rect 66530 425728 66536 425740
rect 66036 425700 66536 425728
rect 66036 425688 66042 425700
rect 66530 425688 66536 425700
rect 66588 425688 66594 425740
rect 115842 425076 115848 425128
rect 115900 425116 115906 425128
rect 118786 425116 118792 425128
rect 115900 425088 118792 425116
rect 115900 425076 115906 425088
rect 118786 425076 118792 425088
rect 118844 425076 118850 425128
rect 115842 424328 115848 424380
rect 115900 424368 115906 424380
rect 144914 424368 144920 424380
rect 115900 424340 144920 424368
rect 115900 424328 115906 424340
rect 144914 424328 144920 424340
rect 144972 424328 144978 424380
rect 44082 423648 44088 423700
rect 44140 423688 44146 423700
rect 66714 423688 66720 423700
rect 44140 423660 66720 423688
rect 44140 423648 44146 423660
rect 66714 423648 66720 423660
rect 66772 423648 66778 423700
rect 115750 423648 115756 423700
rect 115808 423688 115814 423700
rect 126974 423688 126980 423700
rect 115808 423660 126980 423688
rect 115808 423648 115814 423660
rect 126974 423648 126980 423660
rect 127032 423648 127038 423700
rect 2774 423580 2780 423632
rect 2832 423620 2838 423632
rect 4798 423620 4804 423632
rect 2832 423592 4804 423620
rect 2832 423580 2838 423592
rect 4798 423580 4804 423592
rect 4856 423580 4862 423632
rect 115842 423580 115848 423632
rect 115900 423620 115906 423632
rect 122926 423620 122932 423632
rect 115900 423592 122932 423620
rect 115900 423580 115906 423592
rect 122926 423580 122932 423592
rect 122984 423620 122990 423632
rect 124122 423620 124128 423632
rect 122984 423592 124128 423620
rect 122984 423580 122990 423592
rect 124122 423580 124128 423592
rect 124180 423580 124186 423632
rect 60734 423444 60740 423496
rect 60792 423484 60798 423496
rect 61838 423484 61844 423496
rect 60792 423456 61844 423484
rect 60792 423444 60798 423456
rect 61838 423444 61844 423456
rect 61896 423484 61902 423496
rect 66714 423484 66720 423496
rect 61896 423456 66720 423484
rect 61896 423444 61902 423456
rect 66714 423444 66720 423456
rect 66772 423444 66778 423496
rect 49602 422900 49608 422952
rect 49660 422940 49666 422952
rect 60734 422940 60740 422952
rect 49660 422912 60740 422940
rect 49660 422900 49666 422912
rect 60734 422900 60740 422912
rect 60792 422900 60798 422952
rect 124122 422900 124128 422952
rect 124180 422940 124186 422952
rect 148318 422940 148324 422952
rect 124180 422912 148324 422940
rect 124180 422900 124186 422912
rect 148318 422900 148324 422912
rect 148376 422900 148382 422952
rect 50982 422220 50988 422272
rect 51040 422260 51046 422272
rect 66990 422260 66996 422272
rect 51040 422232 66996 422260
rect 51040 422220 51046 422232
rect 66990 422220 66996 422232
rect 67048 422220 67054 422272
rect 41230 421540 41236 421592
rect 41288 421580 41294 421592
rect 50982 421580 50988 421592
rect 41288 421552 50988 421580
rect 41288 421540 41294 421552
rect 50982 421540 50988 421552
rect 51040 421540 51046 421592
rect 114554 421540 114560 421592
rect 114612 421580 114618 421592
rect 146938 421580 146944 421592
rect 114612 421552 146944 421580
rect 114612 421540 114618 421552
rect 146938 421540 146944 421552
rect 146996 421540 147002 421592
rect 61838 419500 61844 419552
rect 61896 419540 61902 419552
rect 66898 419540 66904 419552
rect 61896 419512 66904 419540
rect 61896 419500 61902 419512
rect 66898 419500 66904 419512
rect 66956 419500 66962 419552
rect 115750 419500 115756 419552
rect 115808 419540 115814 419552
rect 129826 419540 129832 419552
rect 115808 419512 129832 419540
rect 115808 419500 115814 419512
rect 129826 419500 129832 419512
rect 129884 419500 129890 419552
rect 66898 418248 66904 418260
rect 45526 418220 66904 418248
rect 32950 418140 32956 418192
rect 33008 418180 33014 418192
rect 45526 418180 45554 418220
rect 66898 418208 66904 418220
rect 66956 418208 66962 418260
rect 33008 418152 45554 418180
rect 33008 418140 33014 418152
rect 64782 418140 64788 418192
rect 64840 418180 64846 418192
rect 66622 418180 66628 418192
rect 64840 418152 66628 418180
rect 64840 418140 64846 418152
rect 66622 418140 66628 418152
rect 66680 418140 66686 418192
rect 57790 417392 57796 417444
rect 57848 417432 57854 417444
rect 66622 417432 66628 417444
rect 57848 417404 66628 417432
rect 57848 417392 57854 417404
rect 66622 417392 66628 417404
rect 66680 417392 66686 417444
rect 64138 416848 64144 416900
rect 64196 416888 64202 416900
rect 66990 416888 66996 416900
rect 64196 416860 66996 416888
rect 64196 416848 64202 416860
rect 66990 416848 66996 416860
rect 67048 416848 67054 416900
rect 115842 416780 115848 416832
rect 115900 416820 115906 416832
rect 143534 416820 143540 416832
rect 115900 416792 143540 416820
rect 115900 416780 115906 416792
rect 143534 416780 143540 416792
rect 143592 416780 143598 416832
rect 116210 416712 116216 416764
rect 116268 416752 116274 416764
rect 118970 416752 118976 416764
rect 116268 416724 118976 416752
rect 116268 416712 116274 416724
rect 118970 416712 118976 416724
rect 119028 416712 119034 416764
rect 115842 415692 115848 415744
rect 115900 415732 115906 415744
rect 116210 415732 116216 415744
rect 115900 415704 116216 415732
rect 115900 415692 115906 415704
rect 116210 415692 116216 415704
rect 116268 415692 116274 415744
rect 53558 415420 53564 415472
rect 53616 415460 53622 415472
rect 59998 415460 60004 415472
rect 53616 415432 60004 415460
rect 53616 415420 53622 415432
rect 59998 415420 60004 415432
rect 60056 415420 60062 415472
rect 115842 414808 115848 414860
rect 115900 414848 115906 414860
rect 117314 414848 117320 414860
rect 115900 414820 117320 414848
rect 115900 414808 115906 414820
rect 117314 414808 117320 414820
rect 117372 414848 117378 414860
rect 121638 414848 121644 414860
rect 117372 414820 121644 414848
rect 117372 414808 117378 414820
rect 121638 414808 121644 414820
rect 121696 414808 121702 414860
rect 59998 414740 60004 414792
rect 60056 414780 60062 414792
rect 66898 414780 66904 414792
rect 60056 414752 66904 414780
rect 60056 414740 60062 414752
rect 66898 414740 66904 414752
rect 66956 414740 66962 414792
rect 56410 413992 56416 414044
rect 56468 414032 56474 414044
rect 66714 414032 66720 414044
rect 56468 414004 66720 414032
rect 56468 413992 56474 414004
rect 66714 413992 66720 414004
rect 66772 413992 66778 414044
rect 115106 413992 115112 414044
rect 115164 414032 115170 414044
rect 115290 414032 115296 414044
rect 115164 414004 115296 414032
rect 115164 413992 115170 414004
rect 115290 413992 115296 414004
rect 115348 414032 115354 414044
rect 147674 414032 147680 414044
rect 115348 414004 147680 414032
rect 115348 413992 115354 414004
rect 147674 413992 147680 414004
rect 147732 413992 147738 414044
rect 46842 413244 46848 413296
rect 46900 413284 46906 413296
rect 59262 413284 59268 413296
rect 46900 413256 59268 413284
rect 46900 413244 46906 413256
rect 59262 413244 59268 413256
rect 59320 413284 59326 413296
rect 66898 413284 66904 413296
rect 59320 413256 66904 413284
rect 59320 413244 59326 413256
rect 66898 413244 66904 413256
rect 66956 413244 66962 413296
rect 115842 412632 115848 412684
rect 115900 412672 115906 412684
rect 121546 412672 121552 412684
rect 115900 412644 121552 412672
rect 115900 412632 115906 412644
rect 121546 412632 121552 412644
rect 121604 412672 121610 412684
rect 122926 412672 122932 412684
rect 121604 412644 122932 412672
rect 121604 412632 121610 412644
rect 122926 412632 122932 412644
rect 122984 412632 122990 412684
rect 115198 411884 115204 411936
rect 115256 411924 115262 411936
rect 116118 411924 116124 411936
rect 115256 411896 116124 411924
rect 115256 411884 115262 411896
rect 116118 411884 116124 411896
rect 116176 411924 116182 411936
rect 142154 411924 142160 411936
rect 116176 411896 142160 411924
rect 116176 411884 116182 411896
rect 142154 411884 142160 411896
rect 142212 411884 142218 411936
rect 59262 411272 59268 411324
rect 59320 411312 59326 411324
rect 64598 411312 64604 411324
rect 59320 411284 64604 411312
rect 59320 411272 59326 411284
rect 64598 411272 64604 411284
rect 64656 411312 64662 411324
rect 66714 411312 66720 411324
rect 64656 411284 66720 411312
rect 64656 411272 64662 411284
rect 66714 411272 66720 411284
rect 66772 411272 66778 411324
rect 52270 411204 52276 411256
rect 52328 411244 52334 411256
rect 66898 411244 66904 411256
rect 52328 411216 66904 411244
rect 52328 411204 52334 411216
rect 66898 411204 66904 411216
rect 66956 411204 66962 411256
rect 115842 411204 115848 411256
rect 115900 411244 115906 411256
rect 123202 411244 123208 411256
rect 115900 411216 123208 411244
rect 115900 411204 115906 411216
rect 123202 411204 123208 411216
rect 123260 411244 123266 411256
rect 124122 411244 124128 411256
rect 123260 411216 124128 411244
rect 123260 411204 123266 411216
rect 124122 411204 124128 411216
rect 124180 411204 124186 411256
rect 124122 410524 124128 410576
rect 124180 410564 124186 410576
rect 136634 410564 136640 410576
rect 124180 410536 136640 410564
rect 124180 410524 124186 410536
rect 136634 410524 136640 410536
rect 136692 410524 136698 410576
rect 50982 409912 50988 409964
rect 51040 409952 51046 409964
rect 52270 409952 52276 409964
rect 51040 409924 52276 409952
rect 51040 409912 51046 409924
rect 52270 409912 52276 409924
rect 52328 409912 52334 409964
rect 2866 409844 2872 409896
rect 2924 409884 2930 409896
rect 51718 409884 51724 409896
rect 2924 409856 51724 409884
rect 2924 409844 2930 409856
rect 51718 409844 51724 409856
rect 51776 409844 51782 409896
rect 53834 409776 53840 409828
rect 53892 409816 53898 409828
rect 55030 409816 55036 409828
rect 53892 409788 55036 409816
rect 53892 409776 53898 409788
rect 55030 409776 55036 409788
rect 55088 409816 55094 409828
rect 66254 409816 66260 409828
rect 55088 409788 66260 409816
rect 55088 409776 55094 409788
rect 66254 409776 66260 409788
rect 66312 409776 66318 409828
rect 115842 409776 115848 409828
rect 115900 409816 115906 409828
rect 120258 409816 120264 409828
rect 115900 409788 120264 409816
rect 115900 409776 115906 409788
rect 120258 409776 120264 409788
rect 120316 409776 120322 409828
rect 39942 409096 39948 409148
rect 40000 409136 40006 409148
rect 53834 409136 53840 409148
rect 40000 409108 53840 409136
rect 40000 409096 40006 409108
rect 53834 409096 53840 409108
rect 53892 409096 53898 409148
rect 120258 409096 120264 409148
rect 120316 409136 120322 409148
rect 139394 409136 139400 409148
rect 120316 409108 139400 409136
rect 120316 409096 120322 409108
rect 139394 409096 139400 409108
rect 139452 409096 139458 409148
rect 39850 408416 39856 408468
rect 39908 408456 39914 408468
rect 66898 408456 66904 408468
rect 39908 408428 66904 408456
rect 39908 408416 39914 408428
rect 66898 408416 66904 408428
rect 66956 408416 66962 408468
rect 35802 407736 35808 407788
rect 35860 407776 35866 407788
rect 39850 407776 39856 407788
rect 35860 407748 39856 407776
rect 35860 407736 35866 407748
rect 39850 407736 39856 407748
rect 39908 407736 39914 407788
rect 115014 407464 115020 407516
rect 115072 407504 115078 407516
rect 121546 407504 121552 407516
rect 115072 407476 121552 407504
rect 115072 407464 115078 407476
rect 121546 407464 121552 407476
rect 121604 407464 121610 407516
rect 56502 407056 56508 407108
rect 56560 407096 56566 407108
rect 57790 407096 57796 407108
rect 56560 407068 57796 407096
rect 56560 407056 56566 407068
rect 57790 407056 57796 407068
rect 57848 407056 57854 407108
rect 112714 407056 112720 407108
rect 112772 407096 112778 407108
rect 117590 407096 117596 407108
rect 112772 407068 117596 407096
rect 112772 407056 112778 407068
rect 117590 407056 117596 407068
rect 117648 407056 117654 407108
rect 57790 405696 57796 405748
rect 57848 405736 57854 405748
rect 66438 405736 66444 405748
rect 57848 405708 66444 405736
rect 57848 405696 57854 405708
rect 66438 405696 66444 405708
rect 66496 405696 66502 405748
rect 115842 405628 115848 405680
rect 115900 405668 115906 405680
rect 140774 405668 140780 405680
rect 115900 405640 140780 405668
rect 115900 405628 115906 405640
rect 140774 405628 140780 405640
rect 140832 405668 140838 405680
rect 141418 405668 141424 405680
rect 140832 405640 141424 405668
rect 140832 405628 140838 405640
rect 141418 405628 141424 405640
rect 141476 405628 141482 405680
rect 117314 405560 117320 405612
rect 117372 405600 117378 405612
rect 117498 405600 117504 405612
rect 117372 405572 117504 405600
rect 117372 405560 117378 405572
rect 117498 405560 117504 405572
rect 117556 405560 117562 405612
rect 115842 404540 115848 404592
rect 115900 404580 115906 404592
rect 117314 404580 117320 404592
rect 115900 404552 117320 404580
rect 115900 404540 115906 404552
rect 117314 404540 117320 404552
rect 117372 404540 117378 404592
rect 63218 404336 63224 404388
rect 63276 404376 63282 404388
rect 66898 404376 66904 404388
rect 63276 404348 66904 404376
rect 63276 404336 63282 404348
rect 66898 404336 66904 404348
rect 66956 404336 66962 404388
rect 141418 404336 141424 404388
rect 141476 404376 141482 404388
rect 143626 404376 143632 404388
rect 141476 404348 143632 404376
rect 141476 404336 141482 404348
rect 143626 404336 143632 404348
rect 143684 404336 143690 404388
rect 115842 402976 115848 403028
rect 115900 403016 115906 403028
rect 126330 403016 126336 403028
rect 115900 402988 126336 403016
rect 115900 402976 115906 402988
rect 126330 402976 126336 402988
rect 126388 402976 126394 403028
rect 115842 401956 115848 402008
rect 115900 401996 115906 402008
rect 118970 401996 118976 402008
rect 115900 401968 118976 401996
rect 115900 401956 115906 401968
rect 118970 401956 118976 401968
rect 119028 401996 119034 402008
rect 120166 401996 120172 402008
rect 119028 401968 120172 401996
rect 119028 401956 119034 401968
rect 120166 401956 120172 401968
rect 120224 401956 120230 402008
rect 115842 401548 115848 401600
rect 115900 401588 115906 401600
rect 128446 401588 128452 401600
rect 115900 401560 128452 401588
rect 115900 401548 115906 401560
rect 128446 401548 128452 401560
rect 128504 401548 128510 401600
rect 128446 400868 128452 400920
rect 128504 400908 128510 400920
rect 146294 400908 146300 400920
rect 128504 400880 146300 400908
rect 128504 400868 128510 400880
rect 146294 400868 146300 400880
rect 146352 400868 146358 400920
rect 58894 400256 58900 400308
rect 58952 400296 58958 400308
rect 66806 400296 66812 400308
rect 58952 400268 66812 400296
rect 58952 400256 58958 400268
rect 66806 400256 66812 400268
rect 66864 400256 66870 400308
rect 57606 400188 57612 400240
rect 57664 400228 57670 400240
rect 66898 400228 66904 400240
rect 57664 400200 66904 400228
rect 57664 400188 57670 400200
rect 66898 400188 66904 400200
rect 66956 400188 66962 400240
rect 115382 399168 115388 399220
rect 115440 399208 115446 399220
rect 117498 399208 117504 399220
rect 115440 399180 117504 399208
rect 115440 399168 115446 399180
rect 117498 399168 117504 399180
rect 117556 399168 117562 399220
rect 55030 398828 55036 398880
rect 55088 398868 55094 398880
rect 66530 398868 66536 398880
rect 55088 398840 66536 398868
rect 55088 398828 55094 398840
rect 66530 398828 66536 398840
rect 66588 398828 66594 398880
rect 3510 397536 3516 397588
rect 3568 397576 3574 397588
rect 21358 397576 21364 397588
rect 3568 397548 21364 397576
rect 3568 397536 3574 397548
rect 21358 397536 21364 397548
rect 21416 397536 21422 397588
rect 67358 397576 67364 397588
rect 64846 397548 67364 397576
rect 11698 397468 11704 397520
rect 11756 397508 11762 397520
rect 64846 397508 64874 397548
rect 67358 397536 67364 397548
rect 67416 397576 67422 397588
rect 67726 397576 67732 397588
rect 67416 397548 67732 397576
rect 67416 397536 67422 397548
rect 67726 397536 67732 397548
rect 67784 397536 67790 397588
rect 11756 397480 64874 397508
rect 11756 397468 11762 397480
rect 115566 397468 115572 397520
rect 115624 397508 115630 397520
rect 124214 397508 124220 397520
rect 115624 397480 124220 397508
rect 115624 397468 115630 397480
rect 124214 397468 124220 397480
rect 124272 397468 124278 397520
rect 66714 397400 66720 397452
rect 66772 397440 66778 397452
rect 67726 397440 67732 397452
rect 66772 397412 67732 397440
rect 66772 397400 66778 397412
rect 67726 397400 67732 397412
rect 67784 397400 67790 397452
rect 128446 397400 128452 397452
rect 128504 397440 128510 397452
rect 132586 397440 132592 397452
rect 128504 397412 132592 397440
rect 128504 397400 128510 397412
rect 132586 397400 132592 397412
rect 132644 397400 132650 397452
rect 42702 396788 42708 396840
rect 42760 396828 42766 396840
rect 59170 396828 59176 396840
rect 42760 396800 59176 396828
rect 42760 396788 42766 396800
rect 59170 396788 59176 396800
rect 59228 396828 59234 396840
rect 66622 396828 66628 396840
rect 59228 396800 66628 396828
rect 59228 396788 59234 396800
rect 66622 396788 66628 396800
rect 66680 396788 66686 396840
rect 35710 396720 35716 396772
rect 35768 396760 35774 396772
rect 35768 396732 45554 396760
rect 35768 396720 35774 396732
rect 45526 396692 45554 396732
rect 117498 396720 117504 396772
rect 117556 396760 117562 396772
rect 149054 396760 149060 396772
rect 117556 396732 149060 396760
rect 117556 396720 117562 396732
rect 149054 396720 149060 396732
rect 149112 396720 149118 396772
rect 67082 396692 67088 396704
rect 45526 396664 67088 396692
rect 67082 396652 67088 396664
rect 67140 396652 67146 396704
rect 115842 396040 115848 396092
rect 115900 396080 115906 396092
rect 128446 396080 128452 396092
rect 115900 396052 128452 396080
rect 115900 396040 115906 396052
rect 128446 396040 128452 396052
rect 128504 396040 128510 396092
rect 49510 395972 49516 396024
rect 49568 396012 49574 396024
rect 66806 396012 66812 396024
rect 49568 395984 66812 396012
rect 49568 395972 49574 395984
rect 66806 395972 66812 395984
rect 66864 395972 66870 396024
rect 48222 395224 48228 395276
rect 48280 395264 48286 395276
rect 49510 395264 49516 395276
rect 48280 395236 49516 395264
rect 48280 395224 48286 395236
rect 49510 395224 49516 395236
rect 49568 395224 49574 395276
rect 115842 394680 115848 394732
rect 115900 394720 115906 394732
rect 190454 394720 190460 394732
rect 115900 394692 190460 394720
rect 115900 394680 115906 394692
rect 190454 394680 190460 394692
rect 190512 394680 190518 394732
rect 43990 393932 43996 393984
rect 44048 393972 44054 393984
rect 49510 393972 49516 393984
rect 44048 393944 49516 393972
rect 44048 393932 44054 393944
rect 49510 393932 49516 393944
rect 49568 393932 49574 393984
rect 49510 393320 49516 393372
rect 49568 393360 49574 393372
rect 66806 393360 66812 393372
rect 49568 393332 66812 393360
rect 49568 393320 49574 393332
rect 66806 393320 66812 393332
rect 66864 393320 66870 393372
rect 115842 393252 115848 393304
rect 115900 393292 115906 393304
rect 128354 393292 128360 393304
rect 115900 393264 128360 393292
rect 115900 393252 115906 393264
rect 128354 393252 128360 393264
rect 128412 393252 128418 393304
rect 53650 392572 53656 392624
rect 53708 392612 53714 392624
rect 66346 392612 66352 392624
rect 53708 392584 66352 392612
rect 53708 392572 53714 392584
rect 66346 392572 66352 392584
rect 66404 392572 66410 392624
rect 56502 391960 56508 392012
rect 56560 392000 56566 392012
rect 66806 392000 66812 392012
rect 56560 391972 66812 392000
rect 56560 391960 56566 391972
rect 66806 391960 66812 391972
rect 66864 391960 66870 392012
rect 128354 391960 128360 392012
rect 128412 392000 128418 392012
rect 134058 392000 134064 392012
rect 128412 391972 134064 392000
rect 128412 391960 128418 391972
rect 134058 391960 134064 391972
rect 134116 391960 134122 392012
rect 41322 391280 41328 391332
rect 41380 391320 41386 391332
rect 41380 391292 87736 391320
rect 41380 391280 41386 391292
rect 3418 391212 3424 391264
rect 3476 391252 3482 391264
rect 3476 391224 84194 391252
rect 3476 391212 3482 391224
rect 84166 390912 84194 391224
rect 87708 390992 87736 391292
rect 118878 391212 118884 391264
rect 118936 391252 118942 391264
rect 138014 391252 138020 391264
rect 118936 391224 138020 391252
rect 118936 391212 118942 391224
rect 138014 391212 138020 391224
rect 138072 391212 138078 391264
rect 115014 391144 115020 391196
rect 115072 391184 115078 391196
rect 120166 391184 120172 391196
rect 115072 391156 120172 391184
rect 115072 391144 115078 391156
rect 120166 391144 120172 391156
rect 120224 391144 120230 391196
rect 87690 390940 87696 390992
rect 87748 390940 87754 390992
rect 108666 390940 108672 390992
rect 108724 390980 108730 390992
rect 118878 390980 118884 390992
rect 108724 390952 118884 390980
rect 108724 390940 108730 390952
rect 118878 390940 118884 390952
rect 118936 390940 118942 390992
rect 93670 390912 93676 390924
rect 84166 390884 93676 390912
rect 93670 390872 93676 390884
rect 93728 390872 93734 390924
rect 67634 390124 67640 390176
rect 67692 390164 67698 390176
rect 68784 390164 68790 390176
rect 67692 390136 68790 390164
rect 67692 390124 67698 390136
rect 68784 390124 68790 390136
rect 68842 390124 68848 390176
rect 102042 389784 102048 389836
rect 102100 389824 102106 389836
rect 113266 389824 113272 389836
rect 102100 389796 113272 389824
rect 102100 389784 102106 389796
rect 113266 389784 113272 389796
rect 113324 389784 113330 389836
rect 118694 389784 118700 389836
rect 118752 389824 118758 389836
rect 128354 389824 128360 389836
rect 118752 389796 128360 389824
rect 118752 389784 118758 389796
rect 128354 389784 128360 389796
rect 128412 389784 128418 389836
rect 94590 389484 94596 389496
rect 86926 389456 94596 389484
rect 86926 389416 86954 389456
rect 94590 389444 94596 389456
rect 94648 389444 94654 389496
rect 100754 389416 100760 389428
rect 84166 389388 86954 389416
rect 91756 389388 100760 389416
rect 62022 389240 62028 389292
rect 62080 389280 62086 389292
rect 84166 389280 84194 389388
rect 62080 389252 84194 389280
rect 62080 389240 62086 389252
rect 36538 389172 36544 389224
rect 36596 389212 36602 389224
rect 91756 389212 91784 389388
rect 100754 389376 100760 389388
rect 100812 389376 100818 389428
rect 94590 389308 94596 389360
rect 94648 389348 94654 389360
rect 98270 389348 98276 389360
rect 94648 389320 98276 389348
rect 94648 389308 94654 389320
rect 36596 389184 91784 389212
rect 36596 389172 36602 389184
rect 97368 389174 97396 389320
rect 98270 389308 98276 389320
rect 98328 389308 98334 389360
rect 97276 389156 97396 389174
rect 101674 389172 101680 389224
rect 101732 389212 101738 389224
rect 118694 389212 118700 389224
rect 101732 389184 118700 389212
rect 101732 389172 101738 389184
rect 118694 389172 118700 389184
rect 118752 389172 118758 389224
rect 48038 389104 48044 389156
rect 48096 389144 48102 389156
rect 82998 389144 83004 389156
rect 48096 389116 83004 389144
rect 48096 389104 48102 389116
rect 82998 389104 83004 389116
rect 83056 389104 83062 389156
rect 97258 389104 97264 389156
rect 97316 389146 97396 389156
rect 97316 389104 97322 389146
rect 110138 389036 110144 389088
rect 110196 389076 110202 389088
rect 124766 389076 124772 389088
rect 110196 389048 124772 389076
rect 110196 389036 110202 389048
rect 124766 389036 124772 389048
rect 124824 389036 124830 389088
rect 46750 388696 46756 388748
rect 46808 388736 46814 388748
rect 48038 388736 48044 388748
rect 46808 388708 48044 388736
rect 46808 388696 46814 388708
rect 48038 388696 48044 388708
rect 48096 388696 48102 388748
rect 102226 388492 102232 388544
rect 102284 388532 102290 388544
rect 106366 388532 106372 388544
rect 102284 388504 106372 388532
rect 102284 388492 102290 388504
rect 106366 388492 106372 388504
rect 106424 388492 106430 388544
rect 84102 388424 84108 388476
rect 84160 388464 84166 388476
rect 104158 388464 104164 388476
rect 84160 388436 104164 388464
rect 84160 388424 84166 388436
rect 104158 388424 104164 388436
rect 104216 388424 104222 388476
rect 105538 388424 105544 388476
rect 105596 388464 105602 388476
rect 114738 388464 114744 388476
rect 105596 388436 114744 388464
rect 105596 388424 105602 388436
rect 114738 388424 114744 388436
rect 114796 388424 114802 388476
rect 71682 387812 71688 387864
rect 71740 387852 71746 387864
rect 73246 387852 73252 387864
rect 71740 387824 73252 387852
rect 71740 387812 71746 387824
rect 73246 387812 73252 387824
rect 73304 387812 73310 387864
rect 79962 387812 79968 387864
rect 80020 387852 80026 387864
rect 80698 387852 80704 387864
rect 80020 387824 80704 387852
rect 80020 387812 80026 387824
rect 80698 387812 80704 387824
rect 80756 387812 80762 387864
rect 84930 387812 84936 387864
rect 84988 387852 84994 387864
rect 86218 387852 86224 387864
rect 84988 387824 86224 387852
rect 84988 387812 84994 387824
rect 86218 387812 86224 387824
rect 86276 387812 86282 387864
rect 90358 387812 90364 387864
rect 90416 387852 90422 387864
rect 91370 387852 91376 387864
rect 90416 387824 91376 387852
rect 90416 387812 90422 387824
rect 91370 387812 91376 387824
rect 91428 387812 91434 387864
rect 93118 387812 93124 387864
rect 93176 387852 93182 387864
rect 96982 387852 96988 387864
rect 93176 387824 96988 387852
rect 93176 387812 93182 387824
rect 96982 387812 96988 387824
rect 97040 387812 97046 387864
rect 100570 387812 100576 387864
rect 100628 387852 100634 387864
rect 102502 387852 102508 387864
rect 100628 387824 102508 387852
rect 100628 387812 100634 387824
rect 102502 387812 102508 387824
rect 102560 387812 102566 387864
rect 57882 387744 57888 387796
rect 57940 387784 57946 387796
rect 96614 387784 96620 387796
rect 57940 387756 96620 387784
rect 57940 387744 57946 387756
rect 96614 387744 96620 387756
rect 96672 387744 96678 387796
rect 120718 387744 120724 387796
rect 120776 387784 120782 387796
rect 121454 387784 121460 387796
rect 120776 387756 121460 387784
rect 120776 387744 120782 387756
rect 121454 387744 121460 387756
rect 121512 387744 121518 387796
rect 101858 387132 101864 387184
rect 101916 387172 101922 387184
rect 107654 387172 107660 387184
rect 101916 387144 107660 387172
rect 101916 387132 101922 387144
rect 107654 387132 107660 387144
rect 107712 387132 107718 387184
rect 52270 387064 52276 387116
rect 52328 387104 52334 387116
rect 73982 387104 73988 387116
rect 52328 387076 73988 387104
rect 52328 387064 52334 387076
rect 73982 387064 73988 387076
rect 74040 387064 74046 387116
rect 86862 387064 86868 387116
rect 86920 387104 86926 387116
rect 120718 387104 120724 387116
rect 86920 387076 120724 387104
rect 86920 387064 86926 387076
rect 120718 387064 120724 387076
rect 120776 387064 120782 387116
rect 84194 386996 84200 387048
rect 84252 387036 84258 387048
rect 85022 387036 85028 387048
rect 84252 387008 85028 387036
rect 84252 386996 84258 387008
rect 85022 386996 85028 387008
rect 85080 386996 85086 387048
rect 111794 386996 111800 387048
rect 111852 387036 111858 387048
rect 112254 387036 112260 387048
rect 111852 387008 112260 387036
rect 111852 386996 111858 387008
rect 112254 386996 112260 387008
rect 112312 386996 112318 387048
rect 96614 386384 96620 386436
rect 96672 386424 96678 386436
rect 97350 386424 97356 386436
rect 96672 386396 97356 386424
rect 96672 386384 96678 386396
rect 97350 386384 97356 386396
rect 97408 386384 97414 386436
rect 65886 386316 65892 386368
rect 65944 386356 65950 386368
rect 72418 386356 72424 386368
rect 65944 386328 72424 386356
rect 65944 386316 65950 386328
rect 72418 386316 72424 386328
rect 72476 386316 72482 386368
rect 75178 386316 75184 386368
rect 75236 386356 75242 386368
rect 82262 386356 82268 386368
rect 75236 386328 82268 386356
rect 75236 386316 75242 386328
rect 82262 386316 82268 386328
rect 82320 386316 82326 386368
rect 115934 386356 115940 386368
rect 84166 386328 115940 386356
rect 80790 386248 80796 386300
rect 80848 386288 80854 386300
rect 81250 386288 81256 386300
rect 80848 386260 81256 386288
rect 80848 386248 80854 386260
rect 81250 386248 81256 386260
rect 81308 386288 81314 386300
rect 84166 386288 84194 386328
rect 115934 386316 115940 386328
rect 115992 386316 115998 386368
rect 81308 386260 84194 386288
rect 81308 386248 81314 386260
rect 100386 386248 100392 386300
rect 100444 386288 100450 386300
rect 129734 386288 129740 386300
rect 100444 386260 129740 386288
rect 100444 386248 100450 386260
rect 129734 386248 129740 386260
rect 129792 386288 129798 386300
rect 130286 386288 130292 386300
rect 129792 386260 130292 386288
rect 129792 386248 129798 386260
rect 130286 386248 130292 386260
rect 130344 386248 130350 386300
rect 54846 385636 54852 385688
rect 54904 385676 54910 385688
rect 66806 385676 66812 385688
rect 54904 385648 66812 385676
rect 54904 385636 54910 385648
rect 66806 385636 66812 385648
rect 66864 385636 66870 385688
rect 130286 385024 130292 385076
rect 130344 385064 130350 385076
rect 134150 385064 134156 385076
rect 130344 385036 134156 385064
rect 130344 385024 130350 385036
rect 134150 385024 134156 385036
rect 134208 385024 134214 385076
rect 55122 384956 55128 385008
rect 55180 384996 55186 385008
rect 92474 384996 92480 385008
rect 55180 384968 92480 384996
rect 55180 384956 55186 384968
rect 92474 384956 92480 384968
rect 92532 384956 92538 385008
rect 133138 384956 133144 385008
rect 133196 384996 133202 385008
rect 133874 384996 133880 385008
rect 133196 384968 133880 384996
rect 133196 384956 133202 384968
rect 133874 384956 133880 384968
rect 133932 384956 133938 385008
rect 91186 384344 91192 384396
rect 91244 384384 91250 384396
rect 109126 384384 109132 384396
rect 91244 384356 109132 384384
rect 91244 384344 91250 384356
rect 109126 384344 109132 384356
rect 109184 384344 109190 384396
rect 105170 384276 105176 384328
rect 105228 384316 105234 384328
rect 133138 384316 133144 384328
rect 105228 384288 133144 384316
rect 105228 384276 105234 384288
rect 133138 384276 133144 384288
rect 133196 384276 133202 384328
rect 88426 383596 88432 383648
rect 88484 383636 88490 383648
rect 120074 383636 120080 383648
rect 88484 383608 120080 383636
rect 88484 383596 88490 383608
rect 120074 383596 120080 383608
rect 120132 383596 120138 383648
rect 101766 382916 101772 382968
rect 101824 382956 101830 382968
rect 112714 382956 112720 382968
rect 101824 382928 112720 382956
rect 101824 382916 101830 382928
rect 112714 382916 112720 382928
rect 112772 382916 112778 382968
rect 120074 382236 120080 382288
rect 120132 382276 120138 382288
rect 122834 382276 122840 382288
rect 120132 382248 122840 382276
rect 120132 382236 120138 382248
rect 122834 382236 122840 382248
rect 122892 382236 122898 382288
rect 45462 381488 45468 381540
rect 45520 381528 45526 381540
rect 71774 381528 71780 381540
rect 45520 381500 71780 381528
rect 45520 381488 45526 381500
rect 71774 381488 71780 381500
rect 71832 381488 71838 381540
rect 84194 381488 84200 381540
rect 84252 381528 84258 381540
rect 117314 381528 117320 381540
rect 84252 381500 117320 381528
rect 84252 381488 84258 381500
rect 117314 381488 117320 381500
rect 117372 381488 117378 381540
rect 21358 380808 21364 380860
rect 21416 380848 21422 380860
rect 116210 380848 116216 380860
rect 21416 380820 116216 380848
rect 21416 380808 21422 380820
rect 116210 380808 116216 380820
rect 116268 380808 116274 380860
rect 94498 380128 94504 380180
rect 94556 380168 94562 380180
rect 128538 380168 128544 380180
rect 94556 380140 128544 380168
rect 94556 380128 94562 380140
rect 128538 380128 128544 380140
rect 128596 380128 128602 380180
rect 115934 380060 115940 380112
rect 115992 380100 115998 380112
rect 116210 380100 116216 380112
rect 115992 380072 116216 380100
rect 115992 380060 115998 380072
rect 116210 380060 116216 380072
rect 116268 380060 116274 380112
rect 79962 379516 79968 379568
rect 80020 379556 80026 379568
rect 81434 379556 81440 379568
rect 80020 379528 81440 379556
rect 80020 379516 80026 379528
rect 81434 379516 81440 379528
rect 81492 379516 81498 379568
rect 88242 379448 88248 379500
rect 88300 379488 88306 379500
rect 91370 379488 91376 379500
rect 88300 379460 91376 379488
rect 88300 379448 88306 379460
rect 91370 379448 91376 379460
rect 91428 379448 91434 379500
rect 43990 378768 43996 378820
rect 44048 378808 44054 378820
rect 80054 378808 80060 378820
rect 44048 378780 80060 378808
rect 44048 378768 44054 378780
rect 80054 378768 80060 378780
rect 80112 378768 80118 378820
rect 100478 378768 100484 378820
rect 100536 378808 100542 378820
rect 129734 378808 129740 378820
rect 100536 378780 129740 378808
rect 100536 378768 100542 378780
rect 129734 378768 129740 378780
rect 129792 378768 129798 378820
rect 97810 378224 97816 378276
rect 97868 378264 97874 378276
rect 102318 378264 102324 378276
rect 97868 378236 102324 378264
rect 97868 378224 97874 378236
rect 102318 378224 102324 378236
rect 102376 378224 102382 378276
rect 92290 378088 92296 378140
rect 92348 378128 92354 378140
rect 93118 378128 93124 378140
rect 92348 378100 93124 378128
rect 92348 378088 92354 378100
rect 93118 378088 93124 378100
rect 93176 378088 93182 378140
rect 87690 377476 87696 377528
rect 87748 377516 87754 377528
rect 118694 377516 118700 377528
rect 87748 377488 118700 377516
rect 87748 377476 87754 377488
rect 118694 377476 118700 377488
rect 118752 377476 118758 377528
rect 33042 377408 33048 377460
rect 33100 377448 33106 377460
rect 92290 377448 92296 377460
rect 33100 377420 92296 377448
rect 33100 377408 33106 377420
rect 92290 377408 92296 377420
rect 92348 377408 92354 377460
rect 41322 374620 41328 374672
rect 41380 374660 41386 374672
rect 76006 374660 76012 374672
rect 41380 374632 76012 374660
rect 41380 374620 41386 374632
rect 76006 374620 76012 374632
rect 76064 374620 76070 374672
rect 86770 374620 86776 374672
rect 86828 374660 86834 374672
rect 95326 374660 95332 374672
rect 86828 374632 95332 374660
rect 86828 374620 86834 374632
rect 95326 374620 95332 374632
rect 95384 374620 95390 374672
rect 101950 373260 101956 373312
rect 102008 373300 102014 373312
rect 113174 373300 113180 373312
rect 102008 373272 113180 373300
rect 102008 373260 102014 373272
rect 113174 373260 113180 373272
rect 113232 373260 113238 373312
rect 3418 371220 3424 371272
rect 3476 371260 3482 371272
rect 3476 371232 106228 371260
rect 3476 371220 3482 371232
rect 106200 371204 106228 371232
rect 106182 371192 106188 371204
rect 106095 371164 106188 371192
rect 106182 371152 106188 371164
rect 106240 371192 106246 371204
rect 118970 371192 118976 371204
rect 106240 371164 118976 371192
rect 106240 371152 106246 371164
rect 118970 371152 118976 371164
rect 119028 371152 119034 371204
rect 50798 369112 50804 369164
rect 50856 369152 50862 369164
rect 75914 369152 75920 369164
rect 50856 369124 75920 369152
rect 50856 369112 50862 369124
rect 75914 369112 75920 369124
rect 75972 369112 75978 369164
rect 80698 369112 80704 369164
rect 80756 369152 80762 369164
rect 102134 369152 102140 369164
rect 80756 369124 102140 369152
rect 80756 369112 80762 369124
rect 102134 369112 102140 369124
rect 102192 369112 102198 369164
rect 85574 367752 85580 367804
rect 85632 367792 85638 367804
rect 106918 367792 106924 367804
rect 85632 367764 106924 367792
rect 85632 367752 85638 367764
rect 106918 367752 106924 367764
rect 106976 367752 106982 367804
rect 74534 366324 74540 366376
rect 74592 366364 74598 366376
rect 108298 366364 108304 366376
rect 74592 366336 108304 366364
rect 74592 366324 74598 366336
rect 108298 366324 108304 366336
rect 108356 366324 108362 366376
rect 269758 364352 269764 364404
rect 269816 364392 269822 364404
rect 580166 364392 580172 364404
rect 269816 364364 580172 364392
rect 269816 364352 269822 364364
rect 580166 364352 580172 364364
rect 580224 364352 580230 364404
rect 86218 363604 86224 363656
rect 86276 363644 86282 363656
rect 112438 363644 112444 363656
rect 86276 363616 112444 363644
rect 86276 363604 86282 363616
rect 112438 363604 112444 363616
rect 112496 363604 112502 363656
rect 77294 360816 77300 360868
rect 77352 360856 77358 360868
rect 110598 360856 110604 360868
rect 77352 360828 110604 360856
rect 77352 360816 77358 360828
rect 110598 360816 110604 360828
rect 110656 360816 110662 360868
rect 3326 358708 3332 358760
rect 3384 358748 3390 358760
rect 11698 358748 11704 358760
rect 3384 358720 11704 358748
rect 3384 358708 3390 358720
rect 11698 358708 11704 358720
rect 11756 358708 11762 358760
rect 3418 355308 3424 355360
rect 3476 355348 3482 355360
rect 33778 355348 33784 355360
rect 3476 355320 33784 355348
rect 3476 355308 3482 355320
rect 33778 355308 33784 355320
rect 33836 355308 33842 355360
rect 574738 351908 574744 351960
rect 574796 351948 574802 351960
rect 580166 351948 580172 351960
rect 574796 351920 580172 351948
rect 574796 351908 574802 351920
rect 580166 351908 580172 351920
rect 580224 351908 580230 351960
rect 3326 345040 3332 345092
rect 3384 345080 3390 345092
rect 18598 345080 18604 345092
rect 3384 345052 18604 345080
rect 3384 345040 3390 345052
rect 18598 345040 18604 345052
rect 18656 345040 18662 345092
rect 123478 343612 123484 343664
rect 123536 343652 123542 343664
rect 124122 343652 124128 343664
rect 123536 343624 124128 343652
rect 123536 343612 123542 343624
rect 124122 343612 124128 343624
rect 124180 343652 124186 343664
rect 260834 343652 260840 343664
rect 124180 343624 260840 343652
rect 124180 343612 124186 343624
rect 260834 343612 260840 343624
rect 260892 343612 260898 343664
rect 97718 342252 97724 342304
rect 97776 342292 97782 342304
rect 267826 342292 267832 342304
rect 97776 342264 267832 342292
rect 97776 342252 97782 342264
rect 267826 342252 267832 342264
rect 267884 342252 267890 342304
rect 124858 340892 124864 340944
rect 124916 340932 124922 340944
rect 125502 340932 125508 340944
rect 124916 340904 125508 340932
rect 124916 340892 124922 340904
rect 125502 340892 125508 340904
rect 125560 340932 125566 340944
rect 263594 340932 263600 340944
rect 125560 340904 263600 340932
rect 125560 340892 125566 340904
rect 263594 340892 263600 340904
rect 263652 340892 263658 340944
rect 83550 339464 83556 339516
rect 83608 339504 83614 339516
rect 259822 339504 259828 339516
rect 83608 339476 259828 339504
rect 83608 339464 83614 339476
rect 259822 339464 259828 339476
rect 259880 339464 259886 339516
rect 23382 338104 23388 338156
rect 23440 338144 23446 338156
rect 222194 338144 222200 338156
rect 23440 338116 222200 338144
rect 23440 338104 23446 338116
rect 222194 338104 222200 338116
rect 222252 338104 222258 338156
rect 153838 336812 153844 336864
rect 153896 336852 153902 336864
rect 233878 336852 233884 336864
rect 153896 336824 233884 336852
rect 153896 336812 153902 336824
rect 233878 336812 233884 336824
rect 233936 336812 233942 336864
rect 93118 336744 93124 336796
rect 93176 336784 93182 336796
rect 93670 336784 93676 336796
rect 93176 336756 93676 336784
rect 93176 336744 93182 336756
rect 93670 336744 93676 336756
rect 93728 336784 93734 336796
rect 255958 336784 255964 336796
rect 93728 336756 255964 336784
rect 93728 336744 93734 336756
rect 255958 336744 255964 336756
rect 256016 336744 256022 336796
rect 87598 335792 87604 335844
rect 87656 335832 87662 335844
rect 88242 335832 88248 335844
rect 87656 335804 88248 335832
rect 87656 335792 87662 335804
rect 88242 335792 88248 335804
rect 88300 335792 88306 335844
rect 88242 335316 88248 335368
rect 88300 335356 88306 335368
rect 256694 335356 256700 335368
rect 88300 335328 256700 335356
rect 88300 335316 88306 335328
rect 256694 335316 256700 335328
rect 256752 335316 256758 335368
rect 100018 333956 100024 334008
rect 100076 333996 100082 334008
rect 100570 333996 100576 334008
rect 100076 333968 100576 333996
rect 100076 333956 100082 333968
rect 100570 333956 100576 333968
rect 100628 333996 100634 334008
rect 246298 333996 246304 334008
rect 100628 333968 246304 333996
rect 100628 333956 100634 333968
rect 246298 333956 246304 333968
rect 246356 333956 246362 334008
rect 148410 332664 148416 332716
rect 148468 332704 148474 332716
rect 266446 332704 266452 332716
rect 148468 332676 266452 332704
rect 148468 332664 148474 332676
rect 266446 332664 266452 332676
rect 266504 332664 266510 332716
rect 99282 332596 99288 332648
rect 99340 332636 99346 332648
rect 244918 332636 244924 332648
rect 99340 332608 244924 332636
rect 99340 332596 99346 332608
rect 244918 332596 244924 332608
rect 244976 332596 244982 332648
rect 115198 331304 115204 331356
rect 115256 331344 115262 331356
rect 115382 331344 115388 331356
rect 115256 331316 115388 331344
rect 115256 331304 115262 331316
rect 115382 331304 115388 331316
rect 115440 331344 115446 331356
rect 244182 331344 244188 331356
rect 115440 331316 244188 331344
rect 115440 331304 115446 331316
rect 244182 331304 244188 331316
rect 244240 331304 244246 331356
rect 57606 331236 57612 331288
rect 57664 331276 57670 331288
rect 57882 331276 57888 331288
rect 57664 331248 57888 331276
rect 57664 331236 57670 331248
rect 57882 331236 57888 331248
rect 57940 331276 57946 331288
rect 266354 331276 266360 331288
rect 57940 331248 266360 331276
rect 57940 331236 57946 331248
rect 266354 331236 266360 331248
rect 266412 331236 266418 331288
rect 93670 331168 93676 331220
rect 93728 331208 93734 331220
rect 94038 331208 94044 331220
rect 93728 331180 94044 331208
rect 93728 331168 93734 331180
rect 94038 331168 94044 331180
rect 94096 331168 94102 331220
rect 166350 329808 166356 329860
rect 166408 329848 166414 329860
rect 227806 329848 227812 329860
rect 166408 329820 227812 329848
rect 166408 329808 166414 329820
rect 227806 329808 227812 329820
rect 227864 329808 227870 329860
rect 104802 328720 104808 328772
rect 104860 328760 104866 328772
rect 110506 328760 110512 328772
rect 104860 328732 110512 328760
rect 104860 328720 104866 328732
rect 110506 328720 110512 328732
rect 110564 328720 110570 328772
rect 192478 328516 192484 328568
rect 192536 328556 192542 328568
rect 250438 328556 250444 328568
rect 192536 328528 250444 328556
rect 192536 328516 192542 328528
rect 250438 328516 250444 328528
rect 250496 328516 250502 328568
rect 151078 328448 151084 328500
rect 151136 328488 151142 328500
rect 212534 328488 212540 328500
rect 151136 328460 212540 328488
rect 151136 328448 151142 328460
rect 212534 328448 212540 328460
rect 212592 328448 212598 328500
rect 81434 327700 81440 327752
rect 81492 327740 81498 327752
rect 91278 327740 91284 327752
rect 81492 327712 91284 327740
rect 81492 327700 81498 327712
rect 91278 327700 91284 327712
rect 91336 327700 91342 327752
rect 105722 327700 105728 327752
rect 105780 327740 105786 327752
rect 129826 327740 129832 327752
rect 105780 327712 129832 327740
rect 105780 327700 105786 327712
rect 129826 327700 129832 327712
rect 129884 327740 129890 327752
rect 251818 327740 251824 327752
rect 129884 327712 251824 327740
rect 129884 327700 129890 327712
rect 251818 327700 251824 327712
rect 251876 327700 251882 327752
rect 162118 327088 162124 327140
rect 162176 327128 162182 327140
rect 212626 327128 212632 327140
rect 162176 327100 212632 327128
rect 162176 327088 162182 327100
rect 212626 327088 212632 327100
rect 212684 327088 212690 327140
rect 85390 327020 85396 327072
rect 85448 327060 85454 327072
rect 88334 327060 88340 327072
rect 85448 327032 88340 327060
rect 85448 327020 85454 327032
rect 88334 327020 88340 327032
rect 88392 327020 88398 327072
rect 103514 327020 103520 327072
rect 103572 327060 103578 327072
rect 110690 327060 110696 327072
rect 103572 327032 110696 327060
rect 103572 327020 103578 327032
rect 110690 327020 110696 327032
rect 110748 327020 110754 327072
rect 114002 325728 114008 325780
rect 114060 325768 114066 325780
rect 249058 325768 249064 325780
rect 114060 325740 249064 325768
rect 114060 325728 114066 325740
rect 249058 325728 249064 325740
rect 249116 325728 249122 325780
rect 61378 325660 61384 325712
rect 61436 325700 61442 325712
rect 61436 325672 67634 325700
rect 61436 325660 61442 325672
rect 67606 325632 67634 325672
rect 110690 325660 110696 325712
rect 110748 325700 110754 325712
rect 270586 325700 270592 325712
rect 110748 325672 270592 325700
rect 110748 325660 110754 325672
rect 270586 325660 270592 325672
rect 270644 325660 270650 325712
rect 67726 325632 67732 325644
rect 67606 325604 67732 325632
rect 67726 325592 67732 325604
rect 67784 325592 67790 325644
rect 108482 324980 108488 325032
rect 108540 325020 108546 325032
rect 125594 325020 125600 325032
rect 108540 324992 125600 325020
rect 108540 324980 108546 324992
rect 125594 324980 125600 324992
rect 125652 325020 125658 325032
rect 259638 325020 259644 325032
rect 125652 324992 259644 325020
rect 125652 324980 125658 324992
rect 259638 324980 259644 324992
rect 259696 324980 259702 325032
rect 67726 324912 67732 324964
rect 67784 324952 67790 324964
rect 252738 324952 252744 324964
rect 67784 324924 252744 324952
rect 67784 324912 67790 324924
rect 252738 324912 252744 324924
rect 252796 324912 252802 324964
rect 113818 323552 113824 323604
rect 113876 323592 113882 323604
rect 121638 323592 121644 323604
rect 113876 323564 121644 323592
rect 113876 323552 113882 323564
rect 121638 323552 121644 323564
rect 121696 323592 121702 323604
rect 262214 323592 262220 323604
rect 121696 323564 262220 323592
rect 121696 323552 121702 323564
rect 262214 323552 262220 323564
rect 262272 323552 262278 323604
rect 256786 322980 256792 322992
rect 59832 322952 256792 322980
rect 53558 322872 53564 322924
rect 53616 322912 53622 322924
rect 59354 322912 59360 322924
rect 53616 322884 59360 322912
rect 53616 322872 53622 322884
rect 59354 322872 59360 322884
rect 59412 322912 59418 322924
rect 59832 322912 59860 322952
rect 256786 322940 256792 322952
rect 256844 322940 256850 322992
rect 59412 322884 59860 322912
rect 59412 322872 59418 322884
rect 89438 322872 89444 322924
rect 89496 322912 89502 322924
rect 93854 322912 93860 322924
rect 89496 322884 93860 322912
rect 89496 322872 89502 322884
rect 93854 322872 93860 322884
rect 93912 322872 93918 322924
rect 78490 322736 78496 322788
rect 78548 322776 78554 322788
rect 84378 322776 84384 322788
rect 78548 322748 84384 322776
rect 78548 322736 78554 322748
rect 84378 322736 84384 322748
rect 84436 322736 84442 322788
rect 180058 321648 180064 321700
rect 180116 321688 180122 321700
rect 245010 321688 245016 321700
rect 180116 321660 245016 321688
rect 180116 321648 180122 321660
rect 245010 321648 245016 321660
rect 245068 321648 245074 321700
rect 137370 321580 137376 321632
rect 137428 321620 137434 321632
rect 254210 321620 254216 321632
rect 137428 321592 254216 321620
rect 137428 321580 137434 321592
rect 254210 321580 254216 321592
rect 254268 321580 254274 321632
rect 127066 321512 127072 321564
rect 127124 321552 127130 321564
rect 264238 321552 264244 321564
rect 127124 321524 264244 321552
rect 127124 321512 127130 321524
rect 264238 321512 264244 321524
rect 264296 321512 264302 321564
rect 263778 321036 263784 321088
rect 263836 321076 263842 321088
rect 264238 321076 264244 321088
rect 263836 321048 264244 321076
rect 263836 321036 263842 321048
rect 264238 321036 264244 321048
rect 264296 321036 264302 321088
rect 92198 320900 92204 320952
rect 92256 320940 92262 320952
rect 123018 320940 123024 320952
rect 92256 320912 123024 320940
rect 92256 320900 92262 320912
rect 123018 320900 123024 320912
rect 123076 320940 123082 320952
rect 125318 320940 125324 320952
rect 123076 320912 125324 320940
rect 123076 320900 123082 320912
rect 125318 320900 125324 320912
rect 125376 320900 125382 320952
rect 64598 320832 64604 320884
rect 64656 320872 64662 320884
rect 75178 320872 75184 320884
rect 64656 320844 75184 320872
rect 64656 320832 64662 320844
rect 75178 320832 75184 320844
rect 75236 320832 75242 320884
rect 89806 320832 89812 320884
rect 89864 320872 89870 320884
rect 127066 320872 127072 320884
rect 89864 320844 127072 320872
rect 89864 320832 89870 320844
rect 127066 320832 127072 320844
rect 127124 320832 127130 320884
rect 53098 320152 53104 320204
rect 53156 320192 53162 320204
rect 63494 320192 63500 320204
rect 53156 320164 63500 320192
rect 53156 320152 53162 320164
rect 63494 320152 63500 320164
rect 63552 320192 63558 320204
rect 64138 320192 64144 320204
rect 63552 320164 64144 320192
rect 63552 320152 63558 320164
rect 64138 320152 64144 320164
rect 64196 320152 64202 320204
rect 125318 320152 125324 320204
rect 125376 320192 125382 320204
rect 261018 320192 261024 320204
rect 125376 320164 261024 320192
rect 125376 320152 125382 320164
rect 261018 320152 261024 320164
rect 261076 320152 261082 320204
rect 98362 319472 98368 319524
rect 98420 319512 98426 319524
rect 106274 319512 106280 319524
rect 98420 319484 106280 319512
rect 98420 319472 98426 319484
rect 106274 319472 106280 319484
rect 106332 319472 106338 319524
rect 63494 319404 63500 319456
rect 63552 319444 63558 319456
rect 251910 319444 251916 319456
rect 63552 319416 251916 319444
rect 63552 319404 63558 319416
rect 251910 319404 251916 319416
rect 251968 319404 251974 319456
rect 68462 318588 68468 318640
rect 68520 318628 68526 318640
rect 69106 318628 69112 318640
rect 68520 318600 69112 318628
rect 68520 318588 68526 318600
rect 69106 318588 69112 318600
rect 69164 318588 69170 318640
rect 95878 317432 95884 317484
rect 95936 317472 95942 317484
rect 116578 317472 116584 317484
rect 95936 317444 116584 317472
rect 95936 317432 95942 317444
rect 116578 317432 116584 317444
rect 116636 317432 116642 317484
rect 74534 316888 74540 316940
rect 74592 316928 74598 316940
rect 81526 316928 81532 316940
rect 74592 316900 81532 316928
rect 74592 316888 74598 316900
rect 81526 316888 81532 316900
rect 81584 316888 81590 316940
rect 99282 316752 99288 316804
rect 99340 316792 99346 316804
rect 117406 316792 117412 316804
rect 99340 316764 117412 316792
rect 99340 316752 99346 316764
rect 117406 316752 117412 316764
rect 117464 316792 117470 316804
rect 131022 316792 131028 316804
rect 117464 316764 131028 316792
rect 117464 316752 117470 316764
rect 131022 316752 131028 316764
rect 131080 316752 131086 316804
rect 82906 316684 82912 316736
rect 82964 316724 82970 316736
rect 124306 316724 124312 316736
rect 82964 316696 124312 316724
rect 82964 316684 82970 316696
rect 124306 316684 124312 316696
rect 124364 316724 124370 316736
rect 125410 316724 125416 316736
rect 124364 316696 125416 316724
rect 124364 316684 124370 316696
rect 125410 316684 125416 316696
rect 125468 316684 125474 316736
rect 185578 316072 185584 316124
rect 185636 316112 185642 316124
rect 267734 316112 267740 316124
rect 185636 316084 267740 316112
rect 185636 316072 185642 316084
rect 267734 316072 267740 316084
rect 267792 316072 267798 316124
rect 131022 316004 131028 316056
rect 131080 316044 131086 316056
rect 250530 316044 250536 316056
rect 131080 316016 250536 316044
rect 131080 316004 131086 316016
rect 250530 316004 250536 316016
rect 250588 316004 250594 316056
rect 273346 315460 273352 315512
rect 273404 315500 273410 315512
rect 273898 315500 273904 315512
rect 273404 315472 273904 315500
rect 273404 315460 273410 315472
rect 273898 315460 273904 315472
rect 273956 315460 273962 315512
rect 97902 315256 97908 315308
rect 97960 315296 97966 315308
rect 273346 315296 273352 315308
rect 97960 315268 273352 315296
rect 97960 315256 97966 315268
rect 273346 315256 273352 315268
rect 273404 315256 273410 315308
rect 96614 314644 96620 314696
rect 96672 314684 96678 314696
rect 97902 314684 97908 314696
rect 96672 314656 97908 314684
rect 96672 314644 96678 314656
rect 97902 314644 97908 314656
rect 97960 314644 97966 314696
rect 151262 314644 151268 314696
rect 151320 314684 151326 314696
rect 247678 314684 247684 314696
rect 151320 314656 247684 314684
rect 151320 314644 151326 314656
rect 247678 314644 247684 314656
rect 247736 314644 247742 314696
rect 186314 313352 186320 313404
rect 186372 313392 186378 313404
rect 265066 313392 265072 313404
rect 186372 313364 265072 313392
rect 186372 313352 186378 313364
rect 265066 313352 265072 313364
rect 265124 313352 265130 313404
rect 105630 313284 105636 313336
rect 105688 313324 105694 313336
rect 106182 313324 106188 313336
rect 105688 313296 106188 313324
rect 105688 313284 105694 313296
rect 106182 313284 106188 313296
rect 106240 313324 106246 313336
rect 252830 313324 252836 313336
rect 106240 313296 252836 313324
rect 106240 313284 106246 313296
rect 252830 313284 252836 313296
rect 252888 313284 252894 313336
rect 3418 313216 3424 313268
rect 3476 313256 3482 313268
rect 7558 313256 7564 313268
rect 3476 313228 7564 313256
rect 3476 313216 3482 313228
rect 7558 313216 7564 313228
rect 7616 313216 7622 313268
rect 67266 312536 67272 312588
rect 67324 312576 67330 312588
rect 258166 312576 258172 312588
rect 67324 312548 258172 312576
rect 67324 312536 67330 312548
rect 258166 312536 258172 312548
rect 258224 312536 258230 312588
rect 187142 311856 187148 311908
rect 187200 311896 187206 311908
rect 263870 311896 263876 311908
rect 187200 311868 263876 311896
rect 187200 311856 187206 311868
rect 263870 311856 263876 311868
rect 263928 311856 263934 311908
rect 278038 311856 278044 311908
rect 278096 311896 278102 311908
rect 580166 311896 580172 311908
rect 278096 311868 580172 311896
rect 278096 311856 278102 311868
rect 580166 311856 580172 311868
rect 580224 311856 580230 311908
rect 109678 311108 109684 311160
rect 109736 311148 109742 311160
rect 134058 311148 134064 311160
rect 109736 311120 134064 311148
rect 109736 311108 109742 311120
rect 134058 311108 134064 311120
rect 134116 311148 134122 311160
rect 259546 311148 259552 311160
rect 134116 311120 259552 311148
rect 134116 311108 134122 311120
rect 259546 311108 259552 311120
rect 259604 311108 259610 311160
rect 189810 310496 189816 310548
rect 189868 310536 189874 310548
rect 261110 310536 261116 310548
rect 189868 310508 261116 310536
rect 189868 310496 189874 310508
rect 261110 310496 261116 310508
rect 261168 310496 261174 310548
rect 104158 310428 104164 310480
rect 104216 310468 104222 310480
rect 108390 310468 108396 310480
rect 104216 310440 108396 310468
rect 104216 310428 104222 310440
rect 108390 310428 108396 310440
rect 108448 310428 108454 310480
rect 97718 309748 97724 309800
rect 97776 309788 97782 309800
rect 117406 309788 117412 309800
rect 97776 309760 117412 309788
rect 97776 309748 97782 309760
rect 117406 309748 117412 309760
rect 117464 309748 117470 309800
rect 148318 309204 148324 309256
rect 148376 309244 148382 309256
rect 238018 309244 238024 309256
rect 148376 309216 238024 309244
rect 148376 309204 148382 309216
rect 238018 309204 238024 309216
rect 238076 309204 238082 309256
rect 122742 309136 122748 309188
rect 122800 309176 122806 309188
rect 220170 309176 220176 309188
rect 122800 309148 220176 309176
rect 122800 309136 122806 309148
rect 220170 309136 220176 309148
rect 220228 309136 220234 309188
rect 67358 309068 67364 309120
rect 67416 309108 67422 309120
rect 186314 309108 186320 309120
rect 67416 309080 186320 309108
rect 67416 309068 67422 309080
rect 186314 309068 186320 309080
rect 186372 309068 186378 309120
rect 188430 307844 188436 307896
rect 188488 307884 188494 307896
rect 254118 307884 254124 307896
rect 188488 307856 254124 307884
rect 188488 307844 188494 307856
rect 254118 307844 254124 307856
rect 254176 307844 254182 307896
rect 22002 307776 22008 307828
rect 22060 307816 22066 307828
rect 202414 307816 202420 307828
rect 22060 307788 202420 307816
rect 22060 307776 22066 307788
rect 202414 307776 202420 307788
rect 202472 307776 202478 307828
rect 202506 307776 202512 307828
rect 202564 307816 202570 307828
rect 262398 307816 262404 307828
rect 202564 307788 262404 307816
rect 202564 307776 202570 307788
rect 262398 307776 262404 307788
rect 262456 307776 262462 307828
rect 182910 306416 182916 306468
rect 182968 306456 182974 306468
rect 210418 306456 210424 306468
rect 182968 306428 210424 306456
rect 182968 306416 182974 306428
rect 210418 306416 210424 306428
rect 210476 306416 210482 306468
rect 175918 306348 175924 306400
rect 175976 306388 175982 306400
rect 241054 306388 241060 306400
rect 175976 306360 241060 306388
rect 175976 306348 175982 306360
rect 241054 306348 241060 306360
rect 241112 306348 241118 306400
rect 65886 305600 65892 305652
rect 65944 305640 65950 305652
rect 151262 305640 151268 305652
rect 65944 305612 151268 305640
rect 65944 305600 65950 305612
rect 151262 305600 151268 305612
rect 151320 305600 151326 305652
rect 232498 305600 232504 305652
rect 232556 305640 232562 305652
rect 269206 305640 269212 305652
rect 232556 305612 269212 305640
rect 232556 305600 232562 305612
rect 269206 305600 269212 305612
rect 269264 305600 269270 305652
rect 192570 305056 192576 305108
rect 192628 305096 192634 305108
rect 255498 305096 255504 305108
rect 192628 305068 255504 305096
rect 192628 305056 192634 305068
rect 255498 305056 255504 305068
rect 255556 305056 255562 305108
rect 3234 304988 3240 305040
rect 3292 305028 3298 305040
rect 32398 305028 32404 305040
rect 3292 305000 32404 305028
rect 3292 304988 3298 305000
rect 32398 304988 32404 305000
rect 32456 304988 32462 305040
rect 152458 304988 152464 305040
rect 152516 305028 152522 305040
rect 216766 305028 216772 305040
rect 152516 305000 216772 305028
rect 152516 304988 152522 305000
rect 216766 304988 216772 305000
rect 216824 304988 216830 305040
rect 113910 304308 113916 304360
rect 113968 304348 113974 304360
rect 123478 304348 123484 304360
rect 113968 304320 123484 304348
rect 113968 304308 113974 304320
rect 123478 304308 123484 304320
rect 123536 304308 123542 304360
rect 85574 304240 85580 304292
rect 85632 304280 85638 304292
rect 95878 304280 95884 304292
rect 85632 304252 95884 304280
rect 85632 304240 85638 304252
rect 95878 304240 95884 304252
rect 95936 304240 95942 304292
rect 96430 304240 96436 304292
rect 96488 304280 96494 304292
rect 108482 304280 108488 304292
rect 96488 304252 108488 304280
rect 96488 304240 96494 304252
rect 108482 304240 108488 304252
rect 108540 304240 108546 304292
rect 114094 304240 114100 304292
rect 114152 304280 114158 304292
rect 125502 304280 125508 304292
rect 114152 304252 125508 304280
rect 114152 304240 114158 304252
rect 125502 304240 125508 304252
rect 125560 304280 125566 304292
rect 135990 304280 135996 304292
rect 125560 304252 135996 304280
rect 125560 304240 125566 304252
rect 135990 304240 135996 304252
rect 136048 304240 136054 304292
rect 246298 304240 246304 304292
rect 246356 304280 246362 304292
rect 251266 304280 251272 304292
rect 246356 304252 251272 304280
rect 246356 304240 246362 304252
rect 251266 304240 251272 304252
rect 251324 304240 251330 304292
rect 250438 304036 250444 304088
rect 250496 304076 250502 304088
rect 253934 304076 253940 304088
rect 250496 304048 253940 304076
rect 250496 304036 250502 304048
rect 253934 304036 253940 304048
rect 253992 304036 253998 304088
rect 142798 303764 142804 303816
rect 142856 303804 142862 303816
rect 216122 303804 216128 303816
rect 142856 303776 216128 303804
rect 142856 303764 142862 303776
rect 216122 303764 216128 303776
rect 216180 303764 216186 303816
rect 170398 303696 170404 303748
rect 170456 303736 170462 303748
rect 214190 303736 214196 303748
rect 170456 303708 214196 303736
rect 170456 303696 170462 303708
rect 214190 303696 214196 303708
rect 214248 303696 214254 303748
rect 215294 303696 215300 303748
rect 215352 303736 215358 303748
rect 228910 303736 228916 303748
rect 215352 303708 228916 303736
rect 215352 303696 215358 303708
rect 228910 303696 228916 303708
rect 228968 303696 228974 303748
rect 213914 303628 213920 303680
rect 213972 303668 213978 303680
rect 229554 303668 229560 303680
rect 213972 303640 229560 303668
rect 213972 303628 213978 303640
rect 229554 303628 229560 303640
rect 229612 303628 229618 303680
rect 233878 303628 233884 303680
rect 233936 303668 233942 303680
rect 237834 303668 237840 303680
rect 233936 303640 237840 303668
rect 233936 303628 233942 303640
rect 237834 303628 237840 303640
rect 237892 303628 237898 303680
rect 240042 303628 240048 303680
rect 240100 303668 240106 303680
rect 250622 303668 250628 303680
rect 240100 303640 250628 303668
rect 240100 303628 240106 303640
rect 250622 303628 250628 303640
rect 250680 303628 250686 303680
rect 149054 303560 149060 303612
rect 149112 303600 149118 303612
rect 240686 303600 240692 303612
rect 149112 303572 240692 303600
rect 149112 303560 149118 303572
rect 240686 303560 240692 303572
rect 240744 303600 240750 303612
rect 247402 303600 247408 303612
rect 240744 303572 247408 303600
rect 240744 303560 240750 303572
rect 247402 303560 247408 303572
rect 247460 303560 247466 303612
rect 141602 302880 141608 302932
rect 141660 302920 141666 302932
rect 149054 302920 149060 302932
rect 141660 302892 149060 302920
rect 141660 302880 141666 302892
rect 149054 302880 149060 302892
rect 149112 302880 149118 302932
rect 245010 302880 245016 302932
rect 245068 302920 245074 302932
rect 252738 302920 252744 302932
rect 245068 302892 252744 302920
rect 245068 302880 245074 302892
rect 252738 302880 252744 302892
rect 252796 302880 252802 302932
rect 256878 302880 256884 302932
rect 256936 302920 256942 302932
rect 274726 302920 274732 302932
rect 256936 302892 274732 302920
rect 256936 302880 256942 302892
rect 274726 302880 274732 302892
rect 274784 302880 274790 302932
rect 250530 302404 250536 302456
rect 250588 302444 250594 302456
rect 256878 302444 256884 302456
rect 250588 302416 256884 302444
rect 250588 302404 250594 302416
rect 256878 302404 256884 302416
rect 256936 302404 256942 302456
rect 77294 302200 77300 302252
rect 77352 302240 77358 302252
rect 78490 302240 78496 302252
rect 77352 302212 78496 302240
rect 77352 302200 77358 302212
rect 78490 302200 78496 302212
rect 78548 302240 78554 302252
rect 131850 302240 131856 302252
rect 78548 302212 131856 302240
rect 78548 302200 78554 302212
rect 131850 302200 131856 302212
rect 131908 302200 131914 302252
rect 191374 302200 191380 302252
rect 191432 302240 191438 302252
rect 211062 302240 211068 302252
rect 191432 302212 211068 302240
rect 191432 302200 191438 302212
rect 211062 302200 211068 302212
rect 211120 302200 211126 302252
rect 255958 302132 255964 302184
rect 256016 302172 256022 302184
rect 259730 302172 259736 302184
rect 256016 302144 259736 302172
rect 256016 302132 256022 302144
rect 259730 302132 259736 302144
rect 259788 302132 259794 302184
rect 249058 301860 249064 301912
rect 249116 301900 249122 301912
rect 255682 301900 255688 301912
rect 249116 301872 255688 301900
rect 249116 301860 249122 301872
rect 255682 301860 255688 301872
rect 255740 301860 255746 301912
rect 79962 301452 79968 301504
rect 80020 301492 80026 301504
rect 103606 301492 103612 301504
rect 80020 301464 103612 301492
rect 80020 301452 80026 301464
rect 103606 301452 103612 301464
rect 103664 301492 103670 301504
rect 189810 301492 189816 301504
rect 103664 301464 189816 301492
rect 103664 301452 103670 301464
rect 189810 301452 189816 301464
rect 189868 301452 189874 301504
rect 193306 301112 193312 301164
rect 193364 301152 193370 301164
rect 193364 301124 200114 301152
rect 193364 301112 193370 301124
rect 186286 301056 195974 301084
rect 186286 300948 186314 301056
rect 195422 300976 195428 301028
rect 195480 300976 195486 301028
rect 180766 300920 186314 300948
rect 178678 300840 178684 300892
rect 178736 300880 178742 300892
rect 180766 300880 180794 300920
rect 178736 300852 180794 300880
rect 178736 300840 178742 300852
rect 190362 300772 190368 300824
rect 190420 300812 190426 300824
rect 195440 300812 195468 300976
rect 195946 300948 195974 301056
rect 200086 301016 200114 301124
rect 211982 301016 211988 301028
rect 200086 300988 211988 301016
rect 211982 300976 211988 300988
rect 212040 300976 212046 301028
rect 208854 300948 208860 300960
rect 195946 300920 208860 300948
rect 208854 300908 208860 300920
rect 208912 300908 208918 300960
rect 219434 300908 219440 300960
rect 219492 300908 219498 300960
rect 244274 300908 244280 300960
rect 244332 300908 244338 300960
rect 190420 300784 195468 300812
rect 219452 300812 219480 300908
rect 244292 300880 244320 300908
rect 270494 300880 270500 300892
rect 244292 300852 270500 300880
rect 270494 300840 270500 300852
rect 270552 300840 270558 300892
rect 219452 300784 229094 300812
rect 190420 300772 190426 300784
rect 179322 300160 179328 300212
rect 179380 300200 179386 300212
rect 190454 300200 190460 300212
rect 179380 300172 190460 300200
rect 179380 300160 179386 300172
rect 190454 300160 190460 300172
rect 190512 300160 190518 300212
rect 126422 300092 126428 300144
rect 126480 300132 126486 300144
rect 190546 300132 190552 300144
rect 126480 300104 190552 300132
rect 126480 300092 126486 300104
rect 190546 300092 190552 300104
rect 190604 300092 190610 300144
rect 229066 300132 229094 300784
rect 252922 300132 252928 300144
rect 229066 300104 252928 300132
rect 252922 300092 252928 300104
rect 252980 300092 252986 300144
rect 252830 299820 252836 299872
rect 252888 299860 252894 299872
rect 253106 299860 253112 299872
rect 252888 299832 253112 299860
rect 252888 299820 252894 299832
rect 253106 299820 253112 299832
rect 253164 299820 253170 299872
rect 56502 299480 56508 299532
rect 56560 299520 56566 299532
rect 159450 299520 159456 299532
rect 56560 299492 159456 299520
rect 56560 299480 56566 299492
rect 159450 299480 159456 299492
rect 159508 299480 159514 299532
rect 255406 299480 255412 299532
rect 255464 299520 255470 299532
rect 287054 299520 287060 299532
rect 255464 299492 287060 299520
rect 255464 299480 255470 299492
rect 287054 299480 287060 299492
rect 287112 299480 287118 299532
rect 146938 299412 146944 299464
rect 146996 299452 147002 299464
rect 191006 299452 191012 299464
rect 146996 299424 191012 299452
rect 146996 299412 147002 299424
rect 191006 299412 191012 299424
rect 191064 299412 191070 299464
rect 580902 299412 580908 299464
rect 580960 299452 580966 299464
rect 583570 299452 583576 299464
rect 580960 299424 583576 299452
rect 580960 299412 580966 299424
rect 583570 299412 583576 299424
rect 583628 299412 583634 299464
rect 255314 298120 255320 298172
rect 255372 298160 255378 298172
rect 288434 298160 288440 298172
rect 255372 298132 288440 298160
rect 255372 298120 255378 298132
rect 288434 298120 288440 298132
rect 288492 298120 288498 298172
rect 160094 298052 160100 298104
rect 160152 298092 160158 298104
rect 161290 298092 161296 298104
rect 160152 298064 161296 298092
rect 160152 298052 160158 298064
rect 161290 298052 161296 298064
rect 161348 298092 161354 298104
rect 191098 298092 191104 298104
rect 161348 298064 191104 298092
rect 161348 298052 161354 298064
rect 191098 298052 191104 298064
rect 191156 298052 191162 298104
rect 255314 297984 255320 298036
rect 255372 298024 255378 298036
rect 255498 298024 255504 298036
rect 255372 297996 255504 298024
rect 255372 297984 255378 297996
rect 255498 297984 255504 297996
rect 255556 297984 255562 298036
rect 255590 296760 255596 296812
rect 255648 296800 255654 296812
rect 260926 296800 260932 296812
rect 255648 296772 260932 296800
rect 255648 296760 255654 296772
rect 260926 296760 260932 296772
rect 260984 296760 260990 296812
rect 82814 296692 82820 296744
rect 82872 296732 82878 296744
rect 84010 296732 84016 296744
rect 82872 296704 84016 296732
rect 82872 296692 82878 296704
rect 84010 296692 84016 296704
rect 84068 296732 84074 296744
rect 184198 296732 184204 296744
rect 84068 296704 184204 296732
rect 84068 296692 84074 296704
rect 184198 296692 184204 296704
rect 184256 296692 184262 296744
rect 255498 296692 255504 296744
rect 255556 296732 255562 296744
rect 282914 296732 282920 296744
rect 255556 296704 282920 296732
rect 255556 296692 255562 296704
rect 282914 296692 282920 296704
rect 282972 296692 282978 296744
rect 124122 295944 124128 295996
rect 124180 295984 124186 295996
rect 192478 295984 192484 295996
rect 124180 295956 192484 295984
rect 124180 295944 124186 295956
rect 192478 295944 192484 295956
rect 192536 295944 192542 295996
rect 256050 295468 256056 295520
rect 256108 295508 256114 295520
rect 258350 295508 258356 295520
rect 256108 295480 258356 295508
rect 256108 295468 256114 295480
rect 258350 295468 258356 295480
rect 258408 295468 258414 295520
rect 69658 295332 69664 295384
rect 69716 295372 69722 295384
rect 156598 295372 156604 295384
rect 69716 295344 156604 295372
rect 69716 295332 69722 295344
rect 156598 295332 156604 295344
rect 156656 295372 156662 295384
rect 190454 295372 190460 295384
rect 156656 295344 190460 295372
rect 156656 295332 156662 295344
rect 190454 295332 190460 295344
rect 190512 295332 190518 295384
rect 255498 295332 255504 295384
rect 255556 295372 255562 295384
rect 284386 295372 284392 295384
rect 255556 295344 284392 295372
rect 255556 295332 255562 295344
rect 284386 295332 284392 295344
rect 284444 295332 284450 295384
rect 120166 295264 120172 295316
rect 120224 295304 120230 295316
rect 190546 295304 190552 295316
rect 120224 295276 190552 295304
rect 120224 295264 120230 295276
rect 190546 295264 190552 295276
rect 190604 295264 190610 295316
rect 180242 294584 180248 294636
rect 180300 294624 180306 294636
rect 193306 294624 193312 294636
rect 180300 294596 193312 294624
rect 180300 294584 180306 294596
rect 193306 294584 193312 294596
rect 193364 294584 193370 294636
rect 117222 294040 117228 294092
rect 117280 294080 117286 294092
rect 120166 294080 120172 294092
rect 117280 294052 120172 294080
rect 117280 294040 117286 294052
rect 120166 294040 120172 294052
rect 120224 294040 120230 294092
rect 255590 294040 255596 294092
rect 255648 294080 255654 294092
rect 267918 294080 267924 294092
rect 255648 294052 267924 294080
rect 255648 294040 255654 294052
rect 267918 294040 267924 294052
rect 267976 294040 267982 294092
rect 69566 293972 69572 294024
rect 69624 294012 69630 294024
rect 70210 294012 70216 294024
rect 69624 293984 70216 294012
rect 69624 293972 69630 293984
rect 70210 293972 70216 293984
rect 70268 294012 70274 294024
rect 126514 294012 126520 294024
rect 70268 293984 126520 294012
rect 70268 293972 70274 293984
rect 126514 293972 126520 293984
rect 126572 293972 126578 294024
rect 255498 293972 255504 294024
rect 255556 294012 255562 294024
rect 273254 294012 273260 294024
rect 255556 293984 273260 294012
rect 255556 293972 255562 293984
rect 273254 293972 273260 293984
rect 273312 293972 273318 294024
rect 59170 293292 59176 293344
rect 59228 293332 59234 293344
rect 87598 293332 87604 293344
rect 59228 293304 87604 293332
rect 59228 293292 59234 293304
rect 87598 293292 87604 293304
rect 87656 293292 87662 293344
rect 84562 293224 84568 293276
rect 84620 293264 84626 293276
rect 93026 293264 93032 293276
rect 84620 293236 93032 293264
rect 84620 293224 84626 293236
rect 93026 293224 93032 293236
rect 93084 293264 93090 293276
rect 124122 293264 124128 293276
rect 93084 293236 124128 293264
rect 93084 293224 93090 293236
rect 124122 293224 124128 293236
rect 124180 293224 124186 293276
rect 169018 293224 169024 293276
rect 169076 293264 169082 293276
rect 192570 293264 192576 293276
rect 169076 293236 192576 293264
rect 169076 293224 169082 293236
rect 192570 293224 192576 293236
rect 192628 293224 192634 293276
rect 255498 293224 255504 293276
rect 255556 293264 255562 293276
rect 270586 293264 270592 293276
rect 255556 293236 270592 293264
rect 255556 293224 255562 293236
rect 270586 293224 270592 293236
rect 270644 293224 270650 293276
rect 71682 292612 71688 292664
rect 71740 292652 71746 292664
rect 71958 292652 71964 292664
rect 71740 292624 71964 292652
rect 71740 292612 71746 292624
rect 71958 292612 71964 292624
rect 72016 292612 72022 292664
rect 3418 292544 3424 292596
rect 3476 292584 3482 292596
rect 18690 292584 18696 292596
rect 3476 292556 18696 292584
rect 3476 292544 3482 292556
rect 18690 292544 18696 292556
rect 18748 292544 18754 292596
rect 36538 292544 36544 292596
rect 36596 292584 36602 292596
rect 58986 292584 58992 292596
rect 36596 292556 58992 292584
rect 36596 292544 36602 292556
rect 58986 292544 58992 292556
rect 59044 292584 59050 292596
rect 59170 292584 59176 292596
rect 59044 292556 59176 292584
rect 59044 292544 59050 292556
rect 59170 292544 59176 292556
rect 59228 292544 59234 292596
rect 122098 292544 122104 292596
rect 122156 292584 122162 292596
rect 193122 292584 193128 292596
rect 122156 292556 193128 292584
rect 122156 292544 122162 292556
rect 193122 292544 193128 292556
rect 193180 292544 193186 292596
rect 255590 292544 255596 292596
rect 255648 292584 255654 292596
rect 280154 292584 280160 292596
rect 255648 292556 280160 292584
rect 255648 292544 255654 292556
rect 280154 292544 280160 292556
rect 280212 292544 280218 292596
rect 101398 292476 101404 292528
rect 101456 292516 101462 292528
rect 193214 292516 193220 292528
rect 101456 292488 193220 292516
rect 101456 292476 101462 292488
rect 193214 292476 193220 292488
rect 193272 292476 193278 292528
rect 101490 291796 101496 291848
rect 101548 291836 101554 291848
rect 114002 291836 114008 291848
rect 101548 291808 114008 291836
rect 101548 291796 101554 291808
rect 114002 291796 114008 291808
rect 114060 291796 114066 291848
rect 255682 291796 255688 291848
rect 255740 291836 255746 291848
rect 269114 291836 269120 291848
rect 255740 291808 269120 291836
rect 255740 291796 255746 291808
rect 269114 291796 269120 291808
rect 269172 291796 269178 291848
rect 91462 291184 91468 291236
rect 91520 291224 91526 291236
rect 97258 291224 97264 291236
rect 91520 291196 97264 291224
rect 91520 291184 91526 291196
rect 97258 291184 97264 291196
rect 97316 291184 97322 291236
rect 255498 291184 255504 291236
rect 255556 291224 255562 291236
rect 262306 291224 262312 291236
rect 255556 291196 262312 291224
rect 255556 291184 255562 291196
rect 262306 291184 262312 291196
rect 262364 291184 262370 291236
rect 255498 290980 255504 291032
rect 255556 291020 255562 291032
rect 259638 291020 259644 291032
rect 255556 290992 259644 291020
rect 255556 290980 255562 290992
rect 259638 290980 259644 290992
rect 259696 290980 259702 291032
rect 82998 289892 83004 289944
rect 83056 289932 83062 289944
rect 84102 289932 84108 289944
rect 83056 289904 84108 289932
rect 83056 289892 83062 289904
rect 84102 289892 84108 289904
rect 84160 289932 84166 289944
rect 103514 289932 103520 289944
rect 84160 289904 103520 289932
rect 84160 289892 84166 289904
rect 103514 289892 103520 289904
rect 103572 289892 103578 289944
rect 94498 289824 94504 289876
rect 94556 289864 94562 289876
rect 193214 289864 193220 289876
rect 94556 289836 193220 289864
rect 94556 289824 94562 289836
rect 193214 289824 193220 289836
rect 193272 289824 193278 289876
rect 255498 289756 255504 289808
rect 255556 289796 255562 289808
rect 262214 289796 262220 289808
rect 255556 289768 262220 289796
rect 255556 289756 255562 289768
rect 262214 289756 262220 289768
rect 262272 289756 262278 289808
rect 82722 289076 82728 289128
rect 82780 289116 82786 289128
rect 94498 289116 94504 289128
rect 82780 289088 94504 289116
rect 82780 289076 82786 289088
rect 94498 289076 94504 289088
rect 94556 289076 94562 289128
rect 45370 288464 45376 288516
rect 45428 288504 45434 288516
rect 79318 288504 79324 288516
rect 45428 288476 79324 288504
rect 45428 288464 45434 288476
rect 79318 288464 79324 288476
rect 79376 288504 79382 288516
rect 79594 288504 79600 288516
rect 79376 288476 79600 288504
rect 79376 288464 79382 288476
rect 79594 288464 79600 288476
rect 79652 288464 79658 288516
rect 95602 288464 95608 288516
rect 95660 288504 95666 288516
rect 96430 288504 96436 288516
rect 95660 288476 96436 288504
rect 95660 288464 95666 288476
rect 96430 288464 96436 288476
rect 96488 288504 96494 288516
rect 112530 288504 112536 288516
rect 96488 288476 112536 288504
rect 96488 288464 96494 288476
rect 112530 288464 112536 288476
rect 112588 288464 112594 288516
rect 142982 288464 142988 288516
rect 143040 288504 143046 288516
rect 186222 288504 186228 288516
rect 143040 288476 186228 288504
rect 143040 288464 143046 288476
rect 186222 288464 186228 288476
rect 186280 288504 186286 288516
rect 191006 288504 191012 288516
rect 186280 288476 191012 288504
rect 186280 288464 186286 288476
rect 191006 288464 191012 288476
rect 191064 288464 191070 288516
rect 78582 288396 78588 288448
rect 78640 288436 78646 288448
rect 168282 288436 168288 288448
rect 78640 288408 168288 288436
rect 78640 288396 78646 288408
rect 168282 288396 168288 288408
rect 168340 288396 168346 288448
rect 18598 288328 18604 288380
rect 18656 288368 18662 288380
rect 71038 288368 71044 288380
rect 18656 288340 71044 288368
rect 18656 288328 18662 288340
rect 71038 288328 71044 288340
rect 71096 288328 71102 288380
rect 168300 288368 168328 288396
rect 180058 288368 180064 288380
rect 168300 288340 180064 288368
rect 180058 288328 180064 288340
rect 180116 288328 180122 288380
rect 255498 288328 255504 288380
rect 255556 288368 255562 288380
rect 262398 288368 262404 288380
rect 255556 288340 262404 288368
rect 255556 288328 255562 288340
rect 262398 288328 262404 288340
rect 262456 288328 262462 288380
rect 127618 287648 127624 287700
rect 127676 287688 127682 287700
rect 137370 287688 137376 287700
rect 127676 287660 137376 287688
rect 127676 287648 127682 287660
rect 137370 287648 137376 287660
rect 137428 287648 137434 287700
rect 159450 287648 159456 287700
rect 159508 287688 159514 287700
rect 166902 287688 166908 287700
rect 159508 287660 166908 287688
rect 159508 287648 159514 287660
rect 166902 287648 166908 287660
rect 166960 287648 166966 287700
rect 95142 287104 95148 287156
rect 95200 287144 95206 287156
rect 127618 287144 127624 287156
rect 95200 287116 127624 287144
rect 95200 287104 95206 287116
rect 127618 287104 127624 287116
rect 127676 287104 127682 287156
rect 60458 287036 60464 287088
rect 60516 287076 60522 287088
rect 79410 287076 79416 287088
rect 60516 287048 79416 287076
rect 60516 287036 60522 287048
rect 79410 287036 79416 287048
rect 79468 287036 79474 287088
rect 96522 287076 96528 287088
rect 96481 287048 96528 287076
rect 96522 287036 96528 287048
rect 96580 287076 96586 287088
rect 162854 287076 162860 287088
rect 96580 287048 162860 287076
rect 96580 287036 96614 287048
rect 162854 287036 162860 287048
rect 162912 287036 162918 287088
rect 166902 287036 166908 287088
rect 166960 287076 166966 287088
rect 191742 287076 191748 287088
rect 166960 287048 191748 287076
rect 166960 287036 166966 287048
rect 191742 287036 191748 287048
rect 191800 287036 191806 287088
rect 255498 287036 255504 287088
rect 255556 287076 255562 287088
rect 258350 287076 258356 287088
rect 255556 287048 258356 287076
rect 255556 287036 255562 287048
rect 258350 287036 258356 287048
rect 258408 287076 258414 287088
rect 259454 287076 259460 287088
rect 258408 287048 259460 287076
rect 258408 287036 258414 287048
rect 259454 287036 259460 287048
rect 259512 287036 259518 287088
rect 92382 286968 92388 287020
rect 92440 287008 92446 287020
rect 93118 287008 93124 287020
rect 92440 286980 93124 287008
rect 92440 286968 92446 286980
rect 93118 286968 93124 286980
rect 93176 286968 93182 287020
rect 94682 286968 94688 287020
rect 94740 287008 94746 287020
rect 96586 287008 96614 287036
rect 94740 286980 96614 287008
rect 94740 286968 94746 286980
rect 255314 286968 255320 287020
rect 255372 287008 255378 287020
rect 255372 286980 255544 287008
rect 255372 286968 255378 286980
rect 255516 286952 255544 286980
rect 255590 286968 255596 287020
rect 255648 287008 255654 287020
rect 261018 287008 261024 287020
rect 255648 286980 261024 287008
rect 255648 286968 255654 286980
rect 261018 286968 261024 286980
rect 261076 286968 261082 287020
rect 255498 286900 255504 286952
rect 255556 286900 255562 286952
rect 176102 286356 176108 286408
rect 176160 286396 176166 286408
rect 188706 286396 188712 286408
rect 176160 286368 188712 286396
rect 176160 286356 176166 286368
rect 188706 286356 188712 286368
rect 188764 286356 188770 286408
rect 71774 286288 71780 286340
rect 71832 286328 71838 286340
rect 77018 286328 77024 286340
rect 71832 286300 77024 286328
rect 71832 286288 71838 286300
rect 77018 286288 77024 286300
rect 77076 286328 77082 286340
rect 188430 286328 188436 286340
rect 77076 286300 188436 286328
rect 77076 286288 77082 286300
rect 188430 286288 188436 286300
rect 188488 286288 188494 286340
rect 255406 286288 255412 286340
rect 255464 286328 255470 286340
rect 267734 286328 267740 286340
rect 255464 286300 267740 286328
rect 255464 286288 255470 286300
rect 267734 286288 267740 286300
rect 267792 286288 267798 286340
rect 64506 285676 64512 285728
rect 64564 285716 64570 285728
rect 80790 285716 80796 285728
rect 64564 285688 80796 285716
rect 64564 285676 64570 285688
rect 80790 285676 80796 285688
rect 80848 285676 80854 285728
rect 69474 284928 69480 284980
rect 69532 284968 69538 284980
rect 69658 284968 69664 284980
rect 69532 284940 69664 284968
rect 69532 284928 69538 284940
rect 69658 284928 69664 284940
rect 69716 284928 69722 284980
rect 82906 284928 82912 284980
rect 82964 284968 82970 284980
rect 83550 284968 83556 284980
rect 82964 284940 83556 284968
rect 82964 284928 82970 284940
rect 83550 284928 83556 284940
rect 83608 284928 83614 284980
rect 63126 284384 63132 284436
rect 63184 284424 63190 284436
rect 72418 284424 72424 284436
rect 63184 284396 72424 284424
rect 63184 284384 63190 284396
rect 72418 284384 72424 284396
rect 72476 284384 72482 284436
rect 86862 284384 86868 284436
rect 86920 284424 86926 284436
rect 98454 284424 98460 284436
rect 86920 284396 98460 284424
rect 86920 284384 86926 284396
rect 98454 284384 98460 284396
rect 98512 284384 98518 284436
rect 158714 284384 158720 284436
rect 158772 284424 158778 284436
rect 191558 284424 191564 284436
rect 158772 284396 191564 284424
rect 158772 284384 158778 284396
rect 191558 284384 191564 284396
rect 191616 284384 191622 284436
rect 255498 284384 255504 284436
rect 255556 284424 255562 284436
rect 266354 284424 266360 284436
rect 255556 284396 266360 284424
rect 255556 284384 255562 284396
rect 266354 284384 266360 284396
rect 266412 284384 266418 284436
rect 68554 284316 68560 284368
rect 68612 284356 68618 284368
rect 164970 284356 164976 284368
rect 68612 284328 164976 284356
rect 68612 284316 68618 284328
rect 164970 284316 164976 284328
rect 165028 284316 165034 284368
rect 255406 284316 255412 284368
rect 255464 284356 255470 284368
rect 269298 284356 269304 284368
rect 255464 284328 269304 284356
rect 255464 284316 255470 284328
rect 269298 284316 269304 284328
rect 269356 284316 269362 284368
rect 89944 283704 89950 283756
rect 90002 283744 90008 283756
rect 91002 283744 91008 283756
rect 90002 283716 91008 283744
rect 90002 283704 90008 283716
rect 91002 283704 91008 283716
rect 91060 283704 91066 283756
rect 53466 283568 53472 283620
rect 53524 283608 53530 283620
rect 57698 283608 57704 283620
rect 53524 283580 57704 283608
rect 53524 283568 53530 283580
rect 57698 283568 57704 283580
rect 57756 283608 57762 283620
rect 66806 283608 66812 283620
rect 57756 283580 66812 283608
rect 57756 283568 57762 283580
rect 66806 283568 66812 283580
rect 66864 283568 66870 283620
rect 68830 283568 68836 283620
rect 68888 283608 68894 283620
rect 169018 283608 169024 283620
rect 68888 283580 169024 283608
rect 68888 283568 68894 283580
rect 169018 283568 169024 283580
rect 169076 283568 169082 283620
rect 66162 283024 66168 283076
rect 66220 283064 66226 283076
rect 66220 283036 70394 283064
rect 66220 283024 66226 283036
rect 69658 282956 69664 283008
rect 69716 282956 69722 283008
rect 70366 282996 70394 283036
rect 81434 282996 81440 283008
rect 70366 282968 81440 282996
rect 81434 282956 81440 282968
rect 81492 282956 81498 283008
rect 89622 282956 89628 283008
rect 89680 282996 89686 283008
rect 89680 282956 89714 282996
rect 63310 282820 63316 282872
rect 63368 282860 63374 282872
rect 63368 282832 64874 282860
rect 63368 282820 63374 282832
rect 64846 282792 64874 282832
rect 69676 282792 69704 282956
rect 89686 282928 89714 282956
rect 89686 282900 128400 282928
rect 128372 282860 128400 282900
rect 178034 282888 178040 282940
rect 178092 282928 178098 282940
rect 179230 282928 179236 282940
rect 178092 282900 179236 282928
rect 178092 282888 178098 282900
rect 179230 282888 179236 282900
rect 179288 282928 179294 282940
rect 191006 282928 191012 282940
rect 179288 282900 191012 282928
rect 179288 282888 179294 282900
rect 191006 282888 191012 282900
rect 191064 282888 191070 282940
rect 255406 282888 255412 282940
rect 255464 282928 255470 282940
rect 270678 282928 270684 282940
rect 255464 282900 270684 282928
rect 255464 282888 255470 282900
rect 270678 282888 270684 282900
rect 270736 282888 270742 282940
rect 192386 282860 192392 282872
rect 128372 282832 192392 282860
rect 192386 282820 192392 282832
rect 192444 282820 192450 282872
rect 255498 282820 255504 282872
rect 255556 282860 255562 282872
rect 262490 282860 262496 282872
rect 255556 282832 262496 282860
rect 255556 282820 255562 282832
rect 262490 282820 262496 282832
rect 262548 282820 262554 282872
rect 64846 282764 69704 282792
rect 69032 282736 69060 282764
rect 69014 282684 69020 282736
rect 69072 282684 69078 282736
rect 255406 282684 255412 282736
rect 255464 282724 255470 282736
rect 258258 282724 258264 282736
rect 255464 282696 258264 282724
rect 255464 282684 255470 282696
rect 258258 282684 258264 282696
rect 258316 282684 258322 282736
rect 97994 282208 98000 282260
rect 98052 282248 98058 282260
rect 98730 282248 98736 282260
rect 98052 282220 98736 282248
rect 98052 282208 98058 282220
rect 98730 282208 98736 282220
rect 98788 282208 98794 282260
rect 100754 281528 100760 281580
rect 100812 281568 100818 281580
rect 149698 281568 149704 281580
rect 100812 281540 149704 281568
rect 100812 281528 100818 281540
rect 149698 281528 149704 281540
rect 149756 281528 149762 281580
rect 107010 281460 107016 281512
rect 107068 281500 107074 281512
rect 158714 281500 158720 281512
rect 107068 281472 158720 281500
rect 107068 281460 107074 281472
rect 158714 281460 158720 281472
rect 158772 281460 158778 281512
rect 162854 281460 162860 281512
rect 162912 281500 162918 281512
rect 164142 281500 164148 281512
rect 162912 281472 164148 281500
rect 162912 281460 162918 281472
rect 164142 281460 164148 281472
rect 164200 281460 164206 281512
rect 255406 281460 255412 281512
rect 255464 281500 255470 281512
rect 265066 281500 265072 281512
rect 255464 281472 265072 281500
rect 255464 281460 255470 281472
rect 265066 281460 265072 281472
rect 265124 281460 265130 281512
rect 100754 281392 100760 281444
rect 100812 281432 100818 281444
rect 135898 281432 135904 281444
rect 100812 281404 135904 281432
rect 100812 281392 100818 281404
rect 135898 281392 135904 281404
rect 135956 281392 135962 281444
rect 164142 280780 164148 280832
rect 164200 280820 164206 280832
rect 191742 280820 191748 280832
rect 164200 280792 191748 280820
rect 164200 280780 164206 280792
rect 191742 280780 191748 280792
rect 191800 280780 191806 280832
rect 10318 280168 10324 280220
rect 10376 280208 10382 280220
rect 67266 280208 67272 280220
rect 10376 280180 67272 280208
rect 10376 280168 10382 280180
rect 67266 280168 67272 280180
rect 67324 280208 67330 280220
rect 68830 280208 68836 280220
rect 67324 280180 68836 280208
rect 67324 280168 67330 280180
rect 68830 280168 68836 280180
rect 68888 280168 68894 280220
rect 255406 280168 255412 280220
rect 255464 280208 255470 280220
rect 262214 280208 262220 280220
rect 255464 280180 262220 280208
rect 255464 280168 255470 280180
rect 262214 280168 262220 280180
rect 262272 280168 262278 280220
rect 126974 280100 126980 280152
rect 127032 280140 127038 280152
rect 127434 280140 127440 280152
rect 127032 280112 127440 280140
rect 127032 280100 127038 280112
rect 127434 280100 127440 280112
rect 127492 280140 127498 280152
rect 185578 280140 185584 280152
rect 127492 280112 185584 280140
rect 127492 280100 127498 280112
rect 185578 280100 185584 280112
rect 185636 280100 185642 280152
rect 100754 280032 100760 280084
rect 100812 280072 100818 280084
rect 142890 280072 142896 280084
rect 100812 280044 142896 280072
rect 100812 280032 100818 280044
rect 142890 280032 142896 280044
rect 142948 280032 142954 280084
rect 7558 279420 7564 279472
rect 7616 279460 7622 279472
rect 34330 279460 34336 279472
rect 7616 279432 34336 279460
rect 7616 279420 7622 279432
rect 34330 279420 34336 279432
rect 34388 279460 34394 279472
rect 65886 279460 65892 279472
rect 34388 279432 65892 279460
rect 34388 279420 34394 279432
rect 65886 279420 65892 279432
rect 65944 279460 65950 279472
rect 66530 279460 66536 279472
rect 65944 279432 66536 279460
rect 65944 279420 65950 279432
rect 66530 279420 66536 279432
rect 66588 279420 66594 279472
rect 102226 279420 102232 279472
rect 102284 279460 102290 279472
rect 127434 279460 127440 279472
rect 102284 279432 127440 279460
rect 102284 279420 102290 279432
rect 127434 279420 127440 279432
rect 127492 279420 127498 279472
rect 255314 278740 255320 278792
rect 255372 278780 255378 278792
rect 266538 278780 266544 278792
rect 255372 278752 266544 278780
rect 255372 278740 255378 278752
rect 266538 278740 266544 278752
rect 266596 278740 266602 278792
rect 47946 278672 47952 278724
rect 48004 278712 48010 278724
rect 48130 278712 48136 278724
rect 48004 278684 48136 278712
rect 48004 278672 48010 278684
rect 48130 278672 48136 278684
rect 48188 278672 48194 278724
rect 99374 278672 99380 278724
rect 99432 278712 99438 278724
rect 102042 278712 102048 278724
rect 99432 278684 102048 278712
rect 99432 278672 99438 278684
rect 102042 278672 102048 278684
rect 102100 278712 102106 278724
rect 122098 278712 122104 278724
rect 102100 278684 122104 278712
rect 102100 278672 102106 278684
rect 122098 278672 122104 278684
rect 122156 278672 122162 278724
rect 255498 278672 255504 278724
rect 255556 278712 255562 278724
rect 263870 278712 263876 278724
rect 255556 278684 263876 278712
rect 255556 278672 255562 278684
rect 263870 278672 263876 278684
rect 263928 278672 263934 278724
rect 152642 278060 152648 278112
rect 152700 278100 152706 278112
rect 188522 278100 188528 278112
rect 152700 278072 188528 278100
rect 152700 278060 152706 278072
rect 188522 278060 188528 278072
rect 188580 278060 188586 278112
rect 47946 277992 47952 278044
rect 48004 278032 48010 278044
rect 66806 278032 66812 278044
rect 48004 278004 66812 278032
rect 48004 277992 48010 278004
rect 66806 277992 66812 278004
rect 66864 277992 66870 278044
rect 98454 277992 98460 278044
rect 98512 278032 98518 278044
rect 177850 278032 177856 278044
rect 98512 278004 177856 278032
rect 98512 277992 98518 278004
rect 177850 277992 177856 278004
rect 177908 277992 177914 278044
rect 255406 277448 255412 277500
rect 255464 277488 255470 277500
rect 259730 277488 259736 277500
rect 255464 277460 259736 277488
rect 255464 277448 255470 277460
rect 259730 277448 259736 277460
rect 259788 277448 259794 277500
rect 188614 277380 188620 277432
rect 188672 277420 188678 277432
rect 191650 277420 191656 277432
rect 188672 277392 191656 277420
rect 188672 277380 188678 277392
rect 191650 277380 191656 277392
rect 191708 277380 191714 277432
rect 55122 277312 55128 277364
rect 55180 277352 55186 277364
rect 66898 277352 66904 277364
rect 55180 277324 66904 277352
rect 55180 277312 55186 277324
rect 66898 277312 66904 277324
rect 66956 277312 66962 277364
rect 177942 277312 177948 277364
rect 178000 277352 178006 277364
rect 187142 277352 187148 277364
rect 178000 277324 187148 277352
rect 178000 277312 178006 277324
rect 187142 277312 187148 277324
rect 187200 277312 187206 277364
rect 255406 277108 255412 277160
rect 255464 277148 255470 277160
rect 259546 277148 259552 277160
rect 255464 277120 259552 277148
rect 255464 277108 255470 277120
rect 259546 277108 259552 277120
rect 259604 277108 259610 277160
rect 100754 276632 100760 276684
rect 100812 276672 100818 276684
rect 118786 276672 118792 276684
rect 100812 276644 118792 276672
rect 100812 276632 100818 276644
rect 118786 276632 118792 276644
rect 118844 276632 118850 276684
rect 169202 276632 169208 276684
rect 169260 276672 169266 276684
rect 190454 276672 190460 276684
rect 169260 276644 190460 276672
rect 169260 276632 169266 276644
rect 190454 276632 190460 276644
rect 190512 276632 190518 276684
rect 61930 276156 61936 276208
rect 61988 276196 61994 276208
rect 66806 276196 66812 276208
rect 61988 276168 66812 276196
rect 61988 276156 61994 276168
rect 66806 276156 66812 276168
rect 66864 276156 66870 276208
rect 255498 276020 255504 276072
rect 255556 276060 255562 276072
rect 273438 276060 273444 276072
rect 255556 276032 273444 276060
rect 255556 276020 255562 276032
rect 273438 276020 273444 276032
rect 273496 276020 273502 276072
rect 64690 275952 64696 276004
rect 64748 275992 64754 276004
rect 66622 275992 66628 276004
rect 64748 275964 66628 275992
rect 64748 275952 64754 275964
rect 66622 275952 66628 275964
rect 66680 275952 66686 276004
rect 255406 275952 255412 276004
rect 255464 275992 255470 276004
rect 267826 275992 267832 276004
rect 255464 275964 267832 275992
rect 255464 275952 255470 275964
rect 267826 275952 267832 275964
rect 267884 275952 267890 276004
rect 100846 275340 100852 275392
rect 100904 275380 100910 275392
rect 148410 275380 148416 275392
rect 100904 275352 148416 275380
rect 100904 275340 100910 275352
rect 148410 275340 148416 275352
rect 148468 275340 148474 275392
rect 54938 275272 54944 275324
rect 54996 275312 55002 275324
rect 61930 275312 61936 275324
rect 54996 275284 61936 275312
rect 54996 275272 55002 275284
rect 61930 275272 61936 275284
rect 61988 275272 61994 275324
rect 100110 275272 100116 275324
rect 100168 275312 100174 275324
rect 181622 275312 181628 275324
rect 100168 275284 181628 275312
rect 100168 275272 100174 275284
rect 181622 275272 181628 275284
rect 181680 275272 181686 275324
rect 255406 274660 255412 274712
rect 255464 274700 255470 274712
rect 281626 274700 281632 274712
rect 255464 274672 281632 274700
rect 255464 274660 255470 274672
rect 281626 274660 281632 274672
rect 281684 274660 281690 274712
rect 100754 274592 100760 274644
rect 100812 274632 100818 274644
rect 146938 274632 146944 274644
rect 100812 274604 146944 274632
rect 100812 274592 100818 274604
rect 146938 274592 146944 274604
rect 146996 274592 147002 274644
rect 255498 274592 255504 274644
rect 255556 274632 255562 274644
rect 269206 274632 269212 274644
rect 255556 274604 269212 274632
rect 255556 274592 255562 274604
rect 269206 274592 269212 274604
rect 269264 274632 269270 274644
rect 274634 274632 274640 274644
rect 269264 274604 274640 274632
rect 269264 274592 269270 274604
rect 274634 274592 274640 274604
rect 274692 274592 274698 274644
rect 255314 274524 255320 274576
rect 255372 274564 255378 274576
rect 258074 274564 258080 274576
rect 255372 274536 258080 274564
rect 255372 274524 255378 274536
rect 258074 274524 258080 274536
rect 258132 274524 258138 274576
rect 134610 273912 134616 273964
rect 134668 273952 134674 273964
rect 156690 273952 156696 273964
rect 134668 273924 156696 273952
rect 134668 273912 134674 273924
rect 156690 273912 156696 273924
rect 156748 273912 156754 273964
rect 180058 273232 180064 273284
rect 180116 273272 180122 273284
rect 191650 273272 191656 273284
rect 180116 273244 191656 273272
rect 180116 273232 180122 273244
rect 191650 273232 191656 273244
rect 191708 273232 191714 273284
rect 100754 273164 100760 273216
rect 100812 273204 100818 273216
rect 105722 273204 105728 273216
rect 100812 273176 105728 273204
rect 100812 273164 100818 273176
rect 105722 273164 105728 273176
rect 105780 273164 105786 273216
rect 255406 273164 255412 273216
rect 255464 273204 255470 273216
rect 263686 273204 263692 273216
rect 255464 273176 263692 273204
rect 255464 273164 255470 273176
rect 263686 273164 263692 273176
rect 263744 273164 263750 273216
rect 106182 272552 106188 272604
rect 106240 272592 106246 272604
rect 142982 272592 142988 272604
rect 106240 272564 142988 272592
rect 106240 272552 106246 272564
rect 142982 272552 142988 272564
rect 143040 272552 143046 272604
rect 146938 272552 146944 272604
rect 146996 272592 147002 272604
rect 180150 272592 180156 272604
rect 146996 272564 180156 272592
rect 146996 272552 147002 272564
rect 180150 272552 180156 272564
rect 180208 272552 180214 272604
rect 46658 272484 46664 272536
rect 46716 272524 46722 272536
rect 52362 272524 52368 272536
rect 46716 272496 52368 272524
rect 46716 272484 46722 272496
rect 52362 272484 52368 272496
rect 52420 272524 52426 272536
rect 66806 272524 66812 272536
rect 52420 272496 66812 272524
rect 52420 272484 52426 272496
rect 66806 272484 66812 272496
rect 66864 272484 66870 272536
rect 124122 272484 124128 272536
rect 124180 272524 124186 272536
rect 175918 272524 175924 272536
rect 124180 272496 175924 272524
rect 124180 272484 124186 272496
rect 175918 272484 175924 272496
rect 175976 272484 175982 272536
rect 101122 272008 101128 272060
rect 101180 272048 101186 272060
rect 101858 272048 101864 272060
rect 101180 272020 101864 272048
rect 101180 272008 101186 272020
rect 101858 272008 101864 272020
rect 101916 272048 101922 272060
rect 104894 272048 104900 272060
rect 101916 272020 104900 272048
rect 101916 272008 101922 272020
rect 104894 272008 104900 272020
rect 104952 272048 104958 272060
rect 106182 272048 106188 272060
rect 104952 272020 106188 272048
rect 104952 272008 104958 272020
rect 106182 272008 106188 272020
rect 106240 272008 106246 272060
rect 187142 271940 187148 271992
rect 187200 271980 187206 271992
rect 191650 271980 191656 271992
rect 187200 271952 191656 271980
rect 187200 271940 187206 271952
rect 191650 271940 191656 271952
rect 191708 271940 191714 271992
rect 181530 271872 181536 271924
rect 181588 271912 181594 271924
rect 191558 271912 191564 271924
rect 181588 271884 191564 271912
rect 181588 271872 181594 271884
rect 191558 271872 191564 271884
rect 191616 271872 191622 271924
rect 565078 271872 565084 271924
rect 565136 271912 565142 271924
rect 580166 271912 580172 271924
rect 565136 271884 580172 271912
rect 565136 271872 565142 271884
rect 580166 271872 580172 271884
rect 580224 271872 580230 271924
rect 99282 271532 99288 271584
rect 99340 271572 99346 271584
rect 105538 271572 105544 271584
rect 99340 271544 105544 271572
rect 99340 271532 99346 271544
rect 105538 271532 105544 271544
rect 105596 271532 105602 271584
rect 148410 271192 148416 271244
rect 148468 271232 148474 271244
rect 188338 271232 188344 271244
rect 148468 271204 188344 271232
rect 148468 271192 148474 271204
rect 188338 271192 188344 271204
rect 188396 271192 188402 271244
rect 53742 271124 53748 271176
rect 53800 271164 53806 271176
rect 66254 271164 66260 271176
rect 53800 271136 66260 271164
rect 53800 271124 53806 271136
rect 66254 271124 66260 271136
rect 66312 271124 66318 271176
rect 141510 271124 141516 271176
rect 141568 271164 141574 271176
rect 187050 271164 187056 271176
rect 141568 271136 187056 271164
rect 141568 271124 141574 271136
rect 187050 271124 187056 271136
rect 187108 271124 187114 271176
rect 255958 271124 255964 271176
rect 256016 271164 256022 271176
rect 266446 271164 266452 271176
rect 256016 271136 266452 271164
rect 256016 271124 256022 271136
rect 266446 271124 266452 271136
rect 266504 271124 266510 271176
rect 100294 270444 100300 270496
rect 100352 270484 100358 270496
rect 106182 270484 106188 270496
rect 100352 270456 106188 270484
rect 100352 270444 100358 270456
rect 106182 270444 106188 270456
rect 106240 270444 106246 270496
rect 56318 269764 56324 269816
rect 56376 269804 56382 269816
rect 66254 269804 66260 269816
rect 56376 269776 66260 269804
rect 56376 269764 56382 269776
rect 66254 269764 66260 269776
rect 66312 269764 66318 269816
rect 126514 269764 126520 269816
rect 126572 269804 126578 269816
rect 159450 269804 159456 269816
rect 126572 269776 159456 269804
rect 126572 269764 126578 269776
rect 159450 269764 159456 269776
rect 159508 269764 159514 269816
rect 255498 269152 255504 269204
rect 255556 269192 255562 269204
rect 261018 269192 261024 269204
rect 255556 269164 261024 269192
rect 255556 269152 255562 269164
rect 261018 269152 261024 269164
rect 261076 269152 261082 269204
rect 166258 269084 166264 269136
rect 166316 269124 166322 269136
rect 191650 269124 191656 269136
rect 166316 269096 191656 269124
rect 166316 269084 166322 269096
rect 191650 269084 191656 269096
rect 191708 269084 191714 269136
rect 255406 269084 255412 269136
rect 255464 269124 255470 269136
rect 268010 269124 268016 269136
rect 255464 269096 268016 269124
rect 255464 269084 255470 269096
rect 268010 269084 268016 269096
rect 268068 269084 268074 269136
rect 115934 268608 115940 268660
rect 115992 268648 115998 268660
rect 116670 268648 116676 268660
rect 115992 268620 116676 268648
rect 115992 268608 115998 268620
rect 116670 268608 116676 268620
rect 116728 268608 116734 268660
rect 101214 268404 101220 268456
rect 101272 268444 101278 268456
rect 113818 268444 113824 268456
rect 101272 268416 113824 268444
rect 101272 268404 101278 268416
rect 113818 268404 113824 268416
rect 113876 268404 113882 268456
rect 44082 268336 44088 268388
rect 44140 268376 44146 268388
rect 53558 268376 53564 268388
rect 44140 268348 53564 268376
rect 44140 268336 44146 268348
rect 53558 268336 53564 268348
rect 53616 268336 53622 268388
rect 100754 268336 100760 268388
rect 100812 268376 100818 268388
rect 115934 268376 115940 268388
rect 100812 268348 115940 268376
rect 100812 268336 100818 268348
rect 115934 268336 115940 268348
rect 115992 268336 115998 268388
rect 145558 268336 145564 268388
rect 145616 268376 145622 268388
rect 166350 268376 166356 268388
rect 145616 268348 166356 268376
rect 145616 268336 145622 268348
rect 166350 268336 166356 268348
rect 166408 268336 166414 268388
rect 255406 267792 255412 267844
rect 255464 267832 255470 267844
rect 267826 267832 267832 267844
rect 255464 267804 267832 267832
rect 255464 267792 255470 267804
rect 267826 267792 267832 267804
rect 267884 267792 267890 267844
rect 53558 267724 53564 267776
rect 53616 267764 53622 267776
rect 66806 267764 66812 267776
rect 53616 267736 66812 267764
rect 53616 267724 53622 267736
rect 66806 267724 66812 267736
rect 66864 267724 66870 267776
rect 164878 267724 164884 267776
rect 164936 267764 164942 267776
rect 191650 267764 191656 267776
rect 164936 267736 191656 267764
rect 164936 267724 164942 267736
rect 191650 267724 191656 267736
rect 191708 267724 191714 267776
rect 255314 267724 255320 267776
rect 255372 267764 255378 267776
rect 273530 267764 273536 267776
rect 255372 267736 273536 267764
rect 255372 267724 255378 267736
rect 273530 267724 273536 267736
rect 273588 267724 273594 267776
rect 3510 267656 3516 267708
rect 3568 267696 3574 267708
rect 36538 267696 36544 267708
rect 3568 267668 36544 267696
rect 3568 267656 3574 267668
rect 36538 267656 36544 267668
rect 36596 267656 36602 267708
rect 100754 267656 100760 267708
rect 100812 267696 100818 267708
rect 122926 267696 122932 267708
rect 100812 267668 122932 267696
rect 100812 267656 100818 267668
rect 122926 267656 122932 267668
rect 122984 267656 122990 267708
rect 255498 267656 255504 267708
rect 255556 267696 255562 267708
rect 277302 267696 277308 267708
rect 255556 267668 277308 267696
rect 255556 267656 255562 267668
rect 277302 267656 277308 267668
rect 277360 267656 277366 267708
rect 142890 266976 142896 267028
rect 142948 267016 142954 267028
rect 173250 267016 173256 267028
rect 142948 266988 173256 267016
rect 142948 266976 142954 266988
rect 173250 266976 173256 266988
rect 173308 266976 173314 267028
rect 173158 266432 173164 266484
rect 173216 266472 173222 266484
rect 191006 266472 191012 266484
rect 173216 266444 191012 266472
rect 173216 266432 173222 266444
rect 191006 266432 191012 266444
rect 191064 266432 191070 266484
rect 63310 266364 63316 266416
rect 63368 266404 63374 266416
rect 66806 266404 66812 266416
rect 63368 266376 66812 266404
rect 63368 266364 63374 266376
rect 66806 266364 66812 266376
rect 66864 266364 66870 266416
rect 122926 266364 122932 266416
rect 122984 266404 122990 266416
rect 131758 266404 131764 266416
rect 122984 266376 131764 266404
rect 122984 266364 122990 266376
rect 131758 266364 131764 266376
rect 131816 266364 131822 266416
rect 157978 266364 157984 266416
rect 158036 266404 158042 266416
rect 191282 266404 191288 266416
rect 158036 266376 191288 266404
rect 158036 266364 158042 266376
rect 191282 266364 191288 266376
rect 191340 266364 191346 266416
rect 255406 266364 255412 266416
rect 255464 266404 255470 266416
rect 265158 266404 265164 266416
rect 255464 266376 265164 266404
rect 255464 266364 255470 266376
rect 265158 266364 265164 266376
rect 265216 266364 265222 266416
rect 277302 266364 277308 266416
rect 277360 266404 277366 266416
rect 277486 266404 277492 266416
rect 277360 266376 277492 266404
rect 277360 266364 277366 266376
rect 277486 266364 277492 266376
rect 277544 266364 277550 266416
rect 100846 266296 100852 266348
rect 100904 266336 100910 266348
rect 142154 266336 142160 266348
rect 100904 266308 142160 266336
rect 100904 266296 100910 266308
rect 142154 266296 142160 266308
rect 142212 266336 142218 266348
rect 143442 266336 143448 266348
rect 142212 266308 143448 266336
rect 142212 266296 142218 266308
rect 143442 266296 143448 266308
rect 143500 266296 143506 266348
rect 254026 266296 254032 266348
rect 254084 266336 254090 266348
rect 263778 266336 263784 266348
rect 254084 266308 263784 266336
rect 254084 266296 254090 266308
rect 263778 266296 263784 266308
rect 263836 266296 263842 266348
rect 143442 265684 143448 265736
rect 143500 265724 143506 265736
rect 152550 265724 152556 265736
rect 143500 265696 152556 265724
rect 143500 265684 143506 265696
rect 152550 265684 152556 265696
rect 152608 265684 152614 265736
rect 41230 265616 41236 265668
rect 41288 265656 41294 265668
rect 50522 265656 50528 265668
rect 41288 265628 50528 265656
rect 41288 265616 41294 265628
rect 50522 265616 50528 265628
rect 50580 265616 50586 265668
rect 105538 265616 105544 265668
rect 105596 265656 105602 265668
rect 115290 265656 115296 265668
rect 105596 265628 115296 265656
rect 105596 265616 105602 265628
rect 115290 265616 115296 265628
rect 115348 265616 115354 265668
rect 140038 265616 140044 265668
rect 140096 265656 140102 265668
rect 182910 265656 182916 265668
rect 140096 265628 182916 265656
rect 140096 265616 140102 265628
rect 182910 265616 182916 265628
rect 182968 265616 182974 265668
rect 61838 265140 61844 265192
rect 61896 265180 61902 265192
rect 65702 265180 65708 265192
rect 61896 265152 65708 265180
rect 61896 265140 61902 265152
rect 65702 265140 65708 265152
rect 65760 265140 65766 265192
rect 255314 265004 255320 265056
rect 255372 265044 255378 265056
rect 263686 265044 263692 265056
rect 255372 265016 263692 265044
rect 255372 265004 255378 265016
rect 263686 265004 263692 265016
rect 263744 265004 263750 265056
rect 167638 264936 167644 264988
rect 167696 264976 167702 264988
rect 191558 264976 191564 264988
rect 167696 264948 191564 264976
rect 167696 264936 167702 264948
rect 191558 264936 191564 264948
rect 191616 264936 191622 264988
rect 100754 264868 100760 264920
rect 100812 264908 100818 264920
rect 139394 264908 139400 264920
rect 100812 264880 139400 264908
rect 100812 264868 100818 264880
rect 139394 264868 139400 264880
rect 139452 264908 139458 264920
rect 144270 264908 144276 264920
rect 139452 264880 144276 264908
rect 139452 264868 139458 264880
rect 144270 264868 144276 264880
rect 144328 264868 144334 264920
rect 98270 264188 98276 264240
rect 98328 264228 98334 264240
rect 115290 264228 115296 264240
rect 98328 264200 115296 264228
rect 98328 264188 98334 264200
rect 115290 264188 115296 264200
rect 115348 264188 115354 264240
rect 147122 264188 147128 264240
rect 147180 264228 147186 264240
rect 176102 264228 176108 264240
rect 147180 264200 176108 264228
rect 147180 264188 147186 264200
rect 176102 264188 176108 264200
rect 176160 264188 176166 264240
rect 255314 263644 255320 263696
rect 255372 263684 255378 263696
rect 271966 263684 271972 263696
rect 255372 263656 271972 263684
rect 255372 263644 255378 263656
rect 271966 263644 271972 263656
rect 272024 263684 272030 263696
rect 273346 263684 273352 263696
rect 272024 263656 273352 263684
rect 272024 263644 272030 263656
rect 273346 263644 273352 263656
rect 273404 263644 273410 263696
rect 3418 263576 3424 263628
rect 3476 263616 3482 263628
rect 3476 263588 52776 263616
rect 3476 263576 3482 263588
rect 52748 263548 52776 263588
rect 99282 263576 99288 263628
rect 99340 263616 99346 263628
rect 101214 263616 101220 263628
rect 99340 263588 101220 263616
rect 99340 263576 99346 263588
rect 101214 263576 101220 263588
rect 101272 263576 101278 263628
rect 255498 263576 255504 263628
rect 255556 263616 255562 263628
rect 278866 263616 278872 263628
rect 255556 263588 278872 263616
rect 255556 263576 255562 263588
rect 278866 263576 278872 263588
rect 278924 263616 278930 263628
rect 282178 263616 282184 263628
rect 278924 263588 282184 263616
rect 278924 263576 278930 263588
rect 282178 263576 282184 263588
rect 282236 263576 282242 263628
rect 53098 263548 53104 263560
rect 52748 263520 53104 263548
rect 53098 263508 53104 263520
rect 53156 263548 53162 263560
rect 66898 263548 66904 263560
rect 53156 263520 66904 263548
rect 53156 263508 53162 263520
rect 66898 263508 66904 263520
rect 66956 263508 66962 263560
rect 101674 263508 101680 263560
rect 101732 263548 101738 263560
rect 103422 263548 103428 263560
rect 101732 263520 103428 263548
rect 101732 263508 101738 263520
rect 103422 263508 103428 263520
rect 103480 263548 103486 263560
rect 117958 263548 117964 263560
rect 103480 263520 117964 263548
rect 103480 263508 103486 263520
rect 117958 263508 117964 263520
rect 118016 263508 118022 263560
rect 255406 263032 255412 263084
rect 255464 263072 255470 263084
rect 258350 263072 258356 263084
rect 255464 263044 258356 263072
rect 255464 263032 255470 263044
rect 258350 263032 258356 263044
rect 258408 263032 258414 263084
rect 7558 262828 7564 262880
rect 7616 262868 7622 262880
rect 32950 262868 32956 262880
rect 7616 262840 32956 262868
rect 7616 262828 7622 262840
rect 32950 262828 32956 262840
rect 33008 262868 33014 262880
rect 65886 262868 65892 262880
rect 33008 262840 65892 262868
rect 33008 262828 33014 262840
rect 65886 262828 65892 262840
rect 65944 262868 65950 262880
rect 66530 262868 66536 262880
rect 65944 262840 66536 262868
rect 65944 262828 65950 262840
rect 66530 262828 66536 262840
rect 66588 262828 66594 262880
rect 141418 262828 141424 262880
rect 141476 262868 141482 262880
rect 153838 262868 153844 262880
rect 141476 262840 153844 262868
rect 141476 262828 141482 262840
rect 153838 262828 153844 262840
rect 153896 262828 153902 262880
rect 121362 262624 121368 262676
rect 121420 262664 121426 262676
rect 121546 262664 121552 262676
rect 121420 262636 121552 262664
rect 121420 262624 121426 262636
rect 121546 262624 121552 262636
rect 121604 262624 121610 262676
rect 177298 262284 177304 262336
rect 177356 262324 177362 262336
rect 191650 262324 191656 262336
rect 177356 262296 191656 262324
rect 177356 262284 177362 262296
rect 191650 262284 191656 262296
rect 191708 262284 191714 262336
rect 100754 262216 100760 262268
rect 100812 262256 100818 262268
rect 121362 262256 121368 262268
rect 100812 262228 121368 262256
rect 100812 262216 100818 262228
rect 121362 262216 121368 262228
rect 121420 262216 121426 262268
rect 126330 262216 126336 262268
rect 126388 262256 126394 262268
rect 191190 262256 191196 262268
rect 126388 262228 191196 262256
rect 126388 262216 126394 262228
rect 191190 262216 191196 262228
rect 191248 262216 191254 262268
rect 255406 262216 255412 262268
rect 255464 262256 255470 262268
rect 265066 262256 265072 262268
rect 255464 262228 265072 262256
rect 255464 262216 255470 262228
rect 265066 262216 265072 262228
rect 265124 262216 265130 262268
rect 255498 262148 255504 262200
rect 255556 262188 255562 262200
rect 285674 262188 285680 262200
rect 255556 262160 285680 262188
rect 255556 262148 255562 262160
rect 285674 262148 285680 262160
rect 285732 262148 285738 262200
rect 255314 262080 255320 262132
rect 255372 262120 255378 262132
rect 263594 262120 263600 262132
rect 255372 262092 263600 262120
rect 255372 262080 255378 262092
rect 263594 262080 263600 262092
rect 263652 262080 263658 262132
rect 103422 261536 103428 261588
rect 103480 261576 103486 261588
rect 109034 261576 109040 261588
rect 103480 261548 109040 261576
rect 103480 261536 103486 261548
rect 109034 261536 109040 261548
rect 109092 261536 109098 261588
rect 56410 261468 56416 261520
rect 56468 261508 56474 261520
rect 66254 261508 66260 261520
rect 56468 261480 66260 261508
rect 56468 261468 56474 261480
rect 66254 261468 66260 261480
rect 66312 261468 66318 261520
rect 108206 261468 108212 261520
rect 108264 261508 108270 261520
rect 143626 261508 143632 261520
rect 108264 261480 143632 261508
rect 108264 261468 108270 261480
rect 143626 261468 143632 261480
rect 143684 261508 143690 261520
rect 180242 261508 180248 261520
rect 143684 261480 180248 261508
rect 143684 261468 143690 261480
rect 180242 261468 180248 261480
rect 180300 261468 180306 261520
rect 171778 260856 171784 260908
rect 171836 260896 171842 260908
rect 191650 260896 191656 260908
rect 171836 260868 191656 260896
rect 171836 260856 171842 260868
rect 191650 260856 191656 260868
rect 191708 260856 191714 260908
rect 100754 260788 100760 260840
rect 100812 260828 100818 260840
rect 108206 260828 108212 260840
rect 100812 260800 108212 260828
rect 100812 260788 100818 260800
rect 108206 260788 108212 260800
rect 108264 260788 108270 260840
rect 255406 260788 255412 260840
rect 255464 260828 255470 260840
rect 287698 260828 287704 260840
rect 255464 260800 287704 260828
rect 255464 260788 255470 260800
rect 287698 260788 287704 260800
rect 287756 260788 287762 260840
rect 55122 260176 55128 260228
rect 55180 260216 55186 260228
rect 59354 260216 59360 260228
rect 55180 260188 59360 260216
rect 55180 260176 55186 260188
rect 59354 260176 59360 260188
rect 59412 260216 59418 260228
rect 66806 260216 66812 260228
rect 59412 260188 66812 260216
rect 59412 260176 59418 260188
rect 66806 260176 66812 260188
rect 66864 260176 66870 260228
rect 46750 260108 46756 260160
rect 46808 260148 46814 260160
rect 55858 260148 55864 260160
rect 46808 260120 55864 260148
rect 46808 260108 46814 260120
rect 55858 260108 55864 260120
rect 55916 260108 55922 260160
rect 57514 260108 57520 260160
rect 57572 260148 57578 260160
rect 66254 260148 66260 260160
rect 57572 260120 66260 260148
rect 57572 260108 57578 260120
rect 66254 260108 66260 260120
rect 66312 260108 66318 260160
rect 144178 260108 144184 260160
rect 144236 260148 144242 260160
rect 178678 260148 178684 260160
rect 144236 260120 178684 260148
rect 144236 260108 144242 260120
rect 178678 260108 178684 260120
rect 178736 260108 178742 260160
rect 289722 260108 289728 260160
rect 289780 260148 289786 260160
rect 582374 260148 582380 260160
rect 289780 260120 582380 260148
rect 289780 260108 289786 260120
rect 582374 260108 582380 260120
rect 582432 260108 582438 260160
rect 101214 259836 101220 259888
rect 101272 259876 101278 259888
rect 102778 259876 102784 259888
rect 101272 259848 102784 259876
rect 101272 259836 101278 259848
rect 102778 259836 102784 259848
rect 102836 259836 102842 259888
rect 174538 259428 174544 259480
rect 174596 259468 174602 259480
rect 191282 259468 191288 259480
rect 174596 259440 191288 259468
rect 174596 259428 174602 259440
rect 191282 259428 191288 259440
rect 191340 259428 191346 259480
rect 255406 259428 255412 259480
rect 255464 259468 255470 259480
rect 288526 259468 288532 259480
rect 255464 259440 288532 259468
rect 255464 259428 255470 259440
rect 288526 259428 288532 259440
rect 288584 259468 288590 259480
rect 289722 259468 289728 259480
rect 288584 259440 289728 259468
rect 288584 259428 288590 259440
rect 289722 259428 289728 259440
rect 289780 259428 289786 259480
rect 59262 259360 59268 259412
rect 59320 259400 59326 259412
rect 66438 259400 66444 259412
rect 59320 259372 66444 259400
rect 59320 259360 59326 259372
rect 66438 259360 66444 259372
rect 66496 259360 66502 259412
rect 100754 259360 100760 259412
rect 100812 259400 100818 259412
rect 126330 259400 126336 259412
rect 100812 259372 126336 259400
rect 100812 259360 100818 259372
rect 126330 259360 126336 259372
rect 126388 259360 126394 259412
rect 50614 258680 50620 258732
rect 50672 258720 50678 258732
rect 57606 258720 57612 258732
rect 50672 258692 57612 258720
rect 50672 258680 50678 258692
rect 57606 258680 57612 258692
rect 57664 258720 57670 258732
rect 66254 258720 66260 258732
rect 57664 258692 66260 258720
rect 57664 258680 57670 258692
rect 66254 258680 66260 258692
rect 66312 258680 66318 258732
rect 278682 258680 278688 258732
rect 278740 258720 278746 258732
rect 582466 258720 582472 258732
rect 278740 258692 582472 258720
rect 278740 258680 278746 258692
rect 582466 258680 582472 258692
rect 582524 258680 582530 258732
rect 100754 258204 100760 258256
rect 100812 258244 100818 258256
rect 105630 258244 105636 258256
rect 100812 258216 105636 258244
rect 100812 258204 100818 258216
rect 105630 258204 105636 258216
rect 105688 258204 105694 258256
rect 175918 258068 175924 258120
rect 175976 258108 175982 258120
rect 190454 258108 190460 258120
rect 175976 258080 190460 258108
rect 175976 258068 175982 258080
rect 190454 258068 190460 258080
rect 190512 258068 190518 258120
rect 255498 258068 255504 258120
rect 255556 258108 255562 258120
rect 277578 258108 277584 258120
rect 255556 258080 277584 258108
rect 255556 258068 255562 258080
rect 277578 258068 277584 258080
rect 277636 258108 277642 258120
rect 278682 258108 278688 258120
rect 277636 258080 278688 258108
rect 277636 258068 277642 258080
rect 278682 258068 278688 258080
rect 278740 258068 278746 258120
rect 190546 258000 190552 258052
rect 190604 258040 190610 258052
rect 193398 258040 193404 258052
rect 190604 258012 193404 258040
rect 190604 258000 190610 258012
rect 193398 258000 193404 258012
rect 193456 258000 193462 258052
rect 268102 258000 268108 258052
rect 268160 258040 268166 258052
rect 582834 258040 582840 258052
rect 268160 258012 582840 258040
rect 268160 258000 268166 258012
rect 582834 258000 582840 258012
rect 582892 258000 582898 258052
rect 100754 257388 100760 257440
rect 100812 257428 100818 257440
rect 101122 257428 101128 257440
rect 100812 257400 101128 257428
rect 100812 257388 100818 257400
rect 101122 257388 101128 257400
rect 101180 257428 101186 257440
rect 105538 257428 105544 257440
rect 101180 257400 105544 257428
rect 101180 257388 101186 257400
rect 105538 257388 105544 257400
rect 105596 257388 105602 257440
rect 113818 257388 113824 257440
rect 113876 257428 113882 257440
rect 138014 257428 138020 257440
rect 113876 257400 138020 257428
rect 113876 257388 113882 257400
rect 138014 257388 138020 257400
rect 138072 257388 138078 257440
rect 152550 257388 152556 257440
rect 152608 257428 152614 257440
rect 178678 257428 178684 257440
rect 152608 257400 178684 257428
rect 152608 257388 152614 257400
rect 178678 257388 178684 257400
rect 178736 257388 178742 257440
rect 50982 257320 50988 257372
rect 51040 257360 51046 257372
rect 59078 257360 59084 257372
rect 51040 257332 59084 257360
rect 51040 257320 51046 257332
rect 59078 257320 59084 257332
rect 59136 257360 59142 257372
rect 66806 257360 66812 257372
rect 59136 257332 66812 257360
rect 59136 257320 59142 257332
rect 66806 257320 66812 257332
rect 66864 257320 66870 257372
rect 137462 257320 137468 257372
rect 137520 257360 137526 257372
rect 173250 257360 173256 257372
rect 137520 257332 173256 257360
rect 137520 257320 137526 257332
rect 173250 257320 173256 257332
rect 173308 257320 173314 257372
rect 255314 257320 255320 257372
rect 255372 257360 255378 257372
rect 268102 257360 268108 257372
rect 255372 257332 268108 257360
rect 255372 257320 255378 257332
rect 268102 257320 268108 257332
rect 268160 257320 268166 257372
rect 185578 256708 185584 256760
rect 185636 256748 185642 256760
rect 191650 256748 191656 256760
rect 185636 256720 191656 256748
rect 185636 256708 185642 256720
rect 191650 256708 191656 256720
rect 191708 256708 191714 256760
rect 255498 256708 255504 256760
rect 255556 256748 255562 256760
rect 270770 256748 270776 256760
rect 255556 256720 270776 256748
rect 255556 256708 255562 256720
rect 270770 256708 270776 256720
rect 270828 256708 270834 256760
rect 101030 256640 101036 256692
rect 101088 256680 101094 256692
rect 141602 256680 141608 256692
rect 101088 256652 141608 256680
rect 101088 256640 101094 256652
rect 141602 256640 141608 256652
rect 141660 256640 141666 256692
rect 255406 256640 255412 256692
rect 255464 256680 255470 256692
rect 266630 256680 266636 256692
rect 255464 256652 266636 256680
rect 255464 256640 255470 256652
rect 266630 256640 266636 256652
rect 266688 256640 266694 256692
rect 39942 255960 39948 256012
rect 40000 256000 40006 256012
rect 51074 256000 51080 256012
rect 40000 255972 51080 256000
rect 40000 255960 40006 255972
rect 51074 255960 51080 255972
rect 51132 255960 51138 256012
rect 137370 255960 137376 256012
rect 137428 256000 137434 256012
rect 186958 256000 186964 256012
rect 137428 255972 186964 256000
rect 137428 255960 137434 255972
rect 186958 255960 186964 255972
rect 187016 255960 187022 256012
rect 273346 255960 273352 256012
rect 273404 256000 273410 256012
rect 580258 256000 580264 256012
rect 273404 255972 580264 256000
rect 273404 255960 273410 255972
rect 580258 255960 580264 255972
rect 580316 255960 580322 256012
rect 51074 255280 51080 255332
rect 51132 255320 51138 255332
rect 51994 255320 52000 255332
rect 51132 255292 52000 255320
rect 51132 255280 51138 255292
rect 51994 255280 52000 255292
rect 52052 255320 52058 255332
rect 66806 255320 66812 255332
rect 52052 255292 66812 255320
rect 52052 255280 52058 255292
rect 66806 255280 66812 255292
rect 66864 255280 66870 255332
rect 108942 255280 108948 255332
rect 109000 255320 109006 255332
rect 111886 255320 111892 255332
rect 109000 255292 111892 255320
rect 109000 255280 109006 255292
rect 111886 255280 111892 255292
rect 111944 255280 111950 255332
rect 181438 255280 181444 255332
rect 181496 255320 181502 255332
rect 190638 255320 190644 255332
rect 181496 255292 190644 255320
rect 181496 255280 181502 255292
rect 190638 255280 190644 255292
rect 190696 255280 190702 255332
rect 255498 255280 255504 255332
rect 255556 255320 255562 255332
rect 272058 255320 272064 255332
rect 255556 255292 272064 255320
rect 255556 255280 255562 255292
rect 272058 255280 272064 255292
rect 272116 255280 272122 255332
rect 3142 255212 3148 255264
rect 3200 255252 3206 255264
rect 10318 255252 10324 255264
rect 3200 255224 10324 255252
rect 3200 255212 3206 255224
rect 10318 255212 10324 255224
rect 10376 255212 10382 255264
rect 266722 255212 266728 255264
rect 266780 255252 266786 255264
rect 583018 255252 583024 255264
rect 266780 255224 583024 255252
rect 266780 255212 266786 255224
rect 583018 255212 583024 255224
rect 583076 255212 583082 255264
rect 109034 255144 109040 255196
rect 109092 255184 109098 255196
rect 113910 255184 113916 255196
rect 109092 255156 113916 255184
rect 109092 255144 109098 255156
rect 113910 255144 113916 255156
rect 113968 255144 113974 255196
rect 273622 255144 273628 255196
rect 273680 255184 273686 255196
rect 583386 255184 583392 255196
rect 273680 255156 583392 255184
rect 273680 255144 273686 255156
rect 583386 255144 583392 255156
rect 583444 255144 583450 255196
rect 255498 254600 255504 254652
rect 255556 254640 255562 254652
rect 266722 254640 266728 254652
rect 255556 254612 266728 254640
rect 255556 254600 255562 254612
rect 266722 254600 266728 254612
rect 266780 254600 266786 254652
rect 57790 254532 57796 254584
rect 57848 254572 57854 254584
rect 59170 254572 59176 254584
rect 57848 254544 59176 254572
rect 57848 254532 57854 254544
rect 59170 254532 59176 254544
rect 59228 254572 59234 254584
rect 66806 254572 66812 254584
rect 59228 254544 66812 254572
rect 59228 254532 59234 254544
rect 66806 254532 66812 254544
rect 66864 254532 66870 254584
rect 100754 254532 100760 254584
rect 100812 254572 100818 254584
rect 106642 254572 106648 254584
rect 100812 254544 106648 254572
rect 100812 254532 100818 254544
rect 106642 254532 106648 254544
rect 106700 254532 106706 254584
rect 121362 254532 121368 254584
rect 121420 254572 121426 254584
rect 184382 254572 184388 254584
rect 121420 254544 184388 254572
rect 121420 254532 121426 254544
rect 184382 254532 184388 254544
rect 184440 254532 184446 254584
rect 255406 254532 255412 254584
rect 255464 254572 255470 254584
rect 273622 254572 273628 254584
rect 255464 254544 273628 254572
rect 255464 254532 255470 254544
rect 273622 254532 273628 254544
rect 273680 254532 273686 254584
rect 100846 253920 100852 253972
rect 100904 253960 100910 253972
rect 109034 253960 109040 253972
rect 100904 253932 109040 253960
rect 100904 253920 100910 253932
rect 109034 253920 109040 253932
rect 109092 253920 109098 253972
rect 110414 253920 110420 253972
rect 110472 253960 110478 253972
rect 111058 253960 111064 253972
rect 110472 253932 111064 253960
rect 110472 253920 110478 253932
rect 111058 253920 111064 253932
rect 111116 253960 111122 253972
rect 151262 253960 151268 253972
rect 111116 253932 151268 253960
rect 111116 253920 111122 253932
rect 151262 253920 151268 253932
rect 151320 253920 151326 253972
rect 169110 253920 169116 253972
rect 169168 253960 169174 253972
rect 191650 253960 191656 253972
rect 169168 253932 191656 253960
rect 169168 253920 169174 253932
rect 191650 253920 191656 253932
rect 191708 253920 191714 253972
rect 63218 253852 63224 253904
rect 63276 253892 63282 253904
rect 66530 253892 66536 253904
rect 63276 253864 66536 253892
rect 63276 253852 63282 253864
rect 66530 253852 66536 253864
rect 66588 253852 66594 253904
rect 100754 253852 100760 253904
rect 100812 253892 100818 253904
rect 140774 253892 140780 253904
rect 100812 253864 140780 253892
rect 100812 253852 100818 253864
rect 140774 253852 140780 253864
rect 140832 253892 140838 253904
rect 141050 253892 141056 253904
rect 140832 253864 141056 253892
rect 140832 253852 140838 253864
rect 141050 253852 141056 253864
rect 141108 253852 141114 253904
rect 255590 253852 255596 253904
rect 255648 253892 255654 253904
rect 255958 253892 255964 253904
rect 255648 253864 255964 253892
rect 255648 253852 255654 253864
rect 255958 253852 255964 253864
rect 256016 253892 256022 253904
rect 583202 253892 583208 253904
rect 256016 253864 583208 253892
rect 256016 253852 256022 253864
rect 583202 253852 583208 253864
rect 583260 253852 583266 253904
rect 100846 253172 100852 253224
rect 100904 253212 100910 253224
rect 126422 253212 126428 253224
rect 100904 253184 126428 253212
rect 100904 253172 100910 253184
rect 126422 253172 126428 253184
rect 126480 253172 126486 253224
rect 255406 253172 255412 253224
rect 255464 253212 255470 253224
rect 269390 253212 269396 253224
rect 255464 253184 269396 253212
rect 255464 253172 255470 253184
rect 269390 253172 269396 253184
rect 269448 253212 269454 253224
rect 269758 253212 269764 253224
rect 269448 253184 269764 253212
rect 269448 253172 269454 253184
rect 269758 253172 269764 253184
rect 269816 253172 269822 253224
rect 186958 252560 186964 252612
rect 187016 252600 187022 252612
rect 191650 252600 191656 252612
rect 187016 252572 191656 252600
rect 187016 252560 187022 252572
rect 191650 252560 191656 252572
rect 191708 252560 191714 252612
rect 103330 251880 103336 251932
rect 103388 251920 103394 251932
rect 111794 251920 111800 251932
rect 103388 251892 111800 251920
rect 103388 251880 103394 251892
rect 111794 251880 111800 251892
rect 111852 251880 111858 251932
rect 256234 251880 256240 251932
rect 256292 251920 256298 251932
rect 256970 251920 256976 251932
rect 256292 251892 256976 251920
rect 256292 251880 256298 251892
rect 256970 251880 256976 251892
rect 257028 251920 257034 251932
rect 278038 251920 278044 251932
rect 257028 251892 278044 251920
rect 257028 251880 257034 251892
rect 278038 251880 278044 251892
rect 278096 251880 278102 251932
rect 106182 251812 106188 251864
rect 106240 251852 106246 251864
rect 115198 251852 115204 251864
rect 106240 251824 115204 251852
rect 106240 251812 106246 251824
rect 115198 251812 115204 251824
rect 115256 251852 115262 251864
rect 120074 251852 120080 251864
rect 115256 251824 120080 251852
rect 115256 251812 115262 251824
rect 120074 251812 120080 251824
rect 120132 251812 120138 251864
rect 263870 251812 263876 251864
rect 263928 251852 263934 251864
rect 583570 251852 583576 251864
rect 263928 251824 583576 251852
rect 263928 251812 263934 251824
rect 583570 251812 583576 251824
rect 583628 251812 583634 251864
rect 64782 251336 64788 251388
rect 64840 251376 64846 251388
rect 65978 251376 65984 251388
rect 64840 251348 65984 251376
rect 64840 251336 64846 251348
rect 65978 251336 65984 251348
rect 66036 251376 66042 251388
rect 66254 251376 66260 251388
rect 66036 251348 66260 251376
rect 66036 251336 66042 251348
rect 66254 251336 66260 251348
rect 66312 251336 66318 251388
rect 185670 251268 185676 251320
rect 185728 251308 185734 251320
rect 190822 251308 190828 251320
rect 185728 251280 190828 251308
rect 185728 251268 185734 251280
rect 190822 251268 190828 251280
rect 190880 251268 190886 251320
rect 255406 251268 255412 251320
rect 255464 251308 255470 251320
rect 263870 251308 263876 251320
rect 255464 251280 263876 251308
rect 255464 251268 255470 251280
rect 263870 251268 263876 251280
rect 263928 251268 263934 251320
rect 163498 251200 163504 251252
rect 163556 251240 163562 251252
rect 191650 251240 191656 251252
rect 163556 251212 191656 251240
rect 163556 251200 163562 251212
rect 191650 251200 191656 251212
rect 191708 251200 191714 251252
rect 58894 251132 58900 251184
rect 58952 251172 58958 251184
rect 61838 251172 61844 251184
rect 58952 251144 61844 251172
rect 58952 251132 58958 251144
rect 61838 251132 61844 251144
rect 61896 251132 61902 251184
rect 106274 251132 106280 251184
rect 106332 251172 106338 251184
rect 109678 251172 109684 251184
rect 106332 251144 109684 251172
rect 106332 251132 106338 251144
rect 109678 251132 109684 251144
rect 109736 251132 109742 251184
rect 57882 251064 57888 251116
rect 57940 251104 57946 251116
rect 66898 251104 66904 251116
rect 57940 251076 66904 251104
rect 57940 251064 57946 251076
rect 66898 251064 66904 251076
rect 66956 251064 66962 251116
rect 61010 250724 61016 250776
rect 61068 250764 61074 250776
rect 61378 250764 61384 250776
rect 61068 250736 61384 250764
rect 61068 250724 61074 250736
rect 61378 250724 61384 250736
rect 61436 250764 61442 250776
rect 66806 250764 66812 250776
rect 61436 250736 66812 250764
rect 61436 250724 61442 250736
rect 66806 250724 66812 250736
rect 66864 250724 66870 250776
rect 262490 250520 262496 250572
rect 262548 250560 262554 250572
rect 273346 250560 273352 250572
rect 262548 250532 273352 250560
rect 262548 250520 262554 250532
rect 273346 250520 273352 250532
rect 273404 250520 273410 250572
rect 101950 250452 101956 250504
rect 102008 250492 102014 250504
rect 114554 250492 114560 250504
rect 102008 250464 114560 250492
rect 102008 250452 102014 250464
rect 114554 250452 114560 250464
rect 114612 250452 114618 250504
rect 153838 250452 153844 250504
rect 153896 250492 153902 250504
rect 162118 250492 162124 250504
rect 153896 250464 162124 250492
rect 153896 250452 153902 250464
rect 162118 250452 162124 250464
rect 162176 250452 162182 250504
rect 164970 250452 164976 250504
rect 165028 250492 165034 250504
rect 192570 250492 192576 250504
rect 165028 250464 192576 250492
rect 165028 250452 165034 250464
rect 192570 250452 192576 250464
rect 192628 250452 192634 250504
rect 265250 250452 265256 250504
rect 265308 250492 265314 250504
rect 582374 250492 582380 250504
rect 265308 250464 582380 250492
rect 265308 250452 265314 250464
rect 582374 250452 582380 250464
rect 582432 250452 582438 250504
rect 255498 249840 255504 249892
rect 255556 249880 255562 249892
rect 262490 249880 262496 249892
rect 255556 249852 262496 249880
rect 255556 249840 255562 249852
rect 262490 249840 262496 249852
rect 262548 249840 262554 249892
rect 57882 249772 57888 249824
rect 57940 249812 57946 249824
rect 57940 249784 59308 249812
rect 57940 249772 57946 249784
rect 59280 249756 59308 249784
rect 100754 249772 100760 249824
rect 100812 249812 100818 249824
rect 106274 249812 106280 249824
rect 100812 249784 106280 249812
rect 100812 249772 100818 249784
rect 106274 249772 106280 249784
rect 106332 249772 106338 249824
rect 115382 249772 115388 249824
rect 115440 249812 115446 249824
rect 159542 249812 159548 249824
rect 115440 249784 159548 249812
rect 115440 249772 115446 249784
rect 159542 249772 159548 249784
rect 159600 249772 159606 249824
rect 170490 249772 170496 249824
rect 170548 249812 170554 249824
rect 191650 249812 191656 249824
rect 170548 249784 191656 249812
rect 170548 249772 170554 249784
rect 191650 249772 191656 249784
rect 191708 249772 191714 249824
rect 255406 249772 255412 249824
rect 255464 249812 255470 249824
rect 265250 249812 265256 249824
rect 255464 249784 265256 249812
rect 255464 249772 255470 249784
rect 265250 249772 265256 249784
rect 265308 249772 265314 249824
rect 59262 249704 59268 249756
rect 59320 249704 59326 249756
rect 100754 249636 100760 249688
rect 100812 249676 100818 249688
rect 101122 249676 101128 249688
rect 100812 249648 101128 249676
rect 100812 249636 100818 249648
rect 101122 249636 101128 249648
rect 101180 249636 101186 249688
rect 101674 249024 101680 249076
rect 101732 249064 101738 249076
rect 103330 249064 103336 249076
rect 101732 249036 103336 249064
rect 101732 249024 101738 249036
rect 103330 249024 103336 249036
rect 103388 249064 103394 249076
rect 140774 249064 140780 249076
rect 103388 249036 140780 249064
rect 103388 249024 103394 249036
rect 140774 249024 140780 249036
rect 140832 249024 140838 249076
rect 160830 249024 160836 249076
rect 160888 249064 160894 249076
rect 169202 249064 169208 249076
rect 160888 249036 169208 249064
rect 160888 249024 160894 249036
rect 169202 249024 169208 249036
rect 169260 249024 169266 249076
rect 192478 248520 192484 248532
rect 180766 248492 192484 248520
rect 55030 248412 55036 248464
rect 55088 248452 55094 248464
rect 57790 248452 57796 248464
rect 55088 248424 57796 248452
rect 55088 248412 55094 248424
rect 57790 248412 57796 248424
rect 57848 248452 57854 248464
rect 66806 248452 66812 248464
rect 57848 248424 66812 248452
rect 57848 248412 57854 248424
rect 66806 248412 66812 248424
rect 66864 248412 66870 248464
rect 106918 248412 106924 248464
rect 106976 248452 106982 248464
rect 180766 248452 180794 248492
rect 192478 248480 192484 248492
rect 192536 248480 192542 248532
rect 255406 248480 255412 248532
rect 255464 248520 255470 248532
rect 278038 248520 278044 248532
rect 255464 248492 278044 248520
rect 255464 248480 255470 248492
rect 278038 248480 278044 248492
rect 278096 248480 278102 248532
rect 106976 248424 180794 248452
rect 106976 248412 106982 248424
rect 188522 248412 188528 248464
rect 188580 248452 188586 248464
rect 191650 248452 191656 248464
rect 188580 248424 191656 248452
rect 188580 248412 188586 248424
rect 191650 248412 191656 248424
rect 191708 248412 191714 248464
rect 255314 248412 255320 248464
rect 255372 248452 255378 248464
rect 266630 248452 266636 248464
rect 255372 248424 266636 248452
rect 255372 248412 255378 248424
rect 266630 248412 266636 248424
rect 266688 248452 266694 248464
rect 582374 248452 582380 248464
rect 266688 248424 582380 248452
rect 266688 248412 266694 248424
rect 582374 248412 582380 248424
rect 582432 248412 582438 248464
rect 42702 248344 42708 248396
rect 42760 248384 42766 248396
rect 61930 248384 61936 248396
rect 42760 248356 61936 248384
rect 42760 248344 42766 248356
rect 61930 248344 61936 248356
rect 61988 248384 61994 248396
rect 66898 248384 66904 248396
rect 61988 248356 66904 248384
rect 61988 248344 61994 248356
rect 66898 248344 66904 248356
rect 66956 248344 66962 248396
rect 99190 248344 99196 248396
rect 99248 248384 99254 248396
rect 108942 248384 108948 248396
rect 99248 248356 108948 248384
rect 99248 248344 99254 248356
rect 108942 248344 108948 248356
rect 109000 248344 109006 248396
rect 108942 247732 108948 247784
rect 109000 247772 109006 247784
rect 166350 247772 166356 247784
rect 109000 247744 166356 247772
rect 109000 247732 109006 247744
rect 166350 247732 166356 247744
rect 166408 247732 166414 247784
rect 105538 247664 105544 247716
rect 105596 247704 105602 247716
rect 117314 247704 117320 247716
rect 105596 247676 117320 247704
rect 105596 247664 105602 247676
rect 117314 247664 117320 247676
rect 117372 247704 117378 247716
rect 177390 247704 177396 247716
rect 117372 247676 177396 247704
rect 117372 247664 117378 247676
rect 177390 247664 177396 247676
rect 177448 247664 177454 247716
rect 255406 247120 255412 247172
rect 255464 247160 255470 247172
rect 272150 247160 272156 247172
rect 255464 247132 272156 247160
rect 255464 247120 255470 247132
rect 272150 247120 272156 247132
rect 272208 247120 272214 247172
rect 184290 247052 184296 247104
rect 184348 247092 184354 247104
rect 191650 247092 191656 247104
rect 184348 247064 191656 247092
rect 184348 247052 184354 247064
rect 191650 247052 191656 247064
rect 191708 247052 191714 247104
rect 256418 247052 256424 247104
rect 256476 247092 256482 247104
rect 256878 247092 256884 247104
rect 256476 247064 256884 247092
rect 256476 247052 256482 247064
rect 256878 247052 256884 247064
rect 256936 247092 256942 247104
rect 582374 247092 582380 247104
rect 256936 247064 582380 247092
rect 256936 247052 256942 247064
rect 582374 247052 582380 247064
rect 582432 247052 582438 247104
rect 101122 246984 101128 247036
rect 101180 247024 101186 247036
rect 111058 247024 111064 247036
rect 101180 246996 111064 247024
rect 101180 246984 101186 246996
rect 111058 246984 111064 246996
rect 111116 246984 111122 247036
rect 56502 246304 56508 246356
rect 56560 246344 56566 246356
rect 66806 246344 66812 246356
rect 56560 246316 66812 246344
rect 56560 246304 56566 246316
rect 66806 246304 66812 246316
rect 66864 246304 66870 246356
rect 101030 246304 101036 246356
rect 101088 246344 101094 246356
rect 104802 246344 104808 246356
rect 101088 246316 104808 246344
rect 101088 246304 101094 246316
rect 104802 246304 104808 246316
rect 104860 246344 104866 246356
rect 128446 246344 128452 246356
rect 104860 246316 128452 246344
rect 104860 246304 104866 246316
rect 128446 246304 128452 246316
rect 128504 246304 128510 246356
rect 140774 246304 140780 246356
rect 140832 246344 140838 246356
rect 193674 246344 193680 246356
rect 140832 246316 193680 246344
rect 140832 246304 140838 246316
rect 193674 246304 193680 246316
rect 193732 246304 193738 246356
rect 255406 245692 255412 245744
rect 255464 245732 255470 245744
rect 287146 245732 287152 245744
rect 255464 245704 287152 245732
rect 255464 245692 255470 245704
rect 287146 245692 287152 245704
rect 287204 245692 287210 245744
rect 187234 245624 187240 245676
rect 187292 245664 187298 245676
rect 190638 245664 190644 245676
rect 187292 245636 190644 245664
rect 187292 245624 187298 245636
rect 190638 245624 190644 245636
rect 190696 245624 190702 245676
rect 48222 244944 48228 244996
rect 48280 244984 48286 244996
rect 57882 244984 57888 244996
rect 48280 244956 57888 244984
rect 48280 244944 48286 244956
rect 57882 244944 57888 244956
rect 57940 244944 57946 244996
rect 53650 244876 53656 244928
rect 53708 244916 53714 244928
rect 67542 244916 67548 244928
rect 53708 244888 67548 244916
rect 53708 244876 53714 244888
rect 67542 244876 67548 244888
rect 67600 244876 67606 244928
rect 102226 244876 102232 244928
rect 102284 244916 102290 244928
rect 113818 244916 113824 244928
rect 102284 244888 113824 244916
rect 102284 244876 102290 244888
rect 113818 244876 113824 244888
rect 113876 244876 113882 244928
rect 255498 244400 255504 244452
rect 255556 244440 255562 244452
rect 258166 244440 258172 244452
rect 255556 244412 258172 244440
rect 255556 244400 255562 244412
rect 258166 244400 258172 244412
rect 258224 244400 258230 244452
rect 108390 244264 108396 244316
rect 108448 244304 108454 244316
rect 165522 244304 165528 244316
rect 108448 244276 165528 244304
rect 108448 244264 108454 244276
rect 165522 244264 165528 244276
rect 165580 244264 165586 244316
rect 255406 244264 255412 244316
rect 255464 244304 255470 244316
rect 285766 244304 285772 244316
rect 255464 244276 285772 244304
rect 255464 244264 255470 244276
rect 285766 244264 285772 244276
rect 285824 244264 285830 244316
rect 69014 243516 69020 243568
rect 69072 243556 69078 243568
rect 169202 243556 169208 243568
rect 69072 243528 169208 243556
rect 69072 243516 69078 243528
rect 169202 243516 169208 243528
rect 169260 243516 169266 243568
rect 49510 242904 49516 242956
rect 49568 242944 49574 242956
rect 55030 242944 55036 242956
rect 49568 242916 55036 242944
rect 49568 242904 49574 242916
rect 55030 242904 55036 242916
rect 55088 242944 55094 242956
rect 66254 242944 66260 242956
rect 55088 242916 66260 242944
rect 55088 242904 55094 242916
rect 66254 242904 66260 242916
rect 66312 242904 66318 242956
rect 67818 242904 67824 242956
rect 67876 242944 67882 242956
rect 68462 242944 68468 242956
rect 67876 242916 68468 242944
rect 67876 242904 67882 242916
rect 68462 242904 68468 242916
rect 68520 242904 68526 242956
rect 108298 242904 108304 242956
rect 108356 242944 108362 242956
rect 161474 242944 161480 242956
rect 108356 242916 161480 242944
rect 108356 242904 108362 242916
rect 161474 242904 161480 242916
rect 161532 242944 161538 242956
rect 161532 242916 195652 242944
rect 161532 242904 161538 242916
rect 169294 242224 169300 242276
rect 169352 242264 169358 242276
rect 169352 242236 195284 242264
rect 169352 242224 169358 242236
rect 54846 242156 54852 242208
rect 54904 242196 54910 242208
rect 62114 242196 62120 242208
rect 54904 242168 62120 242196
rect 54904 242156 54910 242168
rect 62114 242156 62120 242168
rect 62172 242156 62178 242208
rect 153930 242156 153936 242208
rect 153988 242196 153994 242208
rect 153988 242168 180794 242196
rect 153988 242156 153994 242168
rect 96890 241748 96896 241800
rect 96948 241788 96954 241800
rect 99558 241788 99564 241800
rect 96948 241760 99564 241788
rect 96948 241748 96954 241760
rect 99558 241748 99564 241760
rect 99616 241748 99622 241800
rect 101030 241680 101036 241732
rect 101088 241720 101094 241732
rect 104158 241720 104164 241732
rect 101088 241692 104164 241720
rect 101088 241680 101094 241692
rect 104158 241680 104164 241692
rect 104216 241720 104222 241732
rect 107654 241720 107660 241732
rect 104216 241692 107660 241720
rect 104216 241680 104222 241692
rect 107654 241680 107660 241692
rect 107712 241680 107718 241732
rect 70946 241612 70952 241664
rect 71004 241652 71010 241664
rect 127710 241652 127716 241664
rect 71004 241624 127716 241652
rect 71004 241612 71010 241624
rect 127710 241612 127716 241624
rect 127768 241612 127774 241664
rect 154022 241584 154028 241596
rect 113146 241556 154028 241584
rect 66162 241476 66168 241528
rect 66220 241516 66226 241528
rect 69934 241516 69940 241528
rect 66220 241488 69940 241516
rect 66220 241476 66226 241488
rect 69934 241476 69940 241488
rect 69992 241476 69998 241528
rect 95326 241476 95332 241528
rect 95384 241516 95390 241528
rect 96200 241516 96206 241528
rect 95384 241488 96206 241516
rect 95384 241476 95390 241488
rect 96200 241476 96206 241488
rect 96258 241476 96264 241528
rect 52178 241408 52184 241460
rect 52236 241448 52242 241460
rect 76558 241448 76564 241460
rect 52236 241420 76564 241448
rect 52236 241408 52242 241420
rect 76558 241408 76564 241420
rect 76616 241448 76622 241460
rect 76880 241448 76886 241460
rect 76616 241420 76886 241448
rect 76616 241408 76622 241420
rect 76880 241408 76886 241420
rect 76938 241408 76944 241460
rect 81296 241408 81302 241460
rect 81354 241448 81360 241460
rect 112438 241448 112444 241460
rect 81354 241420 112444 241448
rect 81354 241408 81360 241420
rect 112438 241408 112444 241420
rect 112496 241448 112502 241460
rect 113146 241448 113174 241556
rect 154022 241544 154028 241556
rect 154080 241544 154086 241596
rect 180766 241584 180794 242168
rect 195256 241664 195284 242236
rect 195624 241664 195652 242916
rect 193582 241612 193588 241664
rect 193640 241652 193646 241664
rect 193766 241652 193772 241664
rect 193640 241624 193772 241652
rect 193640 241612 193646 241624
rect 193766 241612 193772 241624
rect 193824 241612 193830 241664
rect 195238 241612 195244 241664
rect 195296 241612 195302 241664
rect 195606 241612 195612 241664
rect 195664 241612 195670 241664
rect 249058 241612 249064 241664
rect 249116 241652 249122 241664
rect 256970 241652 256976 241664
rect 249116 241624 256976 241652
rect 249116 241612 249122 241624
rect 256970 241612 256976 241624
rect 257028 241612 257034 241664
rect 196618 241584 196624 241596
rect 180766 241556 196624 241584
rect 196618 241544 196624 241556
rect 196676 241544 196682 241596
rect 255682 241476 255688 241528
rect 255740 241516 255746 241528
rect 256142 241516 256148 241528
rect 255740 241488 256148 241516
rect 255740 241476 255746 241488
rect 256142 241476 256148 241488
rect 256200 241516 256206 241528
rect 582558 241516 582564 241528
rect 256200 241488 582564 241516
rect 256200 241476 256206 241488
rect 582558 241476 582564 241488
rect 582616 241476 582622 241528
rect 112496 241420 113174 241448
rect 112496 241408 112502 241420
rect 181622 241408 181628 241460
rect 181680 241448 181686 241460
rect 252830 241448 252836 241460
rect 181680 241420 252836 241448
rect 181680 241408 181686 241420
rect 252830 241408 252836 241420
rect 252888 241408 252894 241460
rect 256050 241408 256056 241460
rect 256108 241448 256114 241460
rect 565078 241448 565084 241460
rect 256108 241420 565084 241448
rect 256108 241408 256114 241420
rect 565078 241408 565084 241420
rect 565136 241408 565142 241460
rect 95878 241340 95884 241392
rect 95936 241380 95942 241392
rect 100018 241380 100024 241392
rect 95936 241352 100024 241380
rect 95936 241340 95942 241352
rect 100018 241340 100024 241352
rect 100076 241340 100082 241392
rect 165522 241340 165528 241392
rect 165580 241380 165586 241392
rect 199102 241380 199108 241392
rect 165580 241352 199108 241380
rect 165580 241340 165586 241352
rect 199102 241340 199108 241352
rect 199160 241340 199166 241392
rect 3510 241204 3516 241256
rect 3568 241244 3574 241256
rect 7558 241244 7564 241256
rect 3568 241216 7564 241244
rect 3568 241204 3574 241216
rect 7558 241204 7564 241216
rect 7616 241204 7622 241256
rect 64506 240728 64512 240780
rect 64564 240768 64570 240780
rect 77938 240768 77944 240780
rect 64564 240740 77944 240768
rect 64564 240728 64570 240740
rect 77938 240728 77944 240740
rect 77996 240728 78002 240780
rect 116670 240728 116676 240780
rect 116728 240768 116734 240780
rect 155402 240768 155408 240780
rect 116728 240740 155408 240768
rect 116728 240728 116734 240740
rect 155402 240728 155408 240740
rect 155460 240728 155466 240780
rect 224126 240728 224132 240780
rect 224184 240768 224190 240780
rect 256694 240768 256700 240780
rect 224184 240740 256700 240768
rect 224184 240728 224190 240740
rect 256694 240728 256700 240740
rect 256752 240728 256758 240780
rect 86218 240048 86224 240100
rect 86276 240088 86282 240100
rect 87046 240088 87052 240100
rect 86276 240060 87052 240088
rect 86276 240048 86282 240060
rect 87046 240048 87052 240060
rect 87104 240048 87110 240100
rect 98270 240048 98276 240100
rect 98328 240088 98334 240100
rect 197538 240088 197544 240100
rect 98328 240060 197544 240088
rect 98328 240048 98334 240060
rect 197538 240048 197544 240060
rect 197596 240088 197602 240100
rect 197998 240088 198004 240100
rect 197596 240060 198004 240088
rect 197596 240048 197602 240060
rect 197998 240048 198004 240060
rect 198056 240048 198062 240100
rect 242158 240048 242164 240100
rect 242216 240088 242222 240100
rect 242894 240088 242900 240100
rect 242216 240060 242900 240088
rect 242216 240048 242222 240060
rect 242894 240048 242900 240060
rect 242952 240048 242958 240100
rect 243538 240048 243544 240100
rect 243596 240088 243602 240100
rect 244550 240088 244556 240100
rect 243596 240060 244556 240088
rect 243596 240048 243602 240060
rect 244550 240048 244556 240060
rect 244608 240048 244614 240100
rect 251082 240048 251088 240100
rect 251140 240088 251146 240100
rect 254118 240088 254124 240100
rect 251140 240060 254124 240088
rect 251140 240048 251146 240060
rect 254118 240048 254124 240060
rect 254176 240048 254182 240100
rect 254762 240048 254768 240100
rect 254820 240088 254826 240100
rect 256694 240088 256700 240100
rect 254820 240060 256700 240088
rect 254820 240048 254826 240060
rect 256694 240048 256700 240060
rect 256752 240048 256758 240100
rect 45462 239980 45468 240032
rect 45520 240020 45526 240032
rect 71774 240020 71780 240032
rect 45520 239992 71780 240020
rect 45520 239980 45526 239992
rect 71774 239980 71780 239992
rect 71832 240020 71838 240032
rect 72510 240020 72516 240032
rect 71832 239992 72516 240020
rect 71832 239980 71838 239992
rect 72510 239980 72516 239992
rect 72568 239980 72574 240032
rect 77386 239980 77392 240032
rect 77444 240020 77450 240032
rect 82998 240020 83004 240032
rect 77444 239992 83004 240020
rect 77444 239980 77450 239992
rect 82998 239980 83004 239992
rect 83056 239980 83062 240032
rect 75914 239912 75920 239964
rect 75972 239952 75978 239964
rect 77478 239952 77484 239964
rect 75972 239924 77484 239952
rect 75972 239912 75978 239924
rect 77478 239912 77484 239924
rect 77536 239912 77542 239964
rect 88518 239436 88524 239488
rect 88576 239476 88582 239488
rect 97994 239476 98000 239488
rect 88576 239448 98000 239476
rect 88576 239436 88582 239448
rect 97994 239436 98000 239448
rect 98052 239436 98058 239488
rect 234798 239436 234804 239488
rect 234856 239476 234862 239488
rect 237466 239476 237472 239488
rect 234856 239448 237472 239476
rect 234856 239436 234862 239448
rect 237466 239436 237472 239448
rect 237524 239436 237530 239488
rect 74258 239368 74264 239420
rect 74316 239408 74322 239420
rect 167730 239408 167736 239420
rect 74316 239380 167736 239408
rect 74316 239368 74322 239380
rect 167730 239368 167736 239380
rect 167788 239408 167794 239420
rect 202414 239408 202420 239420
rect 167788 239380 202420 239408
rect 167788 239368 167794 239380
rect 202414 239368 202420 239380
rect 202472 239368 202478 239420
rect 74902 238864 74908 238876
rect 70320 238836 74908 238864
rect 41322 238688 41328 238740
rect 41380 238728 41386 238740
rect 69658 238728 69664 238740
rect 41380 238700 69664 238728
rect 41380 238688 41386 238700
rect 69658 238688 69664 238700
rect 69716 238728 69722 238740
rect 70320 238728 70348 238836
rect 74902 238824 74908 238836
rect 74960 238824 74966 238876
rect 226978 238756 226984 238808
rect 227036 238796 227042 238808
rect 231578 238796 231584 238808
rect 227036 238768 231584 238796
rect 227036 238756 227042 238768
rect 231578 238756 231584 238768
rect 231636 238756 231642 238808
rect 244918 238756 244924 238808
rect 244976 238796 244982 238808
rect 253014 238796 253020 238808
rect 244976 238768 253020 238796
rect 244976 238756 244982 238768
rect 253014 238756 253020 238768
rect 253072 238756 253078 238808
rect 69716 238700 70348 238728
rect 69716 238688 69722 238700
rect 80330 238688 80336 238740
rect 80388 238728 80394 238740
rect 108390 238728 108396 238740
rect 80388 238700 108396 238728
rect 80388 238688 80394 238700
rect 108390 238688 108396 238700
rect 108448 238688 108454 238740
rect 188430 238688 188436 238740
rect 188488 238728 188494 238740
rect 221458 238728 221464 238740
rect 188488 238700 221464 238728
rect 188488 238688 188494 238700
rect 221458 238688 221464 238700
rect 221516 238688 221522 238740
rect 81526 238620 81532 238672
rect 81584 238660 81590 238672
rect 106918 238660 106924 238672
rect 81584 238632 106924 238660
rect 81584 238620 81590 238632
rect 106918 238620 106924 238632
rect 106976 238620 106982 238672
rect 193030 238144 193036 238196
rect 193088 238184 193094 238196
rect 198826 238184 198832 238196
rect 193088 238156 198832 238184
rect 193088 238144 193094 238156
rect 198826 238144 198832 238156
rect 198884 238144 198890 238196
rect 63126 238076 63132 238128
rect 63184 238116 63190 238128
rect 72418 238116 72424 238128
rect 63184 238088 72424 238116
rect 63184 238076 63190 238088
rect 72418 238076 72424 238088
rect 72476 238076 72482 238128
rect 125502 238076 125508 238128
rect 125560 238116 125566 238128
rect 188614 238116 188620 238128
rect 125560 238088 188620 238116
rect 125560 238076 125566 238088
rect 188614 238076 188620 238088
rect 188672 238076 188678 238128
rect 69842 238008 69848 238060
rect 69900 238048 69906 238060
rect 79318 238048 79324 238060
rect 69900 238020 79324 238048
rect 69900 238008 69906 238020
rect 79318 238008 79324 238020
rect 79376 238008 79382 238060
rect 107562 238008 107568 238060
rect 107620 238048 107626 238060
rect 187142 238048 187148 238060
rect 107620 238020 187148 238048
rect 107620 238008 107626 238020
rect 187142 238008 187148 238020
rect 187200 238008 187206 238060
rect 204898 238008 204904 238060
rect 204956 238048 204962 238060
rect 253934 238048 253940 238060
rect 204956 238020 253940 238048
rect 204956 238008 204962 238020
rect 253934 238008 253940 238020
rect 253992 238008 253998 238060
rect 50798 237396 50804 237448
rect 50856 237436 50862 237448
rect 52362 237436 52368 237448
rect 50856 237408 52368 237436
rect 50856 237396 50862 237408
rect 52362 237396 52368 237408
rect 52420 237396 52426 237448
rect 222102 237396 222108 237448
rect 222160 237436 222166 237448
rect 227806 237436 227812 237448
rect 222160 237408 227812 237436
rect 222160 237396 222166 237408
rect 227806 237396 227812 237408
rect 227864 237396 227870 237448
rect 48038 237328 48044 237380
rect 48096 237368 48102 237380
rect 75914 237368 75920 237380
rect 48096 237340 75920 237368
rect 48096 237328 48102 237340
rect 75914 237328 75920 237340
rect 75972 237368 75978 237380
rect 77202 237368 77208 237380
rect 75972 237340 77208 237368
rect 75972 237328 75978 237340
rect 77202 237328 77208 237340
rect 77260 237328 77266 237380
rect 184382 237328 184388 237380
rect 184440 237368 184446 237380
rect 208854 237368 208860 237380
rect 184440 237340 208860 237368
rect 184440 237328 184446 237340
rect 208854 237328 208860 237340
rect 208912 237328 208918 237380
rect 55858 237260 55864 237312
rect 55916 237300 55922 237312
rect 80054 237300 80060 237312
rect 55916 237272 80060 237300
rect 55916 237260 55922 237272
rect 80054 237260 80060 237272
rect 80112 237260 80118 237312
rect 97994 236716 98000 236768
rect 98052 236756 98058 236768
rect 106182 236756 106188 236768
rect 98052 236728 106188 236756
rect 98052 236716 98058 236728
rect 106182 236716 106188 236728
rect 106240 236756 106246 236768
rect 121454 236756 121460 236768
rect 106240 236728 121460 236756
rect 106240 236716 106246 236728
rect 121454 236716 121460 236728
rect 121512 236716 121518 236768
rect 76834 236648 76840 236700
rect 76892 236688 76898 236700
rect 95234 236688 95240 236700
rect 76892 236660 95240 236688
rect 76892 236648 76898 236660
rect 95234 236648 95240 236660
rect 95292 236648 95298 236700
rect 111702 236648 111708 236700
rect 111760 236688 111766 236700
rect 181530 236688 181536 236700
rect 111760 236660 181536 236688
rect 111760 236648 111766 236660
rect 181530 236648 181536 236660
rect 181588 236648 181594 236700
rect 193214 236648 193220 236700
rect 193272 236688 193278 236700
rect 206278 236688 206284 236700
rect 193272 236660 206284 236688
rect 193272 236648 193278 236660
rect 206278 236648 206284 236660
rect 206336 236648 206342 236700
rect 211062 236648 211068 236700
rect 211120 236688 211126 236700
rect 256142 236688 256148 236700
rect 211120 236660 256148 236688
rect 211120 236648 211126 236660
rect 256142 236648 256148 236660
rect 256200 236648 256206 236700
rect 103422 236240 103428 236292
rect 103480 236280 103486 236292
rect 103698 236280 103704 236292
rect 103480 236252 103704 236280
rect 103480 236240 103486 236252
rect 103698 236240 103704 236252
rect 103756 236240 103762 236292
rect 80054 235968 80060 236020
rect 80112 236008 80118 236020
rect 80698 236008 80704 236020
rect 80112 235980 80704 236008
rect 80112 235968 80118 235980
rect 80698 235968 80704 235980
rect 80756 235968 80762 236020
rect 97810 235968 97816 236020
rect 97868 236008 97874 236020
rect 99466 236008 99472 236020
rect 97868 235980 99472 236008
rect 97868 235968 97874 235980
rect 99466 235968 99472 235980
rect 99524 235968 99530 236020
rect 108942 235968 108948 236020
rect 109000 236008 109006 236020
rect 109126 236008 109132 236020
rect 109000 235980 109132 236008
rect 109000 235968 109006 235980
rect 109126 235968 109132 235980
rect 109184 235968 109190 236020
rect 208394 235968 208400 236020
rect 208452 236008 208458 236020
rect 208854 236008 208860 236020
rect 208452 235980 208860 236008
rect 208452 235968 208458 235980
rect 208854 235968 208860 235980
rect 208912 235968 208918 236020
rect 81434 235900 81440 235952
rect 81492 235940 81498 235952
rect 105538 235940 105544 235952
rect 81492 235912 105544 235940
rect 81492 235900 81498 235912
rect 105538 235900 105544 235912
rect 105596 235900 105602 235952
rect 170582 235900 170588 235952
rect 170640 235940 170646 235952
rect 179414 235940 179420 235952
rect 170640 235912 179420 235940
rect 170640 235900 170646 235912
rect 179414 235900 179420 235912
rect 179472 235900 179478 235952
rect 192570 235900 192576 235952
rect 192628 235940 192634 235952
rect 200114 235940 200120 235952
rect 192628 235912 200120 235940
rect 192628 235900 192634 235912
rect 200114 235900 200120 235912
rect 200172 235940 200178 235952
rect 200758 235940 200764 235952
rect 200172 235912 200764 235940
rect 200172 235900 200178 235912
rect 200758 235900 200764 235912
rect 200816 235900 200822 235952
rect 82998 235832 83004 235884
rect 83056 235872 83062 235884
rect 83918 235872 83924 235884
rect 83056 235844 83924 235872
rect 83056 235832 83062 235844
rect 83918 235832 83924 235844
rect 83976 235872 83982 235884
rect 102134 235872 102140 235884
rect 83976 235844 102140 235872
rect 83976 235832 83982 235844
rect 102134 235832 102140 235844
rect 102192 235832 102198 235884
rect 43990 235220 43996 235272
rect 44048 235260 44054 235272
rect 56502 235260 56508 235272
rect 44048 235232 56508 235260
rect 44048 235220 44054 235232
rect 56502 235220 56508 235232
rect 56560 235260 56566 235272
rect 77570 235260 77576 235272
rect 56560 235232 77576 235260
rect 56560 235220 56566 235232
rect 77570 235220 77576 235232
rect 77628 235220 77634 235272
rect 186222 235220 186228 235272
rect 186280 235260 186286 235272
rect 195146 235260 195152 235272
rect 186280 235232 195152 235260
rect 186280 235220 186286 235232
rect 195146 235220 195152 235232
rect 195204 235220 195210 235272
rect 200758 235220 200764 235272
rect 200816 235260 200822 235272
rect 255958 235260 255964 235272
rect 200816 235232 255964 235260
rect 200816 235220 200822 235232
rect 255958 235220 255964 235232
rect 256016 235220 256022 235272
rect 105630 234608 105636 234660
rect 105688 234648 105694 234660
rect 105814 234648 105820 234660
rect 105688 234620 105820 234648
rect 105688 234608 105694 234620
rect 105814 234608 105820 234620
rect 105872 234648 105878 234660
rect 115934 234648 115940 234660
rect 105872 234620 115940 234648
rect 105872 234608 105878 234620
rect 115934 234608 115940 234620
rect 115992 234608 115998 234660
rect 195238 234608 195244 234660
rect 195296 234648 195302 234660
rect 224218 234648 224224 234660
rect 195296 234620 224224 234648
rect 195296 234608 195302 234620
rect 224218 234608 224224 234620
rect 224276 234608 224282 234660
rect 73154 234540 73160 234592
rect 73212 234580 73218 234592
rect 108298 234580 108304 234592
rect 73212 234552 108304 234580
rect 73212 234540 73218 234552
rect 108298 234540 108304 234552
rect 108356 234540 108362 234592
rect 176010 234540 176016 234592
rect 176068 234580 176074 234592
rect 267826 234580 267832 234592
rect 176068 234552 267832 234580
rect 176068 234540 176074 234552
rect 267826 234540 267832 234552
rect 267884 234540 267890 234592
rect 83918 234404 83924 234456
rect 83976 234444 83982 234456
rect 84102 234444 84108 234456
rect 83976 234416 84108 234444
rect 83976 234404 83982 234416
rect 84102 234404 84108 234416
rect 84160 234404 84166 234456
rect 61654 233860 61660 233912
rect 61712 233900 61718 233912
rect 75178 233900 75184 233912
rect 61712 233872 75184 233900
rect 61712 233860 61718 233872
rect 75178 233860 75184 233872
rect 75236 233860 75242 233912
rect 97902 233860 97908 233912
rect 97960 233900 97966 233912
rect 98178 233900 98184 233912
rect 97960 233872 98184 233900
rect 97960 233860 97966 233872
rect 98178 233860 98184 233872
rect 98236 233860 98242 233912
rect 220722 233860 220728 233912
rect 220780 233900 220786 233912
rect 229922 233900 229928 233912
rect 220780 233872 229928 233900
rect 220780 233860 220786 233872
rect 229922 233860 229928 233872
rect 229980 233860 229986 233912
rect 278038 233248 278044 233300
rect 278096 233288 278102 233300
rect 580166 233288 580172 233300
rect 278096 233260 580172 233288
rect 278096 233248 278102 233260
rect 580166 233248 580172 233260
rect 580224 233248 580230 233300
rect 65886 233180 65892 233232
rect 65944 233220 65950 233232
rect 67634 233220 67640 233232
rect 65944 233192 67640 233220
rect 65944 233180 65950 233192
rect 67634 233180 67640 233192
rect 67692 233180 67698 233232
rect 82906 233180 82912 233232
rect 82964 233220 82970 233232
rect 118694 233220 118700 233232
rect 82964 233192 118700 233220
rect 82964 233180 82970 233192
rect 118694 233180 118700 233192
rect 118752 233180 118758 233232
rect 119338 233180 119344 233232
rect 119396 233220 119402 233232
rect 124214 233220 124220 233232
rect 119396 233192 124220 233220
rect 119396 233180 119402 233192
rect 124214 233180 124220 233192
rect 124272 233180 124278 233232
rect 177390 233180 177396 233232
rect 177448 233220 177454 233232
rect 177942 233220 177948 233232
rect 177448 233192 177948 233220
rect 177448 233180 177454 233192
rect 177942 233180 177948 233192
rect 178000 233220 178006 233232
rect 216950 233220 216956 233232
rect 178000 233192 216956 233220
rect 178000 233180 178006 233192
rect 216950 233180 216956 233192
rect 217008 233180 217014 233232
rect 58986 233112 58992 233164
rect 59044 233152 59050 233164
rect 86218 233152 86224 233164
rect 59044 233124 86224 233152
rect 59044 233112 59050 233124
rect 86218 233112 86224 233124
rect 86276 233112 86282 233164
rect 217318 232568 217324 232620
rect 217376 232608 217382 232620
rect 225046 232608 225052 232620
rect 217376 232580 225052 232608
rect 217376 232568 217382 232580
rect 225046 232568 225052 232580
rect 225104 232568 225110 232620
rect 234614 232568 234620 232620
rect 234672 232608 234678 232620
rect 256970 232608 256976 232620
rect 234672 232580 256976 232608
rect 234672 232568 234678 232580
rect 256970 232568 256976 232580
rect 257028 232568 257034 232620
rect 91094 232500 91100 232552
rect 91152 232540 91158 232552
rect 119338 232540 119344 232552
rect 91152 232512 119344 232540
rect 91152 232500 91158 232512
rect 119338 232500 119344 232512
rect 119396 232500 119402 232552
rect 206922 232500 206928 232552
rect 206980 232540 206986 232552
rect 236454 232540 236460 232552
rect 206980 232512 236460 232540
rect 206980 232500 206986 232512
rect 236454 232500 236460 232512
rect 236512 232500 236518 232552
rect 240778 232500 240784 232552
rect 240836 232540 240842 232552
rect 255314 232540 255320 232552
rect 240836 232512 255320 232540
rect 240836 232500 240842 232512
rect 255314 232500 255320 232512
rect 255372 232500 255378 232552
rect 76006 231752 76012 231804
rect 76064 231792 76070 231804
rect 110690 231792 110696 231804
rect 76064 231764 110696 231792
rect 76064 231752 76070 231764
rect 110690 231752 110696 231764
rect 110748 231752 110754 231804
rect 180242 231752 180248 231804
rect 180300 231792 180306 231804
rect 260834 231792 260840 231804
rect 180300 231764 260840 231792
rect 180300 231752 180306 231764
rect 260834 231752 260840 231764
rect 260892 231792 260898 231804
rect 261202 231792 261208 231804
rect 260892 231764 261208 231792
rect 260892 231752 260898 231764
rect 261202 231752 261208 231764
rect 261260 231752 261266 231804
rect 272058 231752 272064 231804
rect 272116 231792 272122 231804
rect 272334 231792 272340 231804
rect 272116 231764 272340 231792
rect 272116 231752 272122 231764
rect 272334 231752 272340 231764
rect 272392 231792 272398 231804
rect 582742 231792 582748 231804
rect 272392 231764 582748 231792
rect 272392 231752 272398 231764
rect 582742 231752 582748 231764
rect 582800 231752 582806 231804
rect 154022 231684 154028 231736
rect 154080 231724 154086 231736
rect 205634 231724 205640 231736
rect 154080 231696 205640 231724
rect 154080 231684 154086 231696
rect 205634 231684 205640 231696
rect 205692 231684 205698 231736
rect 77202 231072 77208 231124
rect 77260 231112 77266 231124
rect 108390 231112 108396 231124
rect 77260 231084 108396 231112
rect 77260 231072 77266 231084
rect 108390 231072 108396 231084
rect 108448 231072 108454 231124
rect 110690 231072 110696 231124
rect 110748 231112 110754 231124
rect 153194 231112 153200 231124
rect 110748 231084 153200 231112
rect 110748 231072 110754 231084
rect 153194 231072 153200 231084
rect 153252 231072 153258 231124
rect 208486 231072 208492 231124
rect 208544 231112 208550 231124
rect 218606 231112 218612 231124
rect 208544 231084 218612 231112
rect 208544 231072 208550 231084
rect 218606 231072 218612 231084
rect 218664 231072 218670 231124
rect 255958 231072 255964 231124
rect 256016 231112 256022 231124
rect 272334 231112 272340 231124
rect 256016 231084 272340 231112
rect 256016 231072 256022 231084
rect 272334 231072 272340 231084
rect 272392 231072 272398 231124
rect 205634 230936 205640 230988
rect 205692 230976 205698 230988
rect 206370 230976 206376 230988
rect 205692 230948 206376 230976
rect 205692 230936 205698 230948
rect 206370 230936 206376 230948
rect 206428 230936 206434 230988
rect 191190 230392 191196 230444
rect 191248 230432 191254 230444
rect 212074 230432 212080 230444
rect 191248 230404 212080 230432
rect 191248 230392 191254 230404
rect 212074 230392 212080 230404
rect 212132 230392 212138 230444
rect 220998 230392 221004 230444
rect 221056 230432 221062 230444
rect 276198 230432 276204 230444
rect 221056 230404 276204 230432
rect 221056 230392 221062 230404
rect 276198 230392 276204 230404
rect 276256 230392 276262 230444
rect 60458 229780 60464 229832
rect 60516 229820 60522 229832
rect 76742 229820 76748 229832
rect 60516 229792 76748 229820
rect 60516 229780 60522 229792
rect 76742 229780 76748 229792
rect 76800 229780 76806 229832
rect 48038 229712 48044 229764
rect 48096 229752 48102 229764
rect 69474 229752 69480 229764
rect 48096 229724 69480 229752
rect 48096 229712 48102 229724
rect 69474 229712 69480 229724
rect 69532 229712 69538 229764
rect 72510 229712 72516 229764
rect 72568 229752 72574 229764
rect 86862 229752 86868 229764
rect 72568 229724 86868 229752
rect 72568 229712 72574 229724
rect 86862 229712 86868 229724
rect 86920 229752 86926 229764
rect 224126 229752 224132 229764
rect 86920 229724 224132 229752
rect 86920 229712 86926 229724
rect 224126 229712 224132 229724
rect 224184 229712 224190 229764
rect 224218 229712 224224 229764
rect 224276 229752 224282 229764
rect 238754 229752 238760 229764
rect 224276 229724 238760 229752
rect 224276 229712 224282 229724
rect 238754 229712 238760 229724
rect 238812 229752 238818 229764
rect 245010 229752 245016 229764
rect 238812 229724 245016 229752
rect 238812 229712 238818 229724
rect 245010 229712 245016 229724
rect 245068 229712 245074 229764
rect 256878 229712 256884 229764
rect 256936 229752 256942 229764
rect 272150 229752 272156 229764
rect 256936 229724 272156 229752
rect 256936 229712 256942 229724
rect 272150 229712 272156 229724
rect 272208 229752 272214 229764
rect 580258 229752 580264 229764
rect 272208 229724 580264 229752
rect 272208 229712 272214 229724
rect 580258 229712 580264 229724
rect 580316 229712 580322 229764
rect 102778 229032 102784 229084
rect 102836 229072 102842 229084
rect 273530 229072 273536 229084
rect 102836 229044 273536 229072
rect 102836 229032 102842 229044
rect 273530 229032 273536 229044
rect 273588 229032 273594 229084
rect 61838 228964 61844 229016
rect 61896 229004 61902 229016
rect 160094 229004 160100 229016
rect 61896 228976 160100 229004
rect 61896 228964 61902 228976
rect 160094 228964 160100 228976
rect 160152 229004 160158 229016
rect 160830 229004 160836 229016
rect 160152 228976 160836 229004
rect 160152 228964 160158 228976
rect 160830 228964 160836 228976
rect 160888 228964 160894 229016
rect 202782 228352 202788 228404
rect 202840 228392 202846 228404
rect 239674 228392 239680 228404
rect 202840 228364 239680 228392
rect 202840 228352 202846 228364
rect 239674 228352 239680 228364
rect 239732 228352 239738 228404
rect 258718 228352 258724 228404
rect 258776 228392 258782 228404
rect 269390 228392 269396 228404
rect 258776 228364 269396 228392
rect 258776 228352 258782 228364
rect 269390 228352 269396 228364
rect 269448 228352 269454 228404
rect 128354 227672 128360 227724
rect 128412 227712 128418 227724
rect 265158 227712 265164 227724
rect 128412 227684 265164 227712
rect 128412 227672 128418 227684
rect 265158 227672 265164 227684
rect 265216 227672 265222 227724
rect 270770 227672 270776 227724
rect 270828 227712 270834 227724
rect 582650 227712 582656 227724
rect 270828 227684 582656 227712
rect 270828 227672 270834 227684
rect 582650 227672 582656 227684
rect 582708 227672 582714 227724
rect 159542 227604 159548 227656
rect 159600 227644 159606 227656
rect 160002 227644 160008 227656
rect 159600 227616 160008 227644
rect 159600 227604 159606 227616
rect 160002 227604 160008 227616
rect 160060 227644 160066 227656
rect 249058 227644 249064 227656
rect 160060 227616 249064 227644
rect 160060 227604 160066 227616
rect 249058 227604 249064 227616
rect 249116 227604 249122 227656
rect 95142 226992 95148 227044
rect 95200 227032 95206 227044
rect 122650 227032 122656 227044
rect 95200 227004 122656 227032
rect 95200 226992 95206 227004
rect 122650 226992 122656 227004
rect 122708 227032 122714 227044
rect 128354 227032 128360 227044
rect 122708 227004 128360 227032
rect 122708 226992 122714 227004
rect 128354 226992 128360 227004
rect 128412 226992 128418 227044
rect 256142 226992 256148 227044
rect 256200 227032 256206 227044
rect 270770 227032 270776 227044
rect 256200 227004 270776 227032
rect 256200 226992 256206 227004
rect 270770 226992 270776 227004
rect 270828 226992 270834 227044
rect 59078 226244 59084 226296
rect 59136 226284 59142 226296
rect 160922 226284 160928 226296
rect 59136 226256 160928 226284
rect 59136 226244 59142 226256
rect 160922 226244 160928 226256
rect 160980 226244 160986 226296
rect 173250 226244 173256 226296
rect 173308 226284 173314 226296
rect 263870 226284 263876 226296
rect 173308 226256 263876 226284
rect 173308 226244 173314 226256
rect 263870 226244 263876 226256
rect 263928 226244 263934 226296
rect 95142 225564 95148 225616
rect 95200 225604 95206 225616
rect 104894 225604 104900 225616
rect 95200 225576 104900 225604
rect 95200 225564 95206 225576
rect 104894 225564 104900 225576
rect 104952 225564 104958 225616
rect 113082 225564 113088 225616
rect 113140 225604 113146 225616
rect 238846 225604 238852 225616
rect 113140 225576 238852 225604
rect 113140 225564 113146 225576
rect 238846 225564 238852 225576
rect 238904 225564 238910 225616
rect 173250 224952 173256 225004
rect 173308 224992 173314 225004
rect 173802 224992 173808 225004
rect 173308 224964 173808 224992
rect 173308 224952 173314 224964
rect 173802 224952 173808 224964
rect 173860 224952 173866 225004
rect 174630 224884 174636 224936
rect 174688 224924 174694 224936
rect 240778 224924 240784 224936
rect 174688 224896 240784 224924
rect 174688 224884 174694 224896
rect 240778 224884 240784 224896
rect 240836 224884 240842 224936
rect 252462 224884 252468 224936
rect 252520 224924 252526 224936
rect 258258 224924 258264 224936
rect 252520 224896 258264 224924
rect 252520 224884 252526 224896
rect 258258 224884 258264 224896
rect 258316 224884 258322 224936
rect 264882 224408 264888 224460
rect 264940 224448 264946 224460
rect 267918 224448 267924 224460
rect 264940 224420 267924 224448
rect 264940 224408 264946 224420
rect 267918 224408 267924 224420
rect 267976 224408 267982 224460
rect 138658 224272 138664 224324
rect 138716 224312 138722 224324
rect 227806 224312 227812 224324
rect 138716 224284 227812 224312
rect 138716 224272 138722 224284
rect 227806 224272 227812 224284
rect 227864 224312 227870 224324
rect 227864 224284 229094 224312
rect 227864 224272 227870 224284
rect 63034 224204 63040 224256
rect 63092 224244 63098 224256
rect 174722 224244 174728 224256
rect 63092 224216 174728 224244
rect 63092 224204 63098 224216
rect 174722 224204 174728 224216
rect 174780 224204 174786 224256
rect 229066 224244 229094 224284
rect 256878 224244 256884 224256
rect 229066 224216 256884 224244
rect 256878 224204 256884 224216
rect 256936 224204 256942 224256
rect 166350 223524 166356 223576
rect 166408 223564 166414 223576
rect 266354 223564 266360 223576
rect 166408 223536 266360 223564
rect 166408 223524 166414 223536
rect 266354 223524 266360 223536
rect 266412 223524 266418 223576
rect 112530 222844 112536 222896
rect 112588 222884 112594 222896
rect 117314 222884 117320 222896
rect 112588 222856 117320 222884
rect 112588 222844 112594 222856
rect 117314 222844 117320 222856
rect 117372 222844 117378 222896
rect 216030 222844 216036 222896
rect 216088 222884 216094 222896
rect 254026 222884 254032 222896
rect 216088 222856 254032 222884
rect 216088 222844 216094 222856
rect 254026 222844 254032 222856
rect 254084 222844 254090 222896
rect 187050 221552 187056 221604
rect 187108 221592 187114 221604
rect 224218 221592 224224 221604
rect 187108 221564 224224 221592
rect 187108 221552 187114 221564
rect 224218 221552 224224 221564
rect 224276 221552 224282 221604
rect 202138 221484 202144 221536
rect 202196 221524 202202 221536
rect 252738 221524 252744 221536
rect 202196 221496 252744 221524
rect 202196 221484 202202 221496
rect 252738 221484 252744 221496
rect 252796 221484 252802 221536
rect 47946 221416 47952 221468
rect 48004 221456 48010 221468
rect 202230 221456 202236 221468
rect 48004 221428 202236 221456
rect 48004 221416 48010 221428
rect 202230 221416 202236 221428
rect 202288 221416 202294 221468
rect 244274 221416 244280 221468
rect 244332 221456 244338 221468
rect 254578 221456 254584 221468
rect 244332 221428 254584 221456
rect 244332 221416 244338 221428
rect 254578 221416 254584 221428
rect 254636 221416 254642 221468
rect 67358 220736 67364 220788
rect 67416 220776 67422 220788
rect 273438 220776 273444 220788
rect 67416 220748 273444 220776
rect 67416 220736 67422 220748
rect 273438 220736 273444 220748
rect 273496 220736 273502 220788
rect 169202 220668 169208 220720
rect 169260 220708 169266 220720
rect 169662 220708 169668 220720
rect 169260 220680 169668 220708
rect 169260 220668 169266 220680
rect 169662 220668 169668 220680
rect 169720 220708 169726 220720
rect 243538 220708 243544 220720
rect 169720 220680 243544 220708
rect 169720 220668 169726 220680
rect 243538 220668 243544 220680
rect 243596 220668 243602 220720
rect 82722 220056 82728 220108
rect 82780 220096 82786 220108
rect 112438 220096 112444 220108
rect 82780 220068 112444 220096
rect 82780 220056 82786 220068
rect 112438 220056 112444 220068
rect 112496 220056 112502 220108
rect 224218 219376 224224 219428
rect 224276 219416 224282 219428
rect 265250 219416 265256 219428
rect 224276 219388 265256 219416
rect 224276 219376 224282 219388
rect 265250 219376 265256 219388
rect 265308 219376 265314 219428
rect 84010 218696 84016 218748
rect 84068 218736 84074 218748
rect 113266 218736 113272 218748
rect 84068 218708 113272 218736
rect 84068 218696 84074 218708
rect 113266 218696 113272 218708
rect 113324 218696 113330 218748
rect 149790 218696 149796 218748
rect 149848 218736 149854 218748
rect 230382 218736 230388 218748
rect 149848 218708 230388 218736
rect 149848 218696 149854 218708
rect 230382 218696 230388 218708
rect 230440 218696 230446 218748
rect 113266 218016 113272 218068
rect 113324 218056 113330 218068
rect 186314 218056 186320 218068
rect 113324 218028 186320 218056
rect 113324 218016 113330 218028
rect 186314 218016 186320 218028
rect 186372 218016 186378 218068
rect 229738 217948 229744 218000
rect 229796 217988 229802 218000
rect 230382 217988 230388 218000
rect 229796 217960 230388 217988
rect 229796 217948 229802 217960
rect 230382 217948 230388 217960
rect 230440 217988 230446 218000
rect 251818 217988 251824 218000
rect 230440 217960 251824 217988
rect 230440 217948 230446 217960
rect 251818 217948 251824 217960
rect 251876 217948 251882 218000
rect 161382 217268 161388 217320
rect 161440 217308 161446 217320
rect 266630 217308 266636 217320
rect 161440 217280 266636 217308
rect 161440 217268 161446 217280
rect 266630 217268 266636 217280
rect 266688 217268 266694 217320
rect 49602 216588 49608 216640
rect 49660 216628 49666 216640
rect 161382 216628 161388 216640
rect 49660 216600 161388 216628
rect 49660 216588 49666 216600
rect 161382 216588 161388 216600
rect 161440 216628 161446 216640
rect 161566 216628 161572 216640
rect 161440 216600 161572 216628
rect 161440 216588 161446 216600
rect 161566 216588 161572 216600
rect 161624 216588 161630 216640
rect 198090 215976 198096 216028
rect 198148 216016 198154 216028
rect 251174 216016 251180 216028
rect 198148 215988 251180 216016
rect 198148 215976 198154 215988
rect 251174 215976 251180 215988
rect 251232 215976 251238 216028
rect 160738 215908 160744 215960
rect 160796 215948 160802 215960
rect 220814 215948 220820 215960
rect 160796 215920 220820 215948
rect 160796 215908 160802 215920
rect 220814 215908 220820 215920
rect 220872 215948 220878 215960
rect 258166 215948 258172 215960
rect 220872 215920 258172 215948
rect 220872 215908 220878 215920
rect 258166 215908 258172 215920
rect 258224 215908 258230 215960
rect 89714 215228 89720 215280
rect 89772 215268 89778 215280
rect 117406 215268 117412 215280
rect 89772 215240 117412 215268
rect 89772 215228 89778 215240
rect 117406 215228 117412 215240
rect 117464 215228 117470 215280
rect 145650 215228 145656 215280
rect 145708 215268 145714 215280
rect 251082 215268 251088 215280
rect 145708 215240 251088 215268
rect 145708 215228 145714 215240
rect 251082 215228 251088 215240
rect 251140 215268 251146 215280
rect 253934 215268 253940 215280
rect 251140 215240 253940 215268
rect 251140 215228 251146 215240
rect 253934 215228 253940 215240
rect 253992 215228 253998 215280
rect 117406 214752 117412 214804
rect 117464 214792 117470 214804
rect 120166 214792 120172 214804
rect 117464 214764 120172 214792
rect 117464 214752 117470 214764
rect 120166 214752 120172 214764
rect 120224 214752 120230 214804
rect 174722 214548 174728 214600
rect 174780 214588 174786 214600
rect 178678 214588 178684 214600
rect 174780 214560 178684 214588
rect 174780 214548 174786 214560
rect 178678 214548 178684 214560
rect 178736 214548 178742 214600
rect 251818 214548 251824 214600
rect 251876 214588 251882 214600
rect 266538 214588 266544 214600
rect 251876 214560 266544 214588
rect 251876 214548 251882 214560
rect 266538 214548 266544 214560
rect 266596 214548 266602 214600
rect 98638 213868 98644 213920
rect 98696 213908 98702 213920
rect 104158 213908 104164 213920
rect 98696 213880 104164 213908
rect 98696 213868 98702 213880
rect 104158 213868 104164 213880
rect 104216 213908 104222 213920
rect 262214 213908 262220 213920
rect 104216 213880 262220 213908
rect 104216 213868 104222 213880
rect 262214 213868 262220 213880
rect 262272 213868 262278 213920
rect 250438 213188 250444 213240
rect 250496 213228 250502 213240
rect 274726 213228 274732 213240
rect 250496 213200 274732 213228
rect 250496 213188 250502 213200
rect 274726 213188 274732 213200
rect 274784 213188 274790 213240
rect 97258 211760 97264 211812
rect 97316 211800 97322 211812
rect 114554 211800 114560 211812
rect 97316 211772 114560 211800
rect 97316 211760 97322 211772
rect 114554 211760 114560 211772
rect 114612 211760 114618 211812
rect 202230 211760 202236 211812
rect 202288 211800 202294 211812
rect 249702 211800 249708 211812
rect 202288 211772 249708 211800
rect 202288 211760 202294 211772
rect 249702 211760 249708 211772
rect 249760 211760 249766 211812
rect 114554 211148 114560 211200
rect 114612 211188 114618 211200
rect 262398 211188 262404 211200
rect 114612 211160 262404 211188
rect 114612 211148 114618 211160
rect 262398 211148 262404 211160
rect 262456 211148 262462 211200
rect 73062 211080 73068 211132
rect 73120 211120 73126 211132
rect 249794 211120 249800 211132
rect 73120 211092 249800 211120
rect 73120 211080 73126 211092
rect 249794 211080 249800 211092
rect 249852 211120 249858 211132
rect 250990 211120 250996 211132
rect 249852 211092 250996 211120
rect 249852 211080 249858 211092
rect 250990 211080 250996 211092
rect 251048 211080 251054 211132
rect 263594 211120 263600 211132
rect 258046 211092 263600 211120
rect 186314 211012 186320 211064
rect 186372 211052 186378 211064
rect 258046 211052 258074 211092
rect 263594 211080 263600 211092
rect 263652 211120 263658 211132
rect 264054 211120 264060 211132
rect 263652 211092 264060 211120
rect 263652 211080 263658 211092
rect 264054 211080 264060 211092
rect 264112 211080 264118 211132
rect 186372 211024 258074 211052
rect 186372 211012 186378 211024
rect 151262 209720 151268 209772
rect 151320 209760 151326 209772
rect 247034 209760 247040 209772
rect 151320 209732 247040 209760
rect 151320 209720 151326 209732
rect 247034 209720 247040 209732
rect 247092 209760 247098 209772
rect 247770 209760 247776 209772
rect 247092 209732 247776 209760
rect 247092 209720 247098 209732
rect 247770 209720 247776 209732
rect 247828 209720 247834 209772
rect 191834 209652 191840 209704
rect 191892 209692 191898 209704
rect 255958 209692 255964 209704
rect 191892 209664 255964 209692
rect 191892 209652 191898 209664
rect 255958 209652 255964 209664
rect 256016 209652 256022 209704
rect 33042 209040 33048 209092
rect 33100 209080 33106 209092
rect 184290 209080 184296 209092
rect 33100 209052 184296 209080
rect 33100 209040 33106 209052
rect 184290 209040 184296 209052
rect 184348 209040 184354 209092
rect 44082 207612 44088 207664
rect 44140 207652 44146 207664
rect 185670 207652 185676 207664
rect 44140 207624 185676 207652
rect 44140 207612 44146 207624
rect 185670 207612 185676 207624
rect 185728 207612 185734 207664
rect 246206 207612 246212 207664
rect 246264 207652 246270 207664
rect 251818 207652 251824 207664
rect 246264 207624 251824 207652
rect 246264 207612 246270 207624
rect 251818 207612 251824 207624
rect 251876 207612 251882 207664
rect 255958 207612 255964 207664
rect 256016 207652 256022 207664
rect 276198 207652 276204 207664
rect 256016 207624 276204 207652
rect 256016 207612 256022 207624
rect 276198 207612 276204 207624
rect 276256 207612 276262 207664
rect 94682 207000 94688 207052
rect 94740 207040 94746 207052
rect 245746 207040 245752 207052
rect 94740 207012 245752 207040
rect 94740 207000 94746 207012
rect 245746 207000 245752 207012
rect 245804 207040 245810 207052
rect 246206 207040 246212 207052
rect 245804 207012 246212 207040
rect 245804 207000 245810 207012
rect 246206 207000 246212 207012
rect 246264 207000 246270 207052
rect 135070 206932 135076 206984
rect 135128 206972 135134 206984
rect 270678 206972 270684 206984
rect 135128 206944 270684 206972
rect 135128 206932 135134 206944
rect 270678 206932 270684 206944
rect 270736 206932 270742 206984
rect 93118 206252 93124 206304
rect 93176 206292 93182 206304
rect 103698 206292 103704 206304
rect 93176 206264 103704 206292
rect 93176 206252 93182 206264
rect 103698 206252 103704 206264
rect 103756 206292 103762 206304
rect 134150 206292 134156 206304
rect 103756 206264 134156 206292
rect 103756 206252 103762 206264
rect 134150 206252 134156 206264
rect 134208 206292 134214 206304
rect 135070 206292 135076 206304
rect 134208 206264 135076 206292
rect 134208 206252 134214 206264
rect 135070 206252 135076 206264
rect 135128 206252 135134 206304
rect 193122 206252 193128 206304
rect 193180 206292 193186 206304
rect 226518 206292 226524 206304
rect 193180 206264 226524 206292
rect 193180 206252 193186 206264
rect 226518 206252 226524 206264
rect 226576 206252 226582 206304
rect 88242 204960 88248 205012
rect 88300 205000 88306 205012
rect 104894 205000 104900 205012
rect 88300 204972 104900 205000
rect 88300 204960 88306 204972
rect 104894 204960 104900 204972
rect 104952 205000 104958 205012
rect 106090 205000 106096 205012
rect 104952 204972 106096 205000
rect 104952 204960 104958 204972
rect 106090 204960 106096 204972
rect 106148 204960 106154 205012
rect 96614 204892 96620 204944
rect 96672 204932 96678 204944
rect 125594 204932 125600 204944
rect 96672 204904 125600 204932
rect 96672 204892 96678 204904
rect 125594 204892 125600 204904
rect 125652 204932 125658 204944
rect 133138 204932 133144 204944
rect 125652 204904 133144 204932
rect 125652 204892 125658 204904
rect 133138 204892 133144 204904
rect 133196 204932 133202 204944
rect 242894 204932 242900 204944
rect 133196 204904 242900 204932
rect 133196 204892 133202 204904
rect 242894 204892 242900 204904
rect 242952 204932 242958 204944
rect 281626 204932 281632 204944
rect 242952 204904 281632 204932
rect 242952 204892 242958 204904
rect 281626 204892 281632 204904
rect 281684 204892 281690 204944
rect 106090 204280 106096 204332
rect 106148 204320 106154 204332
rect 258074 204320 258080 204332
rect 106148 204292 258080 204320
rect 106148 204280 106154 204292
rect 258074 204280 258080 204292
rect 258132 204280 258138 204332
rect 155402 204212 155408 204264
rect 155460 204252 155466 204264
rect 259638 204252 259644 204264
rect 155460 204224 259644 204252
rect 155460 204212 155466 204224
rect 259638 204212 259644 204224
rect 259696 204212 259702 204264
rect 46842 203532 46848 203584
rect 46900 203572 46906 203584
rect 67818 203572 67824 203584
rect 46900 203544 67824 203572
rect 46900 203532 46906 203544
rect 67818 203532 67824 203544
rect 67876 203532 67882 203584
rect 214558 203532 214564 203584
rect 214616 203572 214622 203584
rect 253934 203572 253940 203584
rect 214616 203544 253940 203572
rect 214616 203532 214622 203544
rect 253934 203532 253940 203544
rect 253992 203532 253998 203584
rect 152550 202784 152556 202836
rect 152608 202824 152614 202836
rect 155310 202824 155316 202836
rect 152608 202796 155316 202824
rect 152608 202784 152614 202796
rect 155310 202784 155316 202796
rect 155368 202784 155374 202836
rect 180150 202784 180156 202836
rect 180208 202824 180214 202836
rect 180702 202824 180708 202836
rect 180208 202796 180708 202824
rect 180208 202784 180214 202796
rect 180702 202784 180708 202796
rect 180760 202824 180766 202836
rect 244918 202824 244924 202836
rect 180760 202796 244924 202824
rect 180760 202784 180766 202796
rect 244918 202784 244924 202796
rect 244976 202784 244982 202836
rect 3326 202172 3332 202224
rect 3384 202212 3390 202224
rect 98086 202212 98092 202224
rect 3384 202184 98092 202212
rect 3384 202172 3390 202184
rect 98086 202172 98092 202184
rect 98144 202172 98150 202224
rect 108942 202172 108948 202224
rect 109000 202212 109006 202224
rect 118694 202212 118700 202224
rect 109000 202184 118700 202212
rect 109000 202172 109006 202184
rect 118694 202172 118700 202184
rect 118752 202172 118758 202224
rect 138658 202172 138664 202224
rect 138716 202212 138722 202224
rect 148410 202212 148416 202224
rect 138716 202184 148416 202212
rect 138716 202172 138722 202184
rect 148410 202172 148416 202184
rect 148468 202172 148474 202224
rect 37090 202104 37096 202156
rect 37148 202144 37154 202156
rect 188522 202144 188528 202156
rect 37148 202116 188528 202144
rect 37148 202104 37154 202116
rect 188522 202104 188528 202116
rect 188580 202104 188586 202156
rect 253198 202104 253204 202156
rect 253256 202144 253262 202156
rect 270678 202144 270684 202156
rect 253256 202116 270684 202144
rect 253256 202104 253262 202116
rect 270678 202104 270684 202116
rect 270736 202104 270742 202156
rect 126330 201628 126336 201680
rect 126388 201668 126394 201680
rect 134610 201668 134616 201680
rect 126388 201640 134616 201668
rect 126388 201628 126394 201640
rect 134610 201628 134616 201640
rect 134668 201628 134674 201680
rect 171870 201424 171876 201476
rect 171928 201464 171934 201476
rect 172330 201464 172336 201476
rect 171928 201436 172336 201464
rect 171928 201424 171934 201436
rect 172330 201424 172336 201436
rect 172388 201464 172394 201476
rect 277486 201464 277492 201476
rect 172388 201436 277492 201464
rect 172388 201424 172394 201436
rect 277486 201424 277492 201436
rect 277544 201424 277550 201476
rect 133230 201356 133236 201408
rect 133288 201396 133294 201408
rect 231854 201396 231860 201408
rect 133288 201368 231860 201396
rect 133288 201356 133294 201368
rect 231854 201356 231860 201368
rect 231912 201396 231918 201408
rect 233142 201396 233148 201408
rect 231912 201368 233148 201396
rect 231912 201356 231918 201368
rect 233142 201356 233148 201368
rect 233200 201356 233206 201408
rect 75270 200744 75276 200796
rect 75328 200784 75334 200796
rect 107654 200784 107660 200796
rect 75328 200756 107660 200784
rect 75328 200744 75334 200756
rect 107654 200744 107660 200756
rect 107712 200744 107718 200796
rect 112622 200744 112628 200796
rect 112680 200784 112686 200796
rect 132586 200784 132592 200796
rect 112680 200756 132592 200784
rect 112680 200744 112686 200756
rect 132586 200744 132592 200756
rect 132644 200744 132650 200796
rect 149698 200064 149704 200116
rect 149756 200104 149762 200116
rect 252646 200104 252652 200116
rect 149756 200076 252652 200104
rect 149756 200064 149762 200076
rect 252646 200064 252652 200076
rect 252704 200064 252710 200116
rect 170950 199996 170956 200048
rect 171008 200036 171014 200048
rect 269298 200036 269304 200048
rect 171008 200008 269304 200036
rect 171008 199996 171014 200008
rect 269298 199996 269304 200008
rect 269356 199996 269362 200048
rect 45370 199384 45376 199436
rect 45428 199424 45434 199436
rect 76650 199424 76656 199436
rect 45428 199396 76656 199424
rect 45428 199384 45434 199396
rect 76650 199384 76656 199396
rect 76708 199384 76714 199436
rect 86218 199384 86224 199436
rect 86276 199424 86282 199436
rect 103606 199424 103612 199436
rect 86276 199396 103612 199424
rect 86276 199384 86282 199396
rect 103606 199384 103612 199396
rect 103664 199384 103670 199436
rect 106182 199384 106188 199436
rect 106240 199424 106246 199436
rect 122834 199424 122840 199436
rect 106240 199396 122840 199424
rect 106240 199384 106246 199396
rect 122834 199384 122840 199396
rect 122892 199384 122898 199436
rect 147030 198704 147036 198756
rect 147088 198744 147094 198756
rect 153838 198744 153844 198756
rect 147088 198716 153844 198744
rect 147088 198704 147094 198716
rect 153838 198704 153844 198716
rect 153896 198704 153902 198756
rect 38562 197956 38568 198008
rect 38620 197996 38626 198008
rect 224954 197996 224960 198008
rect 38620 197968 224960 197996
rect 38620 197956 38626 197968
rect 224954 197956 224960 197968
rect 225012 197956 225018 198008
rect 256050 197956 256056 198008
rect 256108 197996 256114 198008
rect 276014 197996 276020 198008
rect 256108 197968 276020 197996
rect 256108 197956 256114 197968
rect 276014 197956 276020 197968
rect 276072 197956 276078 198008
rect 217410 196596 217416 196648
rect 217468 196636 217474 196648
rect 242158 196636 242164 196648
rect 217468 196608 242164 196636
rect 217468 196596 217474 196608
rect 242158 196596 242164 196608
rect 242216 196596 242222 196648
rect 249058 196596 249064 196648
rect 249116 196636 249122 196648
rect 284386 196636 284392 196648
rect 249116 196608 284392 196636
rect 249116 196596 249122 196608
rect 284386 196596 284392 196608
rect 284444 196596 284450 196648
rect 193306 195304 193312 195356
rect 193364 195344 193370 195356
rect 224954 195344 224960 195356
rect 193364 195316 224960 195344
rect 193364 195304 193370 195316
rect 224954 195304 224960 195316
rect 225012 195304 225018 195356
rect 79962 195236 79968 195288
rect 80020 195276 80026 195288
rect 110414 195276 110420 195288
rect 80020 195248 110420 195276
rect 80020 195236 80026 195248
rect 110414 195236 110420 195248
rect 110472 195236 110478 195288
rect 222930 195236 222936 195288
rect 222988 195276 222994 195288
rect 271966 195276 271972 195288
rect 222988 195248 271972 195276
rect 222988 195236 222994 195248
rect 271966 195236 271972 195248
rect 272024 195236 272030 195288
rect 246298 193808 246304 193860
rect 246356 193848 246362 193860
rect 281534 193848 281540 193860
rect 246356 193820 281540 193848
rect 246356 193808 246362 193820
rect 281534 193808 281540 193820
rect 281592 193808 281598 193860
rect 84102 192516 84108 192568
rect 84160 192556 84166 192568
rect 107010 192556 107016 192568
rect 84160 192528 107016 192556
rect 84160 192516 84166 192528
rect 107010 192516 107016 192528
rect 107068 192516 107074 192568
rect 2682 192448 2688 192500
rect 2740 192488 2746 192500
rect 152642 192488 152648 192500
rect 2740 192460 152648 192488
rect 2740 192448 2746 192460
rect 152642 192448 152648 192460
rect 152700 192448 152706 192500
rect 166350 192448 166356 192500
rect 166408 192488 166414 192500
rect 217318 192488 217324 192500
rect 166408 192460 217324 192488
rect 166408 192448 166414 192460
rect 217318 192448 217324 192460
rect 217376 192448 217382 192500
rect 240778 192448 240784 192500
rect 240836 192488 240842 192500
rect 580166 192488 580172 192500
rect 240836 192460 580172 192488
rect 240836 192448 240842 192460
rect 580166 192448 580172 192460
rect 580224 192448 580230 192500
rect 178678 191768 178684 191820
rect 178736 191808 178742 191820
rect 278038 191808 278044 191820
rect 178736 191780 278044 191808
rect 178736 191768 178742 191780
rect 278038 191768 278044 191780
rect 278096 191768 278102 191820
rect 187602 189728 187608 189780
rect 187660 189768 187666 189780
rect 252922 189768 252928 189780
rect 187660 189740 252928 189768
rect 187660 189728 187666 189740
rect 252922 189728 252928 189740
rect 252980 189728 252986 189780
rect 3510 188980 3516 189032
rect 3568 189020 3574 189032
rect 18598 189020 18604 189032
rect 3568 188992 18604 189020
rect 3568 188980 3574 188992
rect 18598 188980 18604 188992
rect 18656 188980 18662 189032
rect 195882 188300 195888 188352
rect 195940 188340 195946 188352
rect 226978 188340 226984 188352
rect 195940 188312 226984 188340
rect 195940 188300 195946 188312
rect 226978 188300 226984 188312
rect 227036 188300 227042 188352
rect 254578 188300 254584 188352
rect 254636 188340 254642 188352
rect 270586 188340 270592 188352
rect 254636 188312 270592 188340
rect 254636 188300 254642 188312
rect 270586 188300 270592 188312
rect 270644 188300 270650 188352
rect 27522 186940 27528 186992
rect 27580 186980 27586 186992
rect 151170 186980 151176 186992
rect 27580 186952 151176 186980
rect 27580 186940 27586 186952
rect 151170 186940 151176 186952
rect 151228 186940 151234 186992
rect 242158 186940 242164 186992
rect 242216 186980 242222 186992
rect 260926 186980 260932 186992
rect 242216 186952 260932 186980
rect 242216 186940 242222 186952
rect 260926 186940 260932 186952
rect 260984 186940 260990 186992
rect 6822 185580 6828 185632
rect 6880 185620 6886 185632
rect 147122 185620 147128 185632
rect 6880 185592 147128 185620
rect 6880 185580 6886 185592
rect 147122 185580 147128 185592
rect 147180 185580 147186 185632
rect 197998 185580 198004 185632
rect 198056 185620 198062 185632
rect 226426 185620 226432 185632
rect 198056 185592 226432 185620
rect 198056 185580 198062 185592
rect 226426 185580 226432 185592
rect 226484 185580 226490 185632
rect 232590 184152 232596 184204
rect 232648 184192 232654 184204
rect 252646 184192 252652 184204
rect 232648 184164 252652 184192
rect 232648 184152 232654 184164
rect 252646 184152 252652 184164
rect 252704 184152 252710 184204
rect 10962 182792 10968 182844
rect 11020 182832 11026 182844
rect 188338 182832 188344 182844
rect 11020 182804 188344 182832
rect 11020 182792 11026 182804
rect 188338 182792 188344 182804
rect 188396 182792 188402 182844
rect 192478 182792 192484 182844
rect 192536 182832 192542 182844
rect 220170 182832 220176 182844
rect 192536 182804 220176 182832
rect 192536 182792 192542 182804
rect 220170 182792 220176 182804
rect 220228 182792 220234 182844
rect 93118 180820 93124 180872
rect 93176 180860 93182 180872
rect 93762 180860 93768 180872
rect 93176 180832 93768 180860
rect 93176 180820 93182 180832
rect 93762 180820 93768 180832
rect 93820 180860 93826 180872
rect 218698 180860 218704 180872
rect 93820 180832 218704 180860
rect 93820 180820 93826 180832
rect 218698 180820 218704 180832
rect 218756 180820 218762 180872
rect 82078 180072 82084 180124
rect 82136 180112 82142 180124
rect 109126 180112 109132 180124
rect 82136 180084 109132 180112
rect 82136 180072 82142 180084
rect 109126 180072 109132 180084
rect 109184 180072 109190 180124
rect 195238 180072 195244 180124
rect 195296 180112 195302 180124
rect 226610 180112 226616 180124
rect 195296 180084 226616 180112
rect 195296 180072 195302 180084
rect 226610 180072 226616 180084
rect 226668 180072 226674 180124
rect 135898 179392 135904 179444
rect 135956 179432 135962 179444
rect 218790 179432 218796 179444
rect 135956 179404 218796 179432
rect 135956 179392 135962 179404
rect 218790 179392 218796 179404
rect 218848 179392 218854 179444
rect 252462 178644 252468 178696
rect 252520 178684 252526 178696
rect 580166 178684 580172 178696
rect 252520 178656 580172 178684
rect 252520 178644 252526 178656
rect 580166 178644 580172 178656
rect 580224 178644 580230 178696
rect 57606 178100 57612 178152
rect 57664 178140 57670 178152
rect 156690 178140 156696 178152
rect 57664 178112 156696 178140
rect 57664 178100 57670 178112
rect 156690 178100 156696 178112
rect 156748 178100 156754 178152
rect 90358 178032 90364 178084
rect 90416 178072 90422 178084
rect 91002 178072 91008 178084
rect 90416 178044 91008 178072
rect 90416 178032 90422 178044
rect 91002 178032 91008 178044
rect 91060 178072 91066 178084
rect 217318 178072 217324 178084
rect 91060 178044 217324 178072
rect 91060 178032 91066 178044
rect 217318 178032 217324 178044
rect 217376 178032 217382 178084
rect 251818 178032 251824 178084
rect 251876 178072 251882 178084
rect 252462 178072 252468 178084
rect 251876 178044 252468 178072
rect 251876 178032 251882 178044
rect 252462 178032 252468 178044
rect 252520 178032 252526 178084
rect 82814 177284 82820 177336
rect 82872 177324 82878 177336
rect 110506 177324 110512 177336
rect 82872 177296 110512 177324
rect 82872 177284 82878 177296
rect 110506 177284 110512 177296
rect 110564 177324 110570 177336
rect 214006 177324 214012 177336
rect 110564 177296 214012 177324
rect 110564 177284 110570 177296
rect 214006 177284 214012 177296
rect 214064 177284 214070 177336
rect 252462 177284 252468 177336
rect 252520 177324 252526 177336
rect 262306 177324 262312 177336
rect 252520 177296 262312 177324
rect 252520 177284 252526 177296
rect 262306 177284 262312 177296
rect 262364 177284 262370 177336
rect 216122 176672 216128 176724
rect 216180 176712 216186 176724
rect 251174 176712 251180 176724
rect 216180 176684 251180 176712
rect 216180 176672 216186 176684
rect 251174 176672 251180 176684
rect 251232 176712 251238 176724
rect 252462 176712 252468 176724
rect 251232 176684 252468 176712
rect 251232 176672 251238 176684
rect 252462 176672 252468 176684
rect 252520 176672 252526 176724
rect 195238 175312 195244 175364
rect 195296 175352 195302 175364
rect 195882 175352 195888 175364
rect 195296 175324 195888 175352
rect 195296 175312 195302 175324
rect 195882 175312 195888 175324
rect 195940 175352 195946 175364
rect 295978 175352 295984 175364
rect 195940 175324 295984 175352
rect 195940 175312 195946 175324
rect 295978 175312 295984 175324
rect 296036 175312 296042 175364
rect 78858 175244 78864 175296
rect 78916 175284 78922 175296
rect 207106 175284 207112 175296
rect 78916 175256 207112 175284
rect 78916 175244 78922 175256
rect 207106 175244 207112 175256
rect 207164 175244 207170 175296
rect 202874 174496 202880 174548
rect 202932 174536 202938 174548
rect 226702 174536 226708 174548
rect 202932 174508 226708 174536
rect 202932 174496 202938 174508
rect 226702 174496 226708 174508
rect 226760 174496 226766 174548
rect 82906 173884 82912 173936
rect 82964 173924 82970 173936
rect 211798 173924 211804 173936
rect 82964 173896 211804 173924
rect 82964 173884 82970 173896
rect 211798 173884 211804 173896
rect 211856 173884 211862 173936
rect 75914 173408 75920 173460
rect 75972 173448 75978 173460
rect 76742 173448 76748 173460
rect 75972 173420 76748 173448
rect 75972 173408 75978 173420
rect 76742 173408 76748 173420
rect 76800 173408 76806 173460
rect 76742 173136 76748 173188
rect 76800 173176 76806 173188
rect 202874 173176 202880 173188
rect 76800 173148 202880 173176
rect 76800 173136 76806 173148
rect 202874 173136 202880 173148
rect 202932 173136 202938 173188
rect 91738 172524 91744 172576
rect 91796 172564 91802 172576
rect 220814 172564 220820 172576
rect 91796 172536 220820 172564
rect 91796 172524 91802 172536
rect 220814 172524 220820 172536
rect 220872 172524 220878 172576
rect 195974 172320 195980 172372
rect 196032 172360 196038 172372
rect 196802 172360 196808 172372
rect 196032 172332 196808 172360
rect 196032 172320 196038 172332
rect 196802 172320 196808 172332
rect 196860 172320 196866 172372
rect 244918 171776 244924 171828
rect 244976 171816 244982 171828
rect 246114 171816 246120 171828
rect 244976 171788 246120 171816
rect 244976 171776 244982 171788
rect 246114 171776 246120 171788
rect 246172 171776 246178 171828
rect 177850 171164 177856 171216
rect 177908 171204 177914 171216
rect 188338 171204 188344 171216
rect 177908 171176 188344 171204
rect 177908 171164 177914 171176
rect 188338 171164 188344 171176
rect 188396 171164 188402 171216
rect 81434 171096 81440 171148
rect 81492 171136 81498 171148
rect 196802 171136 196808 171148
rect 81492 171108 196808 171136
rect 81492 171096 81498 171108
rect 196802 171096 196808 171108
rect 196860 171096 196866 171148
rect 246390 171096 246396 171148
rect 246448 171136 246454 171148
rect 249426 171136 249432 171148
rect 246448 171108 249432 171136
rect 246448 171096 246454 171108
rect 249426 171096 249432 171108
rect 249484 171096 249490 171148
rect 86218 170416 86224 170468
rect 86276 170456 86282 170468
rect 177850 170456 177856 170468
rect 86276 170428 177856 170456
rect 86276 170416 86282 170428
rect 177850 170416 177856 170428
rect 177908 170416 177914 170468
rect 196710 170416 196716 170468
rect 196768 170456 196774 170468
rect 273254 170456 273260 170468
rect 196768 170428 273260 170456
rect 196768 170416 196774 170428
rect 273254 170416 273260 170428
rect 273312 170416 273318 170468
rect 77938 170348 77944 170400
rect 77996 170388 78002 170400
rect 204898 170388 204904 170400
rect 77996 170360 204904 170388
rect 77996 170348 78002 170360
rect 204898 170348 204904 170360
rect 204956 170348 204962 170400
rect 205634 170348 205640 170400
rect 205692 170388 205698 170400
rect 217410 170388 217416 170400
rect 205692 170360 217416 170388
rect 205692 170348 205698 170360
rect 217410 170348 217416 170360
rect 217468 170348 217474 170400
rect 77386 169736 77392 169788
rect 77444 169776 77450 169788
rect 77938 169776 77944 169788
rect 77444 169748 77944 169776
rect 77444 169736 77450 169748
rect 77938 169736 77944 169748
rect 77996 169736 78002 169788
rect 123662 169668 123668 169720
rect 123720 169708 123726 169720
rect 224862 169708 224868 169720
rect 123720 169680 224868 169708
rect 123720 169668 123726 169680
rect 224862 169668 224868 169680
rect 224920 169668 224926 169720
rect 93854 168988 93860 169040
rect 93912 169028 93918 169040
rect 122926 169028 122932 169040
rect 93912 169000 122932 169028
rect 93912 168988 93918 169000
rect 122926 168988 122932 169000
rect 122984 169028 122990 169040
rect 123662 169028 123668 169040
rect 122984 169000 123668 169028
rect 122984 168988 122990 169000
rect 123662 168988 123668 169000
rect 123720 168988 123726 169040
rect 182910 168988 182916 169040
rect 182968 169028 182974 169040
rect 264974 169028 264980 169040
rect 182968 169000 264980 169028
rect 182968 168988 182974 169000
rect 264974 168988 264980 169000
rect 265032 168988 265038 169040
rect 224310 168376 224316 168428
rect 224368 168416 224374 168428
rect 224862 168416 224868 168428
rect 224368 168388 224868 168416
rect 224368 168376 224374 168388
rect 224862 168376 224868 168388
rect 224920 168376 224926 168428
rect 193030 167696 193036 167748
rect 193088 167736 193094 167748
rect 200114 167736 200120 167748
rect 193088 167708 200120 167736
rect 193088 167696 193094 167708
rect 200114 167696 200120 167708
rect 200172 167696 200178 167748
rect 53466 167628 53472 167680
rect 53524 167668 53530 167680
rect 210418 167668 210424 167680
rect 53524 167640 210424 167668
rect 53524 167628 53530 167640
rect 210418 167628 210424 167640
rect 210476 167628 210482 167680
rect 221458 167016 221464 167068
rect 221516 167056 221522 167068
rect 222102 167056 222108 167068
rect 221516 167028 222108 167056
rect 221516 167016 221522 167028
rect 222102 167016 222108 167028
rect 222160 167056 222166 167068
rect 285674 167056 285680 167068
rect 222160 167028 285680 167056
rect 222160 167016 222166 167028
rect 285674 167016 285680 167028
rect 285732 167016 285738 167068
rect 195054 166336 195060 166388
rect 195112 166376 195118 166388
rect 222102 166376 222108 166388
rect 195112 166348 222108 166376
rect 195112 166336 195118 166348
rect 222102 166336 222108 166348
rect 222160 166336 222166 166388
rect 217410 166268 217416 166320
rect 217468 166308 217474 166320
rect 259822 166308 259828 166320
rect 217468 166280 259828 166308
rect 217468 166268 217474 166280
rect 259822 166268 259828 166280
rect 259880 166268 259886 166320
rect 197354 166064 197360 166116
rect 197412 166104 197418 166116
rect 198090 166104 198096 166116
rect 197412 166076 198096 166104
rect 197412 166064 197418 166076
rect 198090 166064 198096 166076
rect 198148 166064 198154 166116
rect 86310 165656 86316 165708
rect 86368 165696 86374 165708
rect 197354 165696 197360 165708
rect 86368 165668 197360 165696
rect 86368 165656 86374 165668
rect 197354 165656 197360 165668
rect 197412 165656 197418 165708
rect 75270 165588 75276 165640
rect 75328 165628 75334 165640
rect 194594 165628 194600 165640
rect 75328 165600 194600 165628
rect 75328 165588 75334 165600
rect 194594 165588 194600 165600
rect 194652 165628 194658 165640
rect 195054 165628 195060 165640
rect 194652 165600 195060 165628
rect 194652 165588 194658 165600
rect 195054 165588 195060 165600
rect 195112 165588 195118 165640
rect 91002 164908 91008 164960
rect 91060 164948 91066 164960
rect 117314 164948 117320 164960
rect 91060 164920 117320 164948
rect 91060 164908 91066 164920
rect 117314 164908 117320 164920
rect 117372 164948 117378 164960
rect 220814 164948 220820 164960
rect 117372 164920 220820 164948
rect 117372 164908 117378 164920
rect 220814 164908 220820 164920
rect 220872 164908 220878 164960
rect 46658 164840 46664 164892
rect 46716 164880 46722 164892
rect 192478 164880 192484 164892
rect 46716 164852 192484 164880
rect 46716 164840 46722 164852
rect 192478 164840 192484 164852
rect 192536 164840 192542 164892
rect 198734 164840 198740 164892
rect 198792 164880 198798 164892
rect 259454 164880 259460 164892
rect 198792 164852 259460 164880
rect 198792 164840 198798 164852
rect 259454 164840 259460 164852
rect 259512 164840 259518 164892
rect 204162 163480 204168 163532
rect 204220 163520 204226 163532
rect 237466 163520 237472 163532
rect 204220 163492 237472 163520
rect 204220 163480 204226 163492
rect 237466 163480 237472 163492
rect 237524 163520 237530 163532
rect 306374 163520 306380 163532
rect 237524 163492 306380 163520
rect 237524 163480 237530 163492
rect 306374 163480 306380 163492
rect 306432 163480 306438 163532
rect 131758 162936 131764 162988
rect 131816 162976 131822 162988
rect 236086 162976 236092 162988
rect 131816 162948 236092 162976
rect 131816 162936 131822 162948
rect 236086 162936 236092 162948
rect 236144 162936 236150 162988
rect 3510 162868 3516 162920
rect 3568 162908 3574 162920
rect 8938 162908 8944 162920
rect 3568 162880 8944 162908
rect 3568 162868 3574 162880
rect 8938 162868 8944 162880
rect 8996 162868 9002 162920
rect 73062 162868 73068 162920
rect 73120 162908 73126 162920
rect 198734 162908 198740 162920
rect 73120 162880 198740 162908
rect 73120 162868 73126 162880
rect 198734 162868 198740 162880
rect 198792 162868 198798 162920
rect 97442 162800 97448 162852
rect 97500 162840 97506 162852
rect 97902 162840 97908 162852
rect 97500 162812 97908 162840
rect 97500 162800 97506 162812
rect 97902 162800 97908 162812
rect 97960 162800 97966 162852
rect 213914 162800 213920 162852
rect 213972 162840 213978 162852
rect 214558 162840 214564 162852
rect 213972 162812 214564 162840
rect 213972 162800 213978 162812
rect 214558 162800 214564 162812
rect 214616 162800 214622 162852
rect 245654 162800 245660 162852
rect 245712 162840 245718 162852
rect 246390 162840 246396 162852
rect 245712 162812 246396 162840
rect 245712 162800 245718 162812
rect 246390 162800 246396 162812
rect 246448 162800 246454 162852
rect 97442 162120 97448 162172
rect 97500 162160 97506 162172
rect 245654 162160 245660 162172
rect 97500 162132 245660 162160
rect 97500 162120 97506 162132
rect 245654 162120 245660 162132
rect 245712 162120 245718 162172
rect 180794 161440 180800 161492
rect 180852 161480 180858 161492
rect 181990 161480 181996 161492
rect 180852 161452 181996 161480
rect 180852 161440 180858 161452
rect 181990 161440 181996 161452
rect 182048 161480 182054 161492
rect 213270 161480 213276 161492
rect 182048 161452 213276 161480
rect 182048 161440 182054 161452
rect 213270 161440 213276 161452
rect 213328 161440 213334 161492
rect 213914 161440 213920 161492
rect 213972 161480 213978 161492
rect 582650 161480 582656 161492
rect 213972 161452 582656 161480
rect 213972 161440 213978 161452
rect 582650 161440 582656 161452
rect 582708 161440 582714 161492
rect 34330 160692 34336 160744
rect 34388 160732 34394 160744
rect 60734 160732 60740 160744
rect 34388 160704 60740 160732
rect 34388 160692 34394 160704
rect 60734 160692 60740 160704
rect 60792 160692 60798 160744
rect 105538 160148 105544 160200
rect 105596 160188 105602 160200
rect 230566 160188 230572 160200
rect 105596 160160 230572 160188
rect 105596 160148 105602 160160
rect 230566 160148 230572 160160
rect 230624 160148 230630 160200
rect 60734 160080 60740 160132
rect 60792 160120 60798 160132
rect 61746 160120 61752 160132
rect 60792 160092 61752 160120
rect 60792 160080 60798 160092
rect 61746 160080 61752 160092
rect 61804 160120 61810 160132
rect 189810 160120 189816 160132
rect 61804 160092 189816 160120
rect 61804 160080 61810 160092
rect 189810 160080 189816 160092
rect 189868 160080 189874 160132
rect 188338 159400 188344 159452
rect 188396 159440 188402 159452
rect 211154 159440 211160 159452
rect 188396 159412 211160 159440
rect 188396 159400 188402 159412
rect 211154 159400 211160 159412
rect 211212 159400 211218 159452
rect 87138 159332 87144 159384
rect 87196 159372 87202 159384
rect 180794 159372 180800 159384
rect 87196 159344 180800 159372
rect 87196 159332 87202 159344
rect 180794 159332 180800 159344
rect 180852 159332 180858 159384
rect 208578 159332 208584 159384
rect 208636 159372 208642 159384
rect 274634 159372 274640 159384
rect 208636 159344 274640 159372
rect 208636 159332 208642 159344
rect 274634 159332 274640 159344
rect 274692 159332 274698 159384
rect 83458 158720 83464 158772
rect 83516 158760 83522 158772
rect 196066 158760 196072 158772
rect 83516 158732 196072 158760
rect 83516 158720 83522 158732
rect 196066 158720 196072 158732
rect 196124 158720 196130 158772
rect 190362 157972 190368 158024
rect 190420 158012 190426 158024
rect 249702 158012 249708 158024
rect 190420 157984 249708 158012
rect 190420 157972 190426 157984
rect 249702 157972 249708 157984
rect 249760 158012 249766 158024
rect 580350 158012 580356 158024
rect 249760 157984 580356 158012
rect 249760 157972 249766 157984
rect 580350 157972 580356 157984
rect 580408 157972 580414 158024
rect 75178 157428 75184 157480
rect 75236 157468 75242 157480
rect 189902 157468 189908 157480
rect 75236 157440 189908 157468
rect 75236 157428 75242 157440
rect 189902 157428 189908 157440
rect 189960 157428 189966 157480
rect 90450 157360 90456 157412
rect 90508 157400 90514 157412
rect 208578 157400 208584 157412
rect 90508 157372 208584 157400
rect 90508 157360 90514 157372
rect 208578 157360 208584 157372
rect 208636 157360 208642 157412
rect 163590 156408 163596 156460
rect 163648 156448 163654 156460
rect 164142 156448 164148 156460
rect 163648 156420 164148 156448
rect 163648 156408 163654 156420
rect 164142 156408 164148 156420
rect 164200 156408 164206 156460
rect 56318 156000 56324 156052
rect 56376 156040 56382 156052
rect 160830 156040 160836 156052
rect 56376 156012 160836 156040
rect 56376 156000 56382 156012
rect 160830 156000 160836 156012
rect 160888 156000 160894 156052
rect 164142 156000 164148 156052
rect 164200 156040 164206 156052
rect 220078 156040 220084 156052
rect 164200 156012 220084 156040
rect 164200 156000 164206 156012
rect 220078 156000 220084 156012
rect 220136 156000 220142 156052
rect 222286 156000 222292 156052
rect 222344 156040 222350 156052
rect 260098 156040 260104 156052
rect 222344 156012 260104 156040
rect 222344 156000 222350 156012
rect 260098 156000 260104 156012
rect 260156 156000 260162 156052
rect 98730 155932 98736 155984
rect 98788 155972 98794 155984
rect 99282 155972 99288 155984
rect 98788 155944 99288 155972
rect 98788 155932 98794 155944
rect 99282 155932 99288 155944
rect 99340 155972 99346 155984
rect 225138 155972 225144 155984
rect 99340 155944 225144 155972
rect 99340 155932 99346 155944
rect 225138 155932 225144 155944
rect 225196 155932 225202 155984
rect 211246 155864 211252 155916
rect 211304 155904 211310 155916
rect 211798 155904 211804 155916
rect 211304 155876 211804 155904
rect 211304 155864 211310 155876
rect 211798 155864 211804 155876
rect 211856 155904 211862 155916
rect 288434 155904 288440 155916
rect 211856 155876 288440 155904
rect 211856 155864 211862 155876
rect 288434 155864 288440 155876
rect 288492 155904 288498 155916
rect 289722 155904 289728 155916
rect 288492 155876 289728 155904
rect 288492 155864 288498 155876
rect 289722 155864 289728 155876
rect 289780 155864 289786 155916
rect 177390 155184 177396 155236
rect 177448 155224 177454 155236
rect 205082 155224 205088 155236
rect 177448 155196 205088 155224
rect 177448 155184 177454 155196
rect 205082 155184 205088 155196
rect 205140 155184 205146 155236
rect 289722 155184 289728 155236
rect 289780 155224 289786 155236
rect 317414 155224 317420 155236
rect 289780 155196 317420 155224
rect 289780 155184 289786 155196
rect 317414 155184 317420 155196
rect 317472 155184 317478 155236
rect 60366 154572 60372 154624
rect 60424 154612 60430 154624
rect 178770 154612 178776 154624
rect 60424 154584 178776 154612
rect 60424 154572 60430 154584
rect 178770 154572 178776 154584
rect 178828 154572 178834 154624
rect 251266 154504 251272 154556
rect 251324 154544 251330 154556
rect 251818 154544 251824 154556
rect 251324 154516 251824 154544
rect 251324 154504 251330 154516
rect 251818 154504 251824 154516
rect 251876 154504 251882 154556
rect 39850 153824 39856 153876
rect 39908 153864 39914 153876
rect 158070 153864 158076 153876
rect 39908 153836 158076 153864
rect 39908 153824 39914 153836
rect 158070 153824 158076 153836
rect 158128 153824 158134 153876
rect 175826 153280 175832 153332
rect 175884 153320 175890 153332
rect 227898 153320 227904 153332
rect 175884 153292 227904 153320
rect 175884 153280 175890 153292
rect 227898 153280 227904 153292
rect 227956 153280 227962 153332
rect 155310 153212 155316 153264
rect 155368 153252 155374 153264
rect 251266 153252 251272 153264
rect 155368 153224 251272 153252
rect 155368 153212 155374 153224
rect 251266 153212 251272 153224
rect 251324 153212 251330 153264
rect 130470 152600 130476 152652
rect 130528 152640 130534 152652
rect 131022 152640 131028 152652
rect 130528 152612 131028 152640
rect 130528 152600 130534 152612
rect 131022 152600 131028 152612
rect 131080 152600 131086 152652
rect 86862 152532 86868 152584
rect 86920 152572 86926 152584
rect 102134 152572 102140 152584
rect 86920 152544 102140 152572
rect 86920 152532 86926 152544
rect 102134 152532 102140 152544
rect 102192 152532 102198 152584
rect 88334 152464 88340 152516
rect 88392 152504 88398 152516
rect 154206 152504 154212 152516
rect 88392 152476 154212 152504
rect 88392 152464 88398 152476
rect 154206 152464 154212 152476
rect 154264 152464 154270 152516
rect 209038 152464 209044 152516
rect 209096 152504 209102 152516
rect 220722 152504 220728 152516
rect 209096 152476 220728 152504
rect 209096 152464 209102 152476
rect 220722 152464 220728 152476
rect 220780 152504 220786 152516
rect 302234 152504 302240 152516
rect 220780 152476 302240 152504
rect 220780 152464 220786 152476
rect 302234 152464 302240 152476
rect 302292 152464 302298 152516
rect 180242 151852 180248 151904
rect 180300 151892 180306 151904
rect 208394 151892 208400 151904
rect 180300 151864 208400 151892
rect 180300 151852 180306 151864
rect 208394 151852 208400 151864
rect 208452 151852 208458 151904
rect 130470 151784 130476 151836
rect 130528 151824 130534 151836
rect 223666 151824 223672 151836
rect 130528 151796 223672 151824
rect 130528 151784 130534 151796
rect 223666 151784 223672 151796
rect 223724 151784 223730 151836
rect 208394 151036 208400 151088
rect 208452 151076 208458 151088
rect 225046 151076 225052 151088
rect 208452 151048 225052 151076
rect 208452 151036 208458 151048
rect 225046 151036 225052 151048
rect 225104 151036 225110 151088
rect 64690 150492 64696 150544
rect 64748 150532 64754 150544
rect 118050 150532 118056 150544
rect 64748 150504 118056 150532
rect 64748 150492 64754 150504
rect 118050 150492 118056 150504
rect 118108 150492 118114 150544
rect 206370 150492 206376 150544
rect 206428 150532 206434 150544
rect 304994 150532 305000 150544
rect 206428 150504 305000 150532
rect 206428 150492 206434 150504
rect 304994 150492 305000 150504
rect 305052 150492 305058 150544
rect 80514 150424 80520 150476
rect 80572 150464 80578 150476
rect 208394 150464 208400 150476
rect 80572 150436 208400 150464
rect 80572 150424 80578 150436
rect 208394 150424 208400 150436
rect 208452 150424 208458 150476
rect 67726 149676 67732 149728
rect 67784 149716 67790 149728
rect 159910 149716 159916 149728
rect 67784 149688 159916 149716
rect 67784 149676 67790 149688
rect 159910 149676 159916 149688
rect 159968 149716 159974 149728
rect 185486 149716 185492 149728
rect 159968 149688 185492 149716
rect 159968 149676 159974 149688
rect 185486 149676 185492 149688
rect 185544 149676 185550 149728
rect 196802 149676 196808 149728
rect 196860 149716 196866 149728
rect 209774 149716 209780 149728
rect 196860 149688 209780 149716
rect 196860 149676 196866 149688
rect 209774 149676 209780 149688
rect 209832 149676 209838 149728
rect 210234 149132 210240 149184
rect 210292 149172 210298 149184
rect 210418 149172 210424 149184
rect 210292 149144 210424 149172
rect 210292 149132 210298 149144
rect 210418 149132 210424 149144
rect 210476 149172 210482 149184
rect 243538 149172 243544 149184
rect 210476 149144 243544 149172
rect 210476 149132 210482 149144
rect 243538 149132 243544 149144
rect 243596 149132 243602 149184
rect 125410 149064 125416 149116
rect 125468 149104 125474 149116
rect 216766 149104 216772 149116
rect 125468 149076 216772 149104
rect 125468 149064 125474 149076
rect 216766 149064 216772 149076
rect 216824 149064 216830 149116
rect 239398 148316 239404 148368
rect 239456 148356 239462 148368
rect 256050 148356 256056 148368
rect 239456 148328 256056 148356
rect 239456 148316 239462 148328
rect 256050 148316 256056 148328
rect 256108 148316 256114 148368
rect 67542 147704 67548 147756
rect 67600 147744 67606 147756
rect 112530 147744 112536 147756
rect 67600 147716 112536 147744
rect 67600 147704 67606 147716
rect 112530 147704 112536 147716
rect 112588 147704 112594 147756
rect 167822 147704 167828 147756
rect 167880 147744 167886 147756
rect 168282 147744 168288 147756
rect 167880 147716 168288 147744
rect 167880 147704 167886 147716
rect 168282 147704 168288 147716
rect 168340 147744 168346 147756
rect 202138 147744 202144 147756
rect 168340 147716 202144 147744
rect 168340 147704 168346 147716
rect 202138 147704 202144 147716
rect 202196 147704 202202 147756
rect 206922 147704 206928 147756
rect 206980 147744 206986 147756
rect 320174 147744 320180 147756
rect 206980 147716 320180 147744
rect 206980 147704 206986 147716
rect 320174 147704 320180 147716
rect 320232 147704 320238 147756
rect 100110 147636 100116 147688
rect 100168 147676 100174 147688
rect 100662 147676 100668 147688
rect 100168 147648 100668 147676
rect 100168 147636 100174 147648
rect 100662 147636 100668 147648
rect 100720 147676 100726 147688
rect 227806 147676 227812 147688
rect 100720 147648 227812 147676
rect 100720 147636 100726 147648
rect 227806 147636 227812 147648
rect 227864 147636 227870 147688
rect 214006 147568 214012 147620
rect 214064 147608 214070 147620
rect 256694 147608 256700 147620
rect 214064 147580 256700 147608
rect 214064 147568 214070 147580
rect 256694 147568 256700 147580
rect 256752 147608 256758 147620
rect 257430 147608 257436 147620
rect 256752 147580 257436 147608
rect 256752 147568 256758 147580
rect 257430 147568 257436 147580
rect 257488 147568 257494 147620
rect 210694 147160 210700 147212
rect 210752 147200 210758 147212
rect 214006 147200 214012 147212
rect 210752 147172 214012 147200
rect 210752 147160 210758 147172
rect 214006 147160 214012 147172
rect 214064 147160 214070 147212
rect 3142 147024 3148 147076
rect 3200 147064 3206 147076
rect 95510 147064 95516 147076
rect 3200 147036 95516 147064
rect 3200 147024 3206 147036
rect 95510 147024 95516 147036
rect 95568 147064 95574 147076
rect 96522 147064 96528 147076
rect 95568 147036 96528 147064
rect 95568 147024 95574 147036
rect 96522 147024 96528 147036
rect 96580 147024 96586 147076
rect 83550 146956 83556 147008
rect 83608 146996 83614 147008
rect 90450 146996 90456 147008
rect 83608 146968 90456 146996
rect 83608 146956 83614 146968
rect 90450 146956 90456 146968
rect 90508 146956 90514 147008
rect 169018 146956 169024 147008
rect 169076 146996 169082 147008
rect 184382 146996 184388 147008
rect 169076 146968 184388 146996
rect 169076 146956 169082 146968
rect 184382 146956 184388 146968
rect 184440 146956 184446 147008
rect 193490 146956 193496 147008
rect 193548 146996 193554 147008
rect 207198 146996 207204 147008
rect 193548 146968 207204 146996
rect 193548 146956 193554 146968
rect 207198 146956 207204 146968
rect 207256 146956 207262 147008
rect 90910 146888 90916 146940
rect 90968 146928 90974 146940
rect 127618 146928 127624 146940
rect 90968 146900 127624 146928
rect 90968 146888 90974 146900
rect 127618 146888 127624 146900
rect 127676 146928 127682 146940
rect 220814 146928 220820 146940
rect 127676 146900 220820 146928
rect 127676 146888 127682 146900
rect 220814 146888 220820 146900
rect 220872 146888 220878 146940
rect 257430 146888 257436 146940
rect 257488 146928 257494 146940
rect 580258 146928 580264 146940
rect 257488 146900 580264 146928
rect 257488 146888 257494 146900
rect 580258 146888 580264 146900
rect 580316 146888 580322 146940
rect 213270 146208 213276 146260
rect 213328 146248 213334 146260
rect 216582 146248 216588 146260
rect 213328 146220 216588 146248
rect 213328 146208 213334 146220
rect 216582 146208 216588 146220
rect 216640 146208 216646 146260
rect 244366 146208 244372 146260
rect 244424 146248 244430 146260
rect 244918 146248 244924 146260
rect 244424 146220 244924 146248
rect 244424 146208 244430 146220
rect 244918 146208 244924 146220
rect 244976 146208 244982 146260
rect 197078 145596 197084 145648
rect 197136 145636 197142 145648
rect 213730 145636 213736 145648
rect 197136 145608 213736 145636
rect 197136 145596 197142 145608
rect 213730 145596 213736 145608
rect 213788 145596 213794 145648
rect 8938 145528 8944 145580
rect 8996 145568 9002 145580
rect 87506 145568 87512 145580
rect 8996 145540 87512 145568
rect 8996 145528 9002 145540
rect 87506 145528 87512 145540
rect 87564 145528 87570 145580
rect 114462 145528 114468 145580
rect 114520 145568 114526 145580
rect 180058 145568 180064 145580
rect 114520 145540 180064 145568
rect 114520 145528 114526 145540
rect 180058 145528 180064 145540
rect 180116 145528 180122 145580
rect 218974 145528 218980 145580
rect 219032 145568 219038 145580
rect 267826 145568 267832 145580
rect 219032 145540 267832 145568
rect 219032 145528 219038 145540
rect 267826 145528 267832 145540
rect 267884 145528 267890 145580
rect 282914 145528 282920 145580
rect 282972 145568 282978 145580
rect 298738 145568 298744 145580
rect 282972 145540 298744 145568
rect 282972 145528 282978 145540
rect 298738 145528 298744 145540
rect 298796 145528 298802 145580
rect 160922 144984 160928 145036
rect 160980 145024 160986 145036
rect 161290 145024 161296 145036
rect 160980 144996 161296 145024
rect 160980 144984 160986 144996
rect 161290 144984 161296 144996
rect 161348 145024 161354 145036
rect 193766 145024 193772 145036
rect 161348 144996 193772 145024
rect 161348 144984 161354 144996
rect 193766 144984 193772 144996
rect 193824 144984 193830 145036
rect 192570 144916 192576 144968
rect 192628 144956 192634 144968
rect 244366 144956 244372 144968
rect 192628 144928 244372 144956
rect 192628 144916 192634 144928
rect 244366 144916 244372 144928
rect 244424 144916 244430 144968
rect 87506 144848 87512 144900
rect 87564 144888 87570 144900
rect 125410 144888 125416 144900
rect 87564 144860 125416 144888
rect 87564 144848 87570 144860
rect 125410 144848 125416 144860
rect 125468 144848 125474 144900
rect 160830 144848 160836 144900
rect 160888 144888 160894 144900
rect 184290 144888 184296 144900
rect 160888 144860 184296 144888
rect 160888 144848 160894 144860
rect 184290 144848 184296 144860
rect 184348 144848 184354 144900
rect 97534 144304 97540 144356
rect 97592 144344 97598 144356
rect 99374 144344 99380 144356
rect 97592 144316 99380 144344
rect 97592 144304 97598 144316
rect 99374 144304 99380 144316
rect 99432 144304 99438 144356
rect 185486 144168 185492 144220
rect 185544 144208 185550 144220
rect 193582 144208 193588 144220
rect 185544 144180 193588 144208
rect 185544 144168 185550 144180
rect 193582 144168 193588 144180
rect 193640 144168 193646 144220
rect 173342 144100 173348 144152
rect 173400 144140 173406 144152
rect 180242 144140 180248 144152
rect 173400 144112 180248 144140
rect 173400 144100 173406 144112
rect 180242 144100 180248 144112
rect 180300 144100 180306 144152
rect 186958 143624 186964 143676
rect 187016 143664 187022 143676
rect 226334 143664 226340 143676
rect 187016 143636 226340 143664
rect 187016 143624 187022 143636
rect 226334 143624 226340 143636
rect 226392 143624 226398 143676
rect 66070 143556 66076 143608
rect 66128 143596 66134 143608
rect 91646 143596 91652 143608
rect 66128 143568 91652 143596
rect 66128 143556 66134 143568
rect 91646 143556 91652 143568
rect 91704 143556 91710 143608
rect 224126 143556 224132 143608
rect 224184 143596 224190 143608
rect 224310 143596 224316 143608
rect 224184 143568 224316 143596
rect 224184 143556 224190 143568
rect 224310 143556 224316 143568
rect 224368 143596 224374 143608
rect 313274 143596 313280 143608
rect 224368 143568 313280 143596
rect 224368 143556 224374 143568
rect 313274 143556 313280 143568
rect 313332 143556 313338 143608
rect 208118 143488 208124 143540
rect 208176 143528 208182 143540
rect 209038 143528 209044 143540
rect 208176 143500 209044 143528
rect 208176 143488 208182 143500
rect 209038 143488 209044 143500
rect 209096 143488 209102 143540
rect 69658 142808 69664 142860
rect 69716 142848 69722 142860
rect 83458 142848 83464 142860
rect 69716 142820 83464 142848
rect 69716 142808 69722 142820
rect 83458 142808 83464 142820
rect 83516 142808 83522 142860
rect 86034 142808 86040 142860
rect 86092 142848 86098 142860
rect 86770 142848 86776 142860
rect 86092 142820 86776 142848
rect 86092 142808 86098 142820
rect 86770 142808 86776 142820
rect 86828 142848 86834 142860
rect 215294 142848 215300 142860
rect 86828 142820 215300 142848
rect 86828 142808 86834 142820
rect 215294 142808 215300 142820
rect 215352 142848 215358 142860
rect 216122 142848 216128 142860
rect 215352 142820 216128 142848
rect 215352 142808 215358 142820
rect 216122 142808 216128 142820
rect 216180 142808 216186 142860
rect 217318 142400 217324 142452
rect 217376 142440 217382 142452
rect 218238 142440 218244 142452
rect 217376 142412 218244 142440
rect 217376 142400 217382 142412
rect 218238 142400 218244 142412
rect 218296 142400 218302 142452
rect 220078 142196 220084 142248
rect 220136 142236 220142 142248
rect 228358 142236 228364 142248
rect 220136 142208 228364 142236
rect 220136 142196 220142 142208
rect 228358 142196 228364 142208
rect 228416 142196 228422 142248
rect 78950 142128 78956 142180
rect 79008 142168 79014 142180
rect 206370 142168 206376 142180
rect 79008 142140 206376 142168
rect 79008 142128 79014 142140
rect 206370 142128 206376 142140
rect 206428 142128 206434 142180
rect 213178 142128 213184 142180
rect 213236 142168 213242 142180
rect 232590 142168 232596 142180
rect 213236 142140 232596 142168
rect 213236 142128 213242 142140
rect 232590 142128 232596 142140
rect 232648 142128 232654 142180
rect 80422 141448 80428 141500
rect 80480 141488 80486 141500
rect 103514 141488 103520 141500
rect 80480 141460 103520 141488
rect 80480 141448 80486 141460
rect 103514 141448 103520 141460
rect 103572 141488 103578 141500
rect 104710 141488 104716 141500
rect 103572 141460 104716 141488
rect 103572 141448 103578 141460
rect 104710 141448 104716 141460
rect 104768 141448 104774 141500
rect 70302 141380 70308 141432
rect 70360 141420 70366 141432
rect 105078 141420 105084 141432
rect 70360 141392 105084 141420
rect 70360 141380 70366 141392
rect 105078 141380 105084 141392
rect 105136 141380 105142 141432
rect 173802 141380 173808 141432
rect 173860 141420 173866 141432
rect 200758 141420 200764 141432
rect 173860 141392 200764 141420
rect 173860 141380 173866 141392
rect 200758 141380 200764 141392
rect 200816 141380 200822 141432
rect 203426 140836 203432 140888
rect 203484 140876 203490 140888
rect 289078 140876 289084 140888
rect 203484 140848 289084 140876
rect 203484 140836 203490 140848
rect 289078 140836 289084 140848
rect 289136 140836 289142 140888
rect 104710 140768 104716 140820
rect 104768 140808 104774 140820
rect 207750 140808 207756 140820
rect 104768 140780 207756 140808
rect 104768 140768 104774 140780
rect 207750 140768 207756 140780
rect 207808 140768 207814 140820
rect 215018 140768 215024 140820
rect 215076 140808 215082 140820
rect 255314 140808 255320 140820
rect 215076 140780 255320 140808
rect 215076 140768 215082 140780
rect 255314 140768 255320 140780
rect 255372 140768 255378 140820
rect 71314 140700 71320 140752
rect 71372 140740 71378 140752
rect 73062 140740 73068 140752
rect 71372 140712 73068 140740
rect 71372 140700 71378 140712
rect 73062 140700 73068 140712
rect 73120 140740 73126 140752
rect 189074 140740 189080 140752
rect 73120 140712 189080 140740
rect 73120 140700 73126 140712
rect 189074 140700 189080 140712
rect 189132 140700 189138 140752
rect 218698 140700 218704 140752
rect 218756 140740 218762 140752
rect 221826 140740 221832 140752
rect 218756 140712 221832 140740
rect 218756 140700 218762 140712
rect 221826 140700 221832 140712
rect 221884 140700 221890 140752
rect 195946 140576 205634 140604
rect 64506 140020 64512 140072
rect 64564 140060 64570 140072
rect 70394 140060 70400 140072
rect 64564 140032 70400 140060
rect 64564 140020 64570 140032
rect 70394 140020 70400 140032
rect 70452 140020 70458 140072
rect 184842 139544 184848 139596
rect 184900 139584 184906 139596
rect 195946 139584 195974 140576
rect 198642 140496 198648 140548
rect 198700 140496 198706 140548
rect 184900 139556 195974 139584
rect 184900 139544 184906 139556
rect 67818 139408 67824 139460
rect 67876 139448 67882 139460
rect 100202 139448 100208 139460
rect 67876 139420 100208 139448
rect 67876 139408 67882 139420
rect 100202 139408 100208 139420
rect 100260 139408 100266 139460
rect 198660 139380 198688 140496
rect 205606 140468 205634 140576
rect 210050 140496 210056 140548
rect 210108 140536 210114 140548
rect 210108 140508 218652 140536
rect 210108 140496 210114 140508
rect 205910 140468 205916 140480
rect 205606 140440 205916 140468
rect 205910 140428 205916 140440
rect 205968 140468 205974 140480
rect 206922 140468 206928 140480
rect 205968 140440 206928 140468
rect 205968 140428 205974 140440
rect 206922 140428 206928 140440
rect 206980 140428 206986 140480
rect 218514 140428 218520 140480
rect 218572 140428 218578 140480
rect 180766 139352 198688 139380
rect 218532 139380 218560 140428
rect 218624 140060 218652 140508
rect 222010 140428 222016 140480
rect 222068 140468 222074 140480
rect 225230 140468 225236 140480
rect 222068 140440 225236 140468
rect 222068 140428 222074 140440
rect 225230 140428 225236 140440
rect 225288 140428 225294 140480
rect 264882 140088 264888 140140
rect 264940 140128 264946 140140
rect 276014 140128 276020 140140
rect 264940 140100 276020 140128
rect 264940 140088 264946 140100
rect 276014 140088 276020 140100
rect 276072 140088 276078 140140
rect 287698 140060 287704 140072
rect 218624 140032 287704 140060
rect 287698 140020 287704 140032
rect 287756 140020 287762 140072
rect 225230 139408 225236 139460
rect 225288 139448 225294 139460
rect 264882 139448 264888 139460
rect 225288 139420 264888 139448
rect 225288 139408 225294 139420
rect 264882 139408 264888 139420
rect 264940 139408 264946 139460
rect 278774 139380 278780 139392
rect 218532 139352 278780 139380
rect 52178 138660 52184 138712
rect 52236 138700 52242 138712
rect 72510 138700 72516 138712
rect 52236 138672 72516 138700
rect 52236 138660 52242 138672
rect 72510 138660 72516 138672
rect 72568 138660 72574 138712
rect 90818 138660 90824 138712
rect 90876 138700 90882 138712
rect 163590 138700 163596 138712
rect 90876 138672 163596 138700
rect 90876 138660 90882 138672
rect 163590 138660 163596 138672
rect 163648 138660 163654 138712
rect 87046 138592 87052 138644
rect 87104 138632 87110 138644
rect 180766 138632 180794 139352
rect 278774 139340 278780 139352
rect 278832 139380 278838 139392
rect 280062 139380 280068 139392
rect 278832 139352 280068 139380
rect 278832 139340 278838 139352
rect 280062 139340 280068 139352
rect 280120 139340 280126 139392
rect 280062 138660 280068 138712
rect 280120 138700 280126 138712
rect 322198 138700 322204 138712
rect 280120 138672 322204 138700
rect 280120 138660 280126 138672
rect 322198 138660 322204 138672
rect 322256 138660 322262 138712
rect 87104 138604 180794 138632
rect 87104 138592 87110 138604
rect 78858 138048 78864 138100
rect 78916 138088 78922 138100
rect 79502 138088 79508 138100
rect 78916 138060 79508 138088
rect 78916 138048 78922 138060
rect 79502 138048 79508 138060
rect 79560 138048 79566 138100
rect 3602 137980 3608 138032
rect 3660 138020 3666 138032
rect 75822 138020 75828 138032
rect 3660 137992 75828 138020
rect 3660 137980 3666 137992
rect 75822 137980 75828 137992
rect 75880 137980 75886 138032
rect 3510 137912 3516 137964
rect 3568 137952 3574 137964
rect 72970 137952 72976 137964
rect 3568 137924 72976 137952
rect 3568 137912 3574 137924
rect 72970 137912 72976 137924
rect 73028 137912 73034 137964
rect 78858 137912 78864 137964
rect 78916 137952 78922 137964
rect 79318 137952 79324 137964
rect 78916 137924 79324 137952
rect 78916 137912 78922 137924
rect 79318 137912 79324 137924
rect 79376 137912 79382 137964
rect 184842 137952 184848 137964
rect 89686 137924 184848 137952
rect 77846 137844 77852 137896
rect 77904 137884 77910 137896
rect 81342 137884 81348 137896
rect 77904 137856 81348 137884
rect 77904 137844 77910 137856
rect 81342 137844 81348 137856
rect 81400 137844 81406 137896
rect 69382 137776 69388 137828
rect 69440 137816 69446 137828
rect 75270 137816 75276 137828
rect 69440 137788 75276 137816
rect 69440 137776 69446 137788
rect 75270 137776 75276 137788
rect 75328 137776 75334 137828
rect 79318 137708 79324 137760
rect 79376 137748 79382 137760
rect 89686 137748 89714 137924
rect 184842 137912 184848 137924
rect 184900 137912 184906 137964
rect 101398 137844 101404 137896
rect 101456 137884 101462 137896
rect 102042 137884 102048 137896
rect 101456 137856 102048 137884
rect 101456 137844 101462 137856
rect 102042 137844 102048 137856
rect 102100 137884 102106 137896
rect 192570 137884 192576 137896
rect 102100 137856 192576 137884
rect 102100 137844 102106 137856
rect 192570 137844 192576 137856
rect 192628 137844 192634 137896
rect 79376 137720 89714 137748
rect 79376 137708 79382 137720
rect 229738 137028 229744 137080
rect 229796 137068 229802 137080
rect 237374 137068 237380 137080
rect 229796 137040 237380 137068
rect 229796 137028 229802 137040
rect 237374 137028 237380 137040
rect 237432 137028 237438 137080
rect 89346 136960 89352 137012
rect 89404 137000 89410 137012
rect 90358 137000 90364 137012
rect 89404 136972 90364 137000
rect 89404 136960 89410 136972
rect 90358 136960 90364 136972
rect 90416 136960 90422 137012
rect 83366 136688 83372 136740
rect 83424 136728 83430 136740
rect 86218 136728 86224 136740
rect 83424 136700 86224 136728
rect 83424 136688 83430 136700
rect 86218 136688 86224 136700
rect 86276 136688 86282 136740
rect 81342 136620 81348 136672
rect 81400 136660 81406 136672
rect 83550 136660 83556 136672
rect 81400 136632 83556 136660
rect 81400 136620 81406 136632
rect 83550 136620 83556 136632
rect 83608 136620 83614 136672
rect 85942 136620 85948 136672
rect 86000 136660 86006 136672
rect 87046 136660 87052 136672
rect 86000 136632 87052 136660
rect 86000 136620 86006 136632
rect 87046 136620 87052 136632
rect 87104 136620 87110 136672
rect 90266 136620 90272 136672
rect 90324 136660 90330 136672
rect 91738 136660 91744 136672
rect 90324 136632 91744 136660
rect 90324 136620 90330 136632
rect 91738 136620 91744 136632
rect 91796 136620 91802 136672
rect 92382 136620 92388 136672
rect 92440 136660 92446 136672
rect 93118 136660 93124 136672
rect 92440 136632 93124 136660
rect 92440 136620 92446 136632
rect 93118 136620 93124 136632
rect 93176 136620 93182 136672
rect 91646 136552 91652 136604
rect 91704 136592 91710 136604
rect 166350 136592 166356 136604
rect 91704 136564 166356 136592
rect 91704 136552 91710 136564
rect 166350 136552 166356 136564
rect 166408 136552 166414 136604
rect 184382 136552 184388 136604
rect 184440 136592 184446 136604
rect 191558 136592 191564 136604
rect 184440 136564 191564 136592
rect 184440 136552 184446 136564
rect 191558 136552 191564 136564
rect 191616 136552 191622 136604
rect 11698 135940 11704 135992
rect 11756 135980 11762 135992
rect 91002 135980 91008 135992
rect 11756 135952 91008 135980
rect 11756 135940 11762 135952
rect 91002 135940 91008 135952
rect 91060 135940 91066 135992
rect 69566 135872 69572 135924
rect 69624 135912 69630 135924
rect 160922 135912 160928 135924
rect 69624 135884 160928 135912
rect 69624 135872 69630 135884
rect 160922 135872 160928 135884
rect 160980 135872 160986 135924
rect 180058 135260 180064 135312
rect 180116 135300 180122 135312
rect 191558 135300 191564 135312
rect 180116 135272 191564 135300
rect 180116 135260 180122 135272
rect 191558 135260 191564 135272
rect 191616 135260 191622 135312
rect 75638 135192 75644 135244
rect 75696 135232 75702 135244
rect 94130 135232 94136 135244
rect 75696 135204 94136 135232
rect 75696 135192 75702 135204
rect 94130 135192 94136 135204
rect 94188 135192 94194 135244
rect 96706 135192 96712 135244
rect 96764 135232 96770 135244
rect 145650 135232 145656 135244
rect 96764 135204 145656 135232
rect 96764 135192 96770 135204
rect 145650 135192 145656 135204
rect 145708 135192 145714 135244
rect 188430 135192 188436 135244
rect 188488 135232 188494 135244
rect 192846 135232 192852 135244
rect 188488 135204 192852 135232
rect 188488 135192 188494 135204
rect 192846 135192 192852 135204
rect 192904 135192 192910 135244
rect 227070 135192 227076 135244
rect 227128 135232 227134 135244
rect 227898 135232 227904 135244
rect 227128 135204 227904 135232
rect 227128 135192 227134 135204
rect 227898 135192 227904 135204
rect 227956 135232 227962 135244
rect 267734 135232 267740 135244
rect 227956 135204 267740 135232
rect 227956 135192 227962 135204
rect 267734 135192 267740 135204
rect 267792 135192 267798 135244
rect 68830 134580 68836 134632
rect 68888 134620 68894 134632
rect 74534 134620 74540 134632
rect 68888 134592 74540 134620
rect 68888 134580 68894 134592
rect 74534 134580 74540 134592
rect 74592 134620 74598 134632
rect 75638 134620 75644 134632
rect 74592 134592 75644 134620
rect 74592 134580 74598 134592
rect 75638 134580 75644 134592
rect 75696 134580 75702 134632
rect 226702 134512 226708 134564
rect 226760 134552 226766 134564
rect 278038 134552 278044 134564
rect 226760 134524 278044 134552
rect 226760 134512 226766 134524
rect 278038 134512 278044 134524
rect 278096 134512 278102 134564
rect 130470 134008 130476 134020
rect 103486 133980 130476 134008
rect 94682 133900 94688 133952
rect 94740 133940 94746 133952
rect 103486 133940 103514 133980
rect 130470 133968 130476 133980
rect 130528 133968 130534 134020
rect 94740 133912 103514 133940
rect 94740 133900 94746 133912
rect 181530 133900 181536 133952
rect 181588 133940 181594 133952
rect 193030 133940 193036 133952
rect 181588 133912 193036 133940
rect 181588 133900 181594 133912
rect 193030 133900 193036 133912
rect 193088 133900 193094 133952
rect 226334 133900 226340 133952
rect 226392 133900 226398 133952
rect 127710 133832 127716 133884
rect 127768 133872 127774 133884
rect 182910 133872 182916 133884
rect 127768 133844 182916 133872
rect 127768 133832 127774 133844
rect 182910 133832 182916 133844
rect 182968 133832 182974 133884
rect 226352 133804 226380 133900
rect 226702 133832 226708 133884
rect 226760 133872 226766 133884
rect 229278 133872 229284 133884
rect 226760 133844 229284 133872
rect 226760 133832 226766 133844
rect 229278 133832 229284 133844
rect 229336 133832 229342 133884
rect 269114 133872 269120 133884
rect 238726 133844 269120 133872
rect 238726 133804 238754 133844
rect 269114 133832 269120 133844
rect 269172 133872 269178 133884
rect 273898 133872 273904 133884
rect 269172 133844 273904 133872
rect 269172 133832 269178 133844
rect 273898 133832 273904 133844
rect 273956 133832 273962 133884
rect 226352 133776 238754 133804
rect 96706 133288 96712 133340
rect 96764 133328 96770 133340
rect 102778 133328 102784 133340
rect 96764 133300 102784 133328
rect 96764 133288 96770 133300
rect 102778 133288 102784 133300
rect 102836 133288 102842 133340
rect 53466 133152 53472 133204
rect 53524 133192 53530 133204
rect 66346 133192 66352 133204
rect 53524 133164 66352 133192
rect 53524 133152 53530 133164
rect 66346 133152 66352 133164
rect 66404 133152 66410 133204
rect 153930 133152 153936 133204
rect 153988 133192 153994 133204
rect 187142 133192 187148 133204
rect 153988 133164 187148 133192
rect 153988 133152 153994 133164
rect 187142 133152 187148 133164
rect 187200 133152 187206 133204
rect 50706 132404 50712 132456
rect 50764 132444 50770 132456
rect 66254 132444 66260 132456
rect 50764 132416 66260 132444
rect 50764 132404 50770 132416
rect 66254 132404 66260 132416
rect 66312 132404 66318 132456
rect 96614 132404 96620 132456
rect 96672 132444 96678 132456
rect 186958 132444 186964 132456
rect 96672 132416 186964 132444
rect 96672 132404 96678 132416
rect 186958 132404 186964 132416
rect 187016 132404 187022 132456
rect 226702 132404 226708 132456
rect 226760 132444 226766 132456
rect 238754 132444 238760 132456
rect 226760 132416 238760 132444
rect 226760 132404 226766 132416
rect 238754 132404 238760 132416
rect 238812 132404 238818 132456
rect 142982 132336 142988 132388
rect 143040 132376 143046 132388
rect 191650 132376 191656 132388
rect 143040 132348 191656 132376
rect 143040 132336 143046 132348
rect 191650 132336 191656 132348
rect 191708 132336 191714 132388
rect 104158 131044 104164 131096
rect 104216 131084 104222 131096
rect 156598 131084 156604 131096
rect 104216 131056 156604 131084
rect 104216 131044 104222 131056
rect 156598 131044 156604 131056
rect 156656 131084 156662 131096
rect 188430 131084 188436 131096
rect 156656 131056 188436 131084
rect 156656 131044 156662 131056
rect 188430 131044 188436 131056
rect 188488 131044 188494 131096
rect 226702 131044 226708 131096
rect 226760 131084 226766 131096
rect 230566 131084 230572 131096
rect 226760 131056 230572 131084
rect 226760 131044 226766 131056
rect 230566 131044 230572 131056
rect 230624 131084 230630 131096
rect 276106 131084 276112 131096
rect 230624 131056 276112 131084
rect 230624 131044 230630 131056
rect 276106 131044 276112 131056
rect 276164 131044 276170 131096
rect 96614 130976 96620 131028
rect 96672 131016 96678 131028
rect 135898 131016 135904 131028
rect 96672 130988 135904 131016
rect 96672 130976 96678 130988
rect 135898 130976 135904 130988
rect 135956 130976 135962 131028
rect 97902 129684 97908 129736
rect 97960 129724 97966 129736
rect 177390 129724 177396 129736
rect 97960 129696 177396 129724
rect 97960 129684 97966 129696
rect 177390 129684 177396 129696
rect 177448 129684 177454 129736
rect 226702 129684 226708 129736
rect 226760 129724 226766 129736
rect 266446 129724 266452 129736
rect 226760 129696 266452 129724
rect 226760 129684 226766 129696
rect 266446 129684 266452 129696
rect 266504 129724 266510 129736
rect 267826 129724 267832 129736
rect 266504 129696 267832 129724
rect 266504 129684 266510 129696
rect 267826 129684 267832 129696
rect 267884 129684 267890 129736
rect 96706 129616 96712 129668
rect 96764 129656 96770 129668
rect 115198 129656 115204 129668
rect 96764 129628 115204 129656
rect 96764 129616 96770 129628
rect 115198 129616 115204 129628
rect 115256 129616 115262 129668
rect 118050 129004 118056 129056
rect 118108 129044 118114 129056
rect 169754 129044 169760 129056
rect 118108 129016 169760 129044
rect 118108 129004 118114 129016
rect 169754 129004 169760 129016
rect 169812 129004 169818 129056
rect 226702 129004 226708 129056
rect 226760 129044 226766 129056
rect 299474 129044 299480 129056
rect 226760 129016 299480 129044
rect 226760 129004 226766 129016
rect 299474 129004 299480 129016
rect 299532 129004 299538 129056
rect 169754 128324 169760 128376
rect 169812 128364 169818 128376
rect 171042 128364 171048 128376
rect 169812 128336 171048 128364
rect 169812 128324 169818 128336
rect 171042 128324 171048 128336
rect 171100 128364 171106 128376
rect 191650 128364 191656 128376
rect 171100 128336 191656 128364
rect 171100 128324 171106 128336
rect 191650 128324 191656 128336
rect 191708 128324 191714 128376
rect 61746 128256 61752 128308
rect 61804 128296 61810 128308
rect 66806 128296 66812 128308
rect 61804 128268 66812 128296
rect 61804 128256 61810 128268
rect 66806 128256 66812 128268
rect 66864 128256 66870 128308
rect 100202 128256 100208 128308
rect 100260 128296 100266 128308
rect 181530 128296 181536 128308
rect 100260 128268 181536 128296
rect 100260 128256 100266 128268
rect 181530 128256 181536 128268
rect 181588 128256 181594 128308
rect 226610 128256 226616 128308
rect 226668 128296 226674 128308
rect 245654 128296 245660 128308
rect 226668 128268 245660 128296
rect 226668 128256 226674 128268
rect 245654 128256 245660 128268
rect 245712 128256 245718 128308
rect 97902 128188 97908 128240
rect 97960 128228 97966 128240
rect 151170 128228 151176 128240
rect 97960 128200 151176 128228
rect 97960 128188 97966 128200
rect 151170 128188 151176 128200
rect 151228 128188 151234 128240
rect 245654 127576 245660 127628
rect 245712 127616 245718 127628
rect 323578 127616 323584 127628
rect 245712 127588 323584 127616
rect 245712 127576 245718 127588
rect 323578 127576 323584 127588
rect 323636 127576 323642 127628
rect 54938 126896 54944 126948
rect 54996 126936 55002 126948
rect 66806 126936 66812 126948
rect 54996 126908 66812 126936
rect 54996 126896 55002 126908
rect 66806 126896 66812 126908
rect 66864 126896 66870 126948
rect 94958 126896 94964 126948
rect 95016 126936 95022 126948
rect 180150 126936 180156 126948
rect 95016 126908 180156 126936
rect 95016 126896 95022 126908
rect 180150 126896 180156 126908
rect 180208 126896 180214 126948
rect 188890 126896 188896 126948
rect 188948 126936 188954 126948
rect 191650 126936 191656 126948
rect 188948 126908 191656 126936
rect 188948 126896 188954 126908
rect 191650 126896 191656 126908
rect 191708 126896 191714 126948
rect 226334 126896 226340 126948
rect 226392 126936 226398 126948
rect 252554 126936 252560 126948
rect 226392 126908 252560 126936
rect 226392 126896 226398 126908
rect 252554 126896 252560 126908
rect 252612 126936 252618 126948
rect 253014 126936 253020 126948
rect 252612 126908 253020 126936
rect 252612 126896 252618 126908
rect 253014 126896 253020 126908
rect 253072 126896 253078 126948
rect 97166 126828 97172 126880
rect 97224 126868 97230 126880
rect 105538 126868 105544 126880
rect 97224 126840 105544 126868
rect 97224 126828 97230 126840
rect 105538 126828 105544 126840
rect 105596 126828 105602 126880
rect 226702 126828 226708 126880
rect 226760 126868 226766 126880
rect 234614 126868 234620 126880
rect 226760 126840 234620 126868
rect 226760 126828 226766 126840
rect 234614 126828 234620 126840
rect 234672 126828 234678 126880
rect 105630 126216 105636 126268
rect 105688 126256 105694 126268
rect 155310 126256 155316 126268
rect 105688 126228 155316 126256
rect 105688 126216 105694 126228
rect 155310 126216 155316 126228
rect 155368 126216 155374 126268
rect 253014 126216 253020 126268
rect 253072 126256 253078 126268
rect 349154 126256 349160 126268
rect 253072 126228 349160 126256
rect 253072 126216 253078 126228
rect 349154 126216 349160 126228
rect 349212 126216 349218 126268
rect 57606 125536 57612 125588
rect 57664 125576 57670 125588
rect 66806 125576 66812 125588
rect 57664 125548 66812 125576
rect 57664 125536 57670 125548
rect 66806 125536 66812 125548
rect 66864 125536 66870 125588
rect 97442 125536 97448 125588
rect 97500 125576 97506 125588
rect 173250 125576 173256 125588
rect 97500 125548 173256 125576
rect 97500 125536 97506 125548
rect 173250 125536 173256 125548
rect 173308 125536 173314 125588
rect 257338 125536 257344 125588
rect 257396 125576 257402 125588
rect 280246 125576 280252 125588
rect 257396 125548 280252 125576
rect 257396 125536 257402 125548
rect 280246 125536 280252 125548
rect 280304 125576 280310 125588
rect 281442 125576 281448 125588
rect 280304 125548 281448 125576
rect 280304 125536 280310 125548
rect 281442 125536 281448 125548
rect 281500 125536 281506 125588
rect 156690 125468 156696 125520
rect 156748 125508 156754 125520
rect 190362 125508 190368 125520
rect 156748 125480 190368 125508
rect 156748 125468 156754 125480
rect 190362 125468 190368 125480
rect 190420 125468 190426 125520
rect 226702 125468 226708 125520
rect 226760 125508 226766 125520
rect 259454 125508 259460 125520
rect 226760 125480 259460 125508
rect 226760 125468 226766 125480
rect 259454 125468 259460 125480
rect 259512 125468 259518 125520
rect 64690 124924 64696 124976
rect 64748 124964 64754 124976
rect 66898 124964 66904 124976
rect 64748 124936 66904 124964
rect 64748 124924 64754 124936
rect 66898 124924 66904 124936
rect 66956 124924 66962 124976
rect 281442 124856 281448 124908
rect 281500 124896 281506 124908
rect 316034 124896 316040 124908
rect 281500 124868 316040 124896
rect 281500 124856 281506 124868
rect 316034 124856 316040 124868
rect 316092 124856 316098 124908
rect 61838 124108 61844 124160
rect 61896 124148 61902 124160
rect 66622 124148 66628 124160
rect 61896 124120 66628 124148
rect 61896 124108 61902 124120
rect 66622 124108 66628 124120
rect 66680 124108 66686 124160
rect 94590 124108 94596 124160
rect 94648 124148 94654 124160
rect 184198 124148 184204 124160
rect 94648 124120 184204 124148
rect 94648 124108 94654 124120
rect 184198 124108 184204 124120
rect 184256 124108 184262 124160
rect 226702 124108 226708 124160
rect 226760 124148 226766 124160
rect 236086 124148 236092 124160
rect 226760 124120 236092 124148
rect 226760 124108 226766 124120
rect 236086 124108 236092 124120
rect 236144 124148 236150 124160
rect 287146 124148 287152 124160
rect 236144 124120 287152 124148
rect 236144 124108 236150 124120
rect 287146 124108 287152 124120
rect 287204 124148 287210 124160
rect 582742 124148 582748 124160
rect 287204 124120 582748 124148
rect 287204 124108 287210 124120
rect 582742 124108 582748 124120
rect 582800 124108 582806 124160
rect 178678 124040 178684 124092
rect 178736 124080 178742 124092
rect 190638 124080 190644 124092
rect 178736 124052 190644 124080
rect 178736 124040 178742 124052
rect 190638 124040 190644 124052
rect 190696 124040 190702 124092
rect 232498 123428 232504 123480
rect 232556 123468 232562 123480
rect 255958 123468 255964 123480
rect 232556 123440 255964 123468
rect 232556 123428 232562 123440
rect 255958 123428 255964 123440
rect 256016 123428 256022 123480
rect 187510 122816 187516 122868
rect 187568 122856 187574 122868
rect 191650 122856 191656 122868
rect 187568 122828 191656 122856
rect 187568 122816 187574 122828
rect 191650 122816 191656 122828
rect 191708 122816 191714 122868
rect 46750 122748 46756 122800
rect 46808 122788 46814 122800
rect 66806 122788 66812 122800
rect 46808 122760 66812 122788
rect 46808 122748 46814 122760
rect 66806 122748 66812 122760
rect 66864 122748 66870 122800
rect 97902 122748 97908 122800
rect 97960 122788 97966 122800
rect 116670 122788 116676 122800
rect 97960 122760 116676 122788
rect 97960 122748 97966 122760
rect 116670 122748 116676 122760
rect 116728 122748 116734 122800
rect 226334 122748 226340 122800
rect 226392 122788 226398 122800
rect 251266 122788 251272 122800
rect 226392 122760 251272 122788
rect 226392 122748 226398 122760
rect 251266 122748 251272 122760
rect 251324 122748 251330 122800
rect 182910 122068 182916 122120
rect 182968 122108 182974 122120
rect 183462 122108 183468 122120
rect 182968 122080 183468 122108
rect 182968 122068 182974 122080
rect 183462 122068 183468 122080
rect 183520 122108 183526 122120
rect 191650 122108 191656 122120
rect 183520 122080 191656 122108
rect 183520 122068 183526 122080
rect 191650 122068 191656 122080
rect 191708 122068 191714 122120
rect 60458 121388 60464 121440
rect 60516 121428 60522 121440
rect 66806 121428 66812 121440
rect 60516 121400 66812 121428
rect 60516 121388 60522 121400
rect 66806 121388 66812 121400
rect 66864 121388 66870 121440
rect 97166 121388 97172 121440
rect 97224 121428 97230 121440
rect 153930 121428 153936 121440
rect 97224 121400 153936 121428
rect 97224 121388 97230 121400
rect 153930 121388 153936 121400
rect 153988 121388 153994 121440
rect 226702 121388 226708 121440
rect 226760 121428 226766 121440
rect 233234 121428 233240 121440
rect 226760 121400 233240 121428
rect 226760 121388 226766 121400
rect 233234 121388 233240 121400
rect 233292 121388 233298 121440
rect 60550 121320 60556 121372
rect 60608 121360 60614 121372
rect 66622 121360 66628 121372
rect 60608 121332 66628 121360
rect 60608 121320 60614 121332
rect 66622 121320 66628 121332
rect 66680 121320 66686 121372
rect 170950 120776 170956 120828
rect 171008 120816 171014 120828
rect 184842 120816 184848 120828
rect 171008 120788 184848 120816
rect 171008 120776 171014 120788
rect 184842 120776 184848 120788
rect 184900 120776 184906 120828
rect 102870 120708 102876 120760
rect 102928 120748 102934 120760
rect 183370 120748 183376 120760
rect 102928 120720 183376 120748
rect 102928 120708 102934 120720
rect 183370 120708 183376 120720
rect 183428 120708 183434 120760
rect 232590 120708 232596 120760
rect 232648 120748 232654 120760
rect 295334 120748 295340 120760
rect 232648 120720 295340 120748
rect 232648 120708 232654 120720
rect 295334 120708 295340 120720
rect 295392 120708 295398 120760
rect 96062 120300 96068 120352
rect 96120 120340 96126 120352
rect 98730 120340 98736 120352
rect 96120 120312 98736 120340
rect 96120 120300 96126 120312
rect 98730 120300 98736 120312
rect 98788 120300 98794 120352
rect 183370 120096 183376 120148
rect 183428 120136 183434 120148
rect 188982 120136 188988 120148
rect 183428 120108 188988 120136
rect 183428 120096 183434 120108
rect 188982 120096 188988 120108
rect 189040 120096 189046 120148
rect 56410 120028 56416 120080
rect 56468 120068 56474 120080
rect 66806 120068 66812 120080
rect 56468 120040 66812 120068
rect 56468 120028 56474 120040
rect 66806 120028 66812 120040
rect 66864 120028 66870 120080
rect 158070 120028 158076 120080
rect 158128 120068 158134 120080
rect 187510 120068 187516 120080
rect 158128 120040 187516 120068
rect 158128 120028 158134 120040
rect 187510 120028 187516 120040
rect 187568 120028 187574 120080
rect 188338 120028 188344 120080
rect 188396 120068 188402 120080
rect 191650 120068 191656 120080
rect 188396 120040 191656 120068
rect 188396 120028 188402 120040
rect 191650 120028 191656 120040
rect 191708 120028 191714 120080
rect 226518 119824 226524 119876
rect 226576 119864 226582 119876
rect 229094 119864 229100 119876
rect 226576 119836 229100 119864
rect 226576 119824 226582 119836
rect 229094 119824 229100 119836
rect 229152 119824 229158 119876
rect 3418 119348 3424 119400
rect 3476 119388 3482 119400
rect 53834 119388 53840 119400
rect 3476 119360 53840 119388
rect 3476 119348 3482 119360
rect 53834 119348 53840 119360
rect 53892 119348 53898 119400
rect 112530 119348 112536 119400
rect 112588 119388 112594 119400
rect 184290 119388 184296 119400
rect 112588 119360 184296 119388
rect 112588 119348 112594 119360
rect 184290 119348 184296 119360
rect 184348 119348 184354 119400
rect 233234 119348 233240 119400
rect 233292 119388 233298 119400
rect 260834 119388 260840 119400
rect 233292 119360 260840 119388
rect 233292 119348 233298 119360
rect 260834 119348 260840 119360
rect 260892 119348 260898 119400
rect 98730 118940 98736 118992
rect 98788 118980 98794 118992
rect 103698 118980 103704 118992
rect 98788 118952 103704 118980
rect 98788 118940 98794 118952
rect 103698 118940 103704 118952
rect 103756 118940 103762 118992
rect 97258 118668 97264 118720
rect 97316 118708 97322 118720
rect 100938 118708 100944 118720
rect 97316 118680 100944 118708
rect 97316 118668 97322 118680
rect 100938 118668 100944 118680
rect 100996 118668 101002 118720
rect 186958 118668 186964 118720
rect 187016 118708 187022 118720
rect 187510 118708 187516 118720
rect 187016 118680 187516 118708
rect 187016 118668 187022 118680
rect 187510 118668 187516 118680
rect 187568 118668 187574 118720
rect 97902 118600 97908 118652
rect 97960 118640 97966 118652
rect 108482 118640 108488 118652
rect 97960 118612 108488 118640
rect 97960 118600 97966 118612
rect 108482 118600 108488 118612
rect 108540 118600 108546 118652
rect 226610 118600 226616 118652
rect 226668 118640 226674 118652
rect 231854 118640 231860 118652
rect 226668 118612 231860 118640
rect 226668 118600 226674 118612
rect 231854 118600 231860 118612
rect 231912 118640 231918 118652
rect 233142 118640 233148 118652
rect 231912 118612 233148 118640
rect 231912 118600 231918 118612
rect 233142 118600 233148 118612
rect 233200 118600 233206 118652
rect 53558 118532 53564 118584
rect 53616 118572 53622 118584
rect 66254 118572 66260 118584
rect 53616 118544 66260 118572
rect 53616 118532 53622 118544
rect 66254 118532 66260 118544
rect 66312 118532 66318 118584
rect 97810 118192 97816 118244
rect 97868 118232 97874 118244
rect 105630 118232 105636 118244
rect 97868 118204 105636 118232
rect 97868 118192 97874 118204
rect 105630 118192 105636 118204
rect 105688 118192 105694 118244
rect 233142 117920 233148 117972
rect 233200 117960 233206 117972
rect 304258 117960 304264 117972
rect 233200 117932 304264 117960
rect 233200 117920 233206 117932
rect 304258 117920 304264 117932
rect 304316 117920 304322 117972
rect 63218 117240 63224 117292
rect 63276 117280 63282 117292
rect 66254 117280 66260 117292
rect 63276 117252 66260 117280
rect 63276 117240 63282 117252
rect 66254 117240 66260 117252
rect 66312 117240 66318 117292
rect 97902 117240 97908 117292
rect 97960 117280 97966 117292
rect 169294 117280 169300 117292
rect 97960 117252 169300 117280
rect 97960 117240 97966 117252
rect 169294 117240 169300 117252
rect 169352 117240 169358 117292
rect 184842 117240 184848 117292
rect 184900 117280 184906 117292
rect 191650 117280 191656 117292
rect 184900 117252 191656 117280
rect 184900 117240 184906 117252
rect 191650 117240 191656 117252
rect 191708 117240 191714 117292
rect 63126 117172 63132 117224
rect 63184 117212 63190 117224
rect 66898 117212 66904 117224
rect 63184 117184 66904 117212
rect 63184 117172 63190 117184
rect 66898 117172 66904 117184
rect 66956 117172 66962 117224
rect 97810 117172 97816 117224
rect 97868 117212 97874 117224
rect 148410 117212 148416 117224
rect 97868 117184 148416 117212
rect 97868 117172 97874 117184
rect 148410 117172 148416 117184
rect 148468 117172 148474 117224
rect 226702 116628 226708 116680
rect 226760 116668 226766 116680
rect 233234 116668 233240 116680
rect 226760 116640 233240 116668
rect 226760 116628 226766 116640
rect 233234 116628 233240 116640
rect 233292 116628 233298 116680
rect 226334 116560 226340 116612
rect 226392 116600 226398 116612
rect 258166 116600 258172 116612
rect 226392 116572 258172 116600
rect 226392 116560 226398 116572
rect 258166 116560 258172 116572
rect 258224 116560 258230 116612
rect 188430 116016 188436 116068
rect 188488 116056 188494 116068
rect 190638 116056 190644 116068
rect 188488 116028 190644 116056
rect 188488 116016 188494 116028
rect 190638 116016 190644 116028
rect 190696 116016 190702 116068
rect 50798 115880 50804 115932
rect 50856 115920 50862 115932
rect 66806 115920 66812 115932
rect 50856 115892 66812 115920
rect 50856 115880 50862 115892
rect 66806 115880 66812 115892
rect 66864 115880 66870 115932
rect 97902 115880 97908 115932
rect 97960 115920 97966 115932
rect 187050 115920 187056 115932
rect 97960 115892 187056 115920
rect 97960 115880 97966 115892
rect 187050 115880 187056 115892
rect 187108 115880 187114 115932
rect 97810 115812 97816 115864
rect 97868 115852 97874 115864
rect 173342 115852 173348 115864
rect 97868 115824 173348 115852
rect 97868 115812 97874 115824
rect 173342 115812 173348 115824
rect 173400 115812 173406 115864
rect 226518 115200 226524 115252
rect 226576 115240 226582 115252
rect 229094 115240 229100 115252
rect 226576 115212 229100 115240
rect 226576 115200 226582 115212
rect 229094 115200 229100 115212
rect 229152 115240 229158 115252
rect 273346 115240 273352 115252
rect 229152 115212 273352 115240
rect 229152 115200 229158 115212
rect 273346 115200 273352 115212
rect 273404 115200 273410 115252
rect 62022 114452 62028 114504
rect 62080 114492 62086 114504
rect 66806 114492 66812 114504
rect 62080 114464 66812 114492
rect 62080 114452 62086 114464
rect 66806 114452 66812 114464
rect 66864 114452 66870 114504
rect 53834 113772 53840 113824
rect 53892 113812 53898 113824
rect 62022 113812 62028 113824
rect 53892 113784 62028 113812
rect 53892 113772 53898 113784
rect 62022 113772 62028 113784
rect 62080 113812 62086 113824
rect 66898 113812 66904 113824
rect 62080 113784 66904 113812
rect 62080 113772 62086 113784
rect 66898 113772 66904 113784
rect 66956 113772 66962 113824
rect 228358 113772 228364 113824
rect 228416 113812 228422 113824
rect 252554 113812 252560 113824
rect 228416 113784 252560 113812
rect 228416 113772 228422 113784
rect 252554 113772 252560 113784
rect 252612 113772 252618 113824
rect 97534 113160 97540 113212
rect 97592 113200 97598 113212
rect 187142 113200 187148 113212
rect 97592 113172 187148 113200
rect 97592 113160 97598 113172
rect 187142 113160 187148 113172
rect 187200 113160 187206 113212
rect 188246 113160 188252 113212
rect 188304 113200 188310 113212
rect 191006 113200 191012 113212
rect 188304 113172 191012 113200
rect 188304 113160 188310 113172
rect 191006 113160 191012 113172
rect 191064 113160 191070 113212
rect 227346 113160 227352 113212
rect 227404 113200 227410 113212
rect 244458 113200 244464 113212
rect 227404 113172 244464 113200
rect 227404 113160 227410 113172
rect 244458 113160 244464 113172
rect 244516 113160 244522 113212
rect 157242 112412 157248 112464
rect 157300 112452 157306 112464
rect 191742 112452 191748 112464
rect 157300 112424 191748 112452
rect 157300 112412 157306 112424
rect 191742 112412 191748 112424
rect 191800 112412 191806 112464
rect 97902 111868 97908 111920
rect 97960 111908 97966 111920
rect 153838 111908 153844 111920
rect 97960 111880 153844 111908
rect 97960 111868 97966 111880
rect 153838 111868 153844 111880
rect 153896 111868 153902 111920
rect 156598 111868 156604 111920
rect 156656 111908 156662 111920
rect 157242 111908 157248 111920
rect 156656 111880 157248 111908
rect 156656 111868 156662 111880
rect 157242 111868 157248 111880
rect 157300 111868 157306 111920
rect 97810 111800 97816 111852
rect 97868 111840 97874 111852
rect 177390 111840 177396 111852
rect 97868 111812 177396 111840
rect 97868 111800 97874 111812
rect 177390 111800 177396 111812
rect 177448 111800 177454 111852
rect 238110 111800 238116 111852
rect 238168 111840 238174 111852
rect 324314 111840 324320 111852
rect 238168 111812 324320 111840
rect 238168 111800 238174 111812
rect 324314 111800 324320 111812
rect 324372 111800 324378 111852
rect 3142 111732 3148 111784
rect 3200 111772 3206 111784
rect 11698 111772 11704 111784
rect 3200 111744 11704 111772
rect 3200 111732 3206 111744
rect 11698 111732 11704 111744
rect 11756 111732 11762 111784
rect 225322 111732 225328 111784
rect 225380 111772 225386 111784
rect 241514 111772 241520 111784
rect 225380 111744 241520 111772
rect 225380 111732 225386 111744
rect 241514 111732 241520 111744
rect 241572 111732 241578 111784
rect 57514 111052 57520 111104
rect 57572 111092 57578 111104
rect 66162 111092 66168 111104
rect 57572 111064 66168 111092
rect 57572 111052 57578 111064
rect 66162 111052 66168 111064
rect 66220 111092 66226 111104
rect 66622 111092 66628 111104
rect 66220 111064 66628 111092
rect 66220 111052 66226 111064
rect 66622 111052 66628 111064
rect 66680 111052 66686 111104
rect 96798 111052 96804 111104
rect 96856 111092 96862 111104
rect 100110 111092 100116 111104
rect 96856 111064 100116 111092
rect 96856 111052 96862 111064
rect 100110 111052 100116 111064
rect 100168 111052 100174 111104
rect 226518 111052 226524 111104
rect 226576 111092 226582 111104
rect 240686 111092 240692 111104
rect 226576 111064 240692 111092
rect 226576 111052 226582 111064
rect 240686 111052 240692 111064
rect 240744 111092 240750 111104
rect 291838 111092 291844 111104
rect 240744 111064 291844 111092
rect 240744 111052 240750 111064
rect 291838 111052 291844 111064
rect 291896 111052 291902 111104
rect 184750 110848 184756 110900
rect 184808 110888 184814 110900
rect 190362 110888 190368 110900
rect 184808 110860 190368 110888
rect 184808 110848 184814 110860
rect 190362 110848 190368 110860
rect 190420 110848 190426 110900
rect 187694 110440 187700 110492
rect 187752 110480 187758 110492
rect 191742 110480 191748 110492
rect 187752 110452 191748 110480
rect 187752 110440 187758 110452
rect 191742 110440 191748 110452
rect 191800 110440 191806 110492
rect 97442 110236 97448 110288
rect 97500 110276 97506 110288
rect 100754 110276 100760 110288
rect 97500 110248 100760 110276
rect 97500 110236 97506 110248
rect 100754 110236 100760 110248
rect 100812 110236 100818 110288
rect 55122 109692 55128 109744
rect 55180 109732 55186 109744
rect 60734 109732 60740 109744
rect 55180 109704 60740 109732
rect 55180 109692 55186 109704
rect 60734 109692 60740 109704
rect 60792 109692 60798 109744
rect 116578 109692 116584 109744
rect 116636 109732 116642 109744
rect 188246 109732 188252 109744
rect 116636 109704 188252 109732
rect 116636 109692 116642 109704
rect 188246 109692 188252 109704
rect 188304 109692 188310 109744
rect 226978 109692 226984 109744
rect 227036 109732 227042 109744
rect 262398 109732 262404 109744
rect 227036 109704 262404 109732
rect 227036 109692 227042 109704
rect 262398 109692 262404 109704
rect 262456 109692 262462 109744
rect 60734 109012 60740 109064
rect 60792 109052 60798 109064
rect 61378 109052 61384 109064
rect 60792 109024 61384 109052
rect 60792 109012 60798 109024
rect 61378 109012 61384 109024
rect 61436 109052 61442 109064
rect 66806 109052 66812 109064
rect 61436 109024 66812 109052
rect 61436 109012 61442 109024
rect 66806 109012 66812 109024
rect 66864 109012 66870 109064
rect 97166 109012 97172 109064
rect 97224 109052 97230 109064
rect 160830 109052 160836 109064
rect 97224 109024 160836 109052
rect 97224 109012 97230 109024
rect 160830 109012 160836 109024
rect 160888 109012 160894 109064
rect 187050 109012 187056 109064
rect 187108 109052 187114 109064
rect 191558 109052 191564 109064
rect 187108 109024 191564 109052
rect 187108 109012 187114 109024
rect 191558 109012 191564 109024
rect 191616 109012 191622 109064
rect 59078 108944 59084 108996
rect 59136 108984 59142 108996
rect 66898 108984 66904 108996
rect 59136 108956 66904 108984
rect 59136 108944 59142 108956
rect 66898 108944 66904 108956
rect 66956 108944 66962 108996
rect 160738 108944 160744 108996
rect 160796 108984 160802 108996
rect 187694 108984 187700 108996
rect 160796 108956 187700 108984
rect 160796 108944 160802 108956
rect 187694 108944 187700 108956
rect 187752 108944 187758 108996
rect 97902 108332 97908 108384
rect 97960 108372 97966 108384
rect 109034 108372 109040 108384
rect 97960 108344 109040 108372
rect 97960 108332 97966 108344
rect 109034 108332 109040 108344
rect 109092 108372 109098 108384
rect 109678 108372 109684 108384
rect 109092 108344 109684 108372
rect 109092 108332 109098 108344
rect 109678 108332 109684 108344
rect 109736 108332 109742 108384
rect 225046 108332 225052 108384
rect 225104 108372 225110 108384
rect 225230 108372 225236 108384
rect 225104 108344 225236 108372
rect 225104 108332 225110 108344
rect 225230 108332 225236 108344
rect 225288 108332 225294 108384
rect 230382 108332 230388 108384
rect 230440 108372 230446 108384
rect 244274 108372 244280 108384
rect 230440 108344 244280 108372
rect 230440 108332 230446 108344
rect 244274 108332 244280 108344
rect 244332 108332 244338 108384
rect 95970 108264 95976 108316
rect 96028 108304 96034 108316
rect 107654 108304 107660 108316
rect 96028 108276 107660 108304
rect 96028 108264 96034 108276
rect 107654 108264 107660 108276
rect 107712 108304 107718 108316
rect 173250 108304 173256 108316
rect 107712 108276 173256 108304
rect 107712 108264 107718 108276
rect 173250 108264 173256 108276
rect 173308 108264 173314 108316
rect 233142 108264 233148 108316
rect 233200 108304 233206 108316
rect 288526 108304 288532 108316
rect 233200 108276 288532 108304
rect 233200 108264 233206 108276
rect 288526 108264 288532 108276
rect 288584 108264 288590 108316
rect 225046 108196 225052 108248
rect 225104 108236 225110 108248
rect 225322 108236 225328 108248
rect 225104 108208 225328 108236
rect 225104 108196 225110 108208
rect 225322 108196 225328 108208
rect 225380 108196 225386 108248
rect 187602 107788 187608 107840
rect 187660 107828 187666 107840
rect 189074 107828 189080 107840
rect 187660 107800 189080 107828
rect 187660 107788 187666 107800
rect 189074 107788 189080 107800
rect 189132 107828 189138 107840
rect 191742 107828 191748 107840
rect 189132 107800 191748 107828
rect 189132 107788 189138 107800
rect 191742 107788 191748 107800
rect 191800 107788 191806 107840
rect 226610 107720 226616 107772
rect 226668 107760 226674 107772
rect 229186 107760 229192 107772
rect 226668 107732 229192 107760
rect 226668 107720 226674 107732
rect 229186 107720 229192 107732
rect 229244 107760 229250 107772
rect 230382 107760 230388 107772
rect 229244 107732 230388 107760
rect 229244 107720 229250 107732
rect 230382 107720 230388 107732
rect 230440 107720 230446 107772
rect 63310 107652 63316 107704
rect 63368 107692 63374 107704
rect 66806 107692 66812 107704
rect 63368 107664 66812 107692
rect 63368 107652 63374 107664
rect 66806 107652 66812 107664
rect 66864 107652 66870 107704
rect 226702 107652 226708 107704
rect 226760 107692 226766 107704
rect 231946 107692 231952 107704
rect 226760 107664 231952 107692
rect 226760 107652 226766 107664
rect 231946 107652 231952 107664
rect 232004 107692 232010 107704
rect 233142 107692 233148 107704
rect 232004 107664 233148 107692
rect 232004 107652 232010 107664
rect 233142 107652 233148 107664
rect 233200 107652 233206 107704
rect 52270 107584 52276 107636
rect 52328 107624 52334 107636
rect 66898 107624 66904 107636
rect 52328 107596 66904 107624
rect 52328 107584 52334 107596
rect 66898 107584 66904 107596
rect 66956 107584 66962 107636
rect 162762 107584 162768 107636
rect 162820 107624 162826 107636
rect 191558 107624 191564 107636
rect 162820 107596 191564 107624
rect 162820 107584 162826 107596
rect 191558 107584 191564 107596
rect 191616 107584 191622 107636
rect 50614 106904 50620 106956
rect 50672 106944 50678 106956
rect 59078 106944 59084 106956
rect 50672 106916 59084 106944
rect 50672 106904 50678 106916
rect 59078 106904 59084 106916
rect 59136 106904 59142 106956
rect 97534 106360 97540 106412
rect 97592 106400 97598 106412
rect 101490 106400 101496 106412
rect 97592 106372 101496 106400
rect 97592 106360 97598 106372
rect 101490 106360 101496 106372
rect 101548 106360 101554 106412
rect 59078 106292 59084 106344
rect 59136 106332 59142 106344
rect 66806 106332 66812 106344
rect 59136 106304 66812 106332
rect 59136 106292 59142 106304
rect 66806 106292 66812 106304
rect 66864 106292 66870 106344
rect 97902 106292 97908 106344
rect 97960 106332 97966 106344
rect 184198 106332 184204 106344
rect 97960 106304 184204 106332
rect 97960 106292 97966 106304
rect 184198 106292 184204 106304
rect 184256 106292 184262 106344
rect 226702 106292 226708 106344
rect 226760 106332 226766 106344
rect 230566 106332 230572 106344
rect 226760 106304 230572 106332
rect 226760 106292 226766 106304
rect 230566 106292 230572 106304
rect 230624 106332 230630 106344
rect 353294 106332 353300 106344
rect 230624 106304 353300 106332
rect 230624 106292 230630 106304
rect 353294 106292 353300 106304
rect 353352 106292 353358 106344
rect 97534 106224 97540 106276
rect 97592 106264 97598 106276
rect 120074 106264 120080 106276
rect 97592 106236 120080 106264
rect 97592 106224 97598 106236
rect 120074 106224 120080 106236
rect 120132 106224 120138 106276
rect 184290 105884 184296 105936
rect 184348 105924 184354 105936
rect 191742 105924 191748 105936
rect 184348 105896 191748 105924
rect 184348 105884 184354 105896
rect 191742 105884 191748 105896
rect 191800 105884 191806 105936
rect 166350 105612 166356 105664
rect 166408 105652 166414 105664
rect 190454 105652 190460 105664
rect 166408 105624 190460 105652
rect 166408 105612 166414 105624
rect 190454 105612 190460 105624
rect 190512 105612 190518 105664
rect 48130 105544 48136 105596
rect 48188 105584 48194 105596
rect 65978 105584 65984 105596
rect 48188 105556 65984 105584
rect 48188 105544 48194 105556
rect 65978 105544 65984 105556
rect 66036 105584 66042 105596
rect 66530 105584 66536 105596
rect 66036 105556 66536 105584
rect 66036 105544 66042 105556
rect 66530 105544 66536 105556
rect 66588 105544 66594 105596
rect 97902 105544 97908 105596
rect 97960 105584 97966 105596
rect 100846 105584 100852 105596
rect 97960 105556 100852 105584
rect 97960 105544 97966 105556
rect 100846 105544 100852 105556
rect 100904 105584 100910 105596
rect 180150 105584 180156 105596
rect 100904 105556 180156 105584
rect 100904 105544 100910 105556
rect 180150 105544 180156 105556
rect 180208 105544 180214 105596
rect 226334 105544 226340 105596
rect 226392 105584 226398 105596
rect 270494 105584 270500 105596
rect 226392 105556 270500 105584
rect 226392 105544 226398 105556
rect 270494 105544 270500 105556
rect 270552 105544 270558 105596
rect 270494 105136 270500 105188
rect 270552 105176 270558 105188
rect 271138 105176 271144 105188
rect 270552 105148 271144 105176
rect 270552 105136 270558 105148
rect 271138 105136 271144 105148
rect 271196 105136 271202 105188
rect 59170 104796 59176 104848
rect 59228 104836 59234 104848
rect 66254 104836 66260 104848
rect 59228 104808 66260 104836
rect 59228 104796 59234 104808
rect 66254 104796 66260 104808
rect 66312 104796 66318 104848
rect 226518 104796 226524 104848
rect 226576 104836 226582 104848
rect 244274 104836 244280 104848
rect 226576 104808 244280 104836
rect 226576 104796 226582 104808
rect 244274 104796 244280 104808
rect 244332 104796 244338 104848
rect 97902 104116 97908 104168
rect 97960 104156 97966 104168
rect 106274 104156 106280 104168
rect 97960 104128 106280 104156
rect 97960 104116 97966 104128
rect 106274 104116 106280 104128
rect 106332 104116 106338 104168
rect 180242 104116 180248 104168
rect 180300 104156 180306 104168
rect 191650 104156 191656 104168
rect 180300 104128 191656 104156
rect 180300 104116 180306 104128
rect 191650 104116 191656 104128
rect 191708 104116 191714 104168
rect 244274 104116 244280 104168
rect 244332 104156 244338 104168
rect 284938 104156 284944 104168
rect 244332 104128 284944 104156
rect 244332 104116 244338 104128
rect 284938 104116 284944 104128
rect 284996 104116 285002 104168
rect 162118 103544 162124 103556
rect 135226 103516 162124 103544
rect 97902 103436 97908 103488
rect 97960 103476 97966 103488
rect 134610 103476 134616 103488
rect 97960 103448 134616 103476
rect 97960 103436 97966 103448
rect 134610 103436 134616 103448
rect 134668 103476 134674 103488
rect 135226 103476 135254 103516
rect 162118 103504 162124 103516
rect 162176 103504 162182 103556
rect 134668 103448 135254 103476
rect 134668 103436 134674 103448
rect 97718 103368 97724 103420
rect 97776 103408 97782 103420
rect 101398 103408 101404 103420
rect 97776 103380 101404 103408
rect 97776 103368 97782 103380
rect 101398 103368 101404 103380
rect 101456 103368 101462 103420
rect 64782 102348 64788 102400
rect 64840 102388 64846 102400
rect 66070 102388 66076 102400
rect 64840 102360 66076 102388
rect 64840 102348 64846 102360
rect 66070 102348 66076 102360
rect 66128 102388 66134 102400
rect 66530 102388 66536 102400
rect 66128 102360 66536 102388
rect 66128 102348 66134 102360
rect 66530 102348 66536 102360
rect 66588 102348 66594 102400
rect 188338 102144 188344 102196
rect 188396 102184 188402 102196
rect 191006 102184 191012 102196
rect 188396 102156 191012 102184
rect 188396 102144 188402 102156
rect 191006 102144 191012 102156
rect 191064 102144 191070 102196
rect 226610 102144 226616 102196
rect 226668 102184 226674 102196
rect 231854 102184 231860 102196
rect 226668 102156 231860 102184
rect 226668 102144 226674 102156
rect 231854 102144 231860 102156
rect 231912 102184 231918 102196
rect 269758 102184 269764 102196
rect 231912 102156 269764 102184
rect 231912 102144 231918 102156
rect 269758 102144 269764 102156
rect 269816 102144 269822 102196
rect 226702 102076 226708 102128
rect 226760 102116 226766 102128
rect 266354 102116 266360 102128
rect 226760 102088 266360 102116
rect 226760 102076 226766 102088
rect 266354 102076 266360 102088
rect 266412 102076 266418 102128
rect 98822 101396 98828 101448
rect 98880 101436 98886 101448
rect 160094 101436 160100 101448
rect 98880 101408 160100 101436
rect 98880 101396 98886 101408
rect 160094 101396 160100 101408
rect 160152 101436 160158 101448
rect 187694 101436 187700 101448
rect 160152 101408 187700 101436
rect 160152 101396 160158 101408
rect 187694 101396 187700 101408
rect 187752 101396 187758 101448
rect 59262 101260 59268 101312
rect 59320 101300 59326 101312
rect 61838 101300 61844 101312
rect 59320 101272 61844 101300
rect 59320 101260 59326 101272
rect 61838 101260 61844 101272
rect 61896 101300 61902 101312
rect 66438 101300 66444 101312
rect 61896 101272 66444 101300
rect 61896 101260 61902 101272
rect 66438 101260 66444 101272
rect 66496 101260 66502 101312
rect 187694 100988 187700 101040
rect 187752 101028 187758 101040
rect 188982 101028 188988 101040
rect 187752 101000 188988 101028
rect 187752 100988 187758 101000
rect 188982 100988 188988 101000
rect 189040 101028 189046 101040
rect 190638 101028 190644 101040
rect 189040 101000 190644 101028
rect 189040 100988 189046 101000
rect 190638 100988 190644 101000
rect 190696 100988 190702 101040
rect 53742 100716 53748 100768
rect 53800 100756 53806 100768
rect 57882 100756 57888 100768
rect 53800 100728 57888 100756
rect 53800 100716 53806 100728
rect 57882 100716 57888 100728
rect 57940 100756 57946 100768
rect 66806 100756 66812 100768
rect 57940 100728 66812 100756
rect 57940 100716 57946 100728
rect 66806 100716 66812 100728
rect 66864 100716 66870 100768
rect 97626 100716 97632 100768
rect 97684 100756 97690 100768
rect 169018 100756 169024 100768
rect 97684 100728 169024 100756
rect 97684 100716 97690 100728
rect 169018 100716 169024 100728
rect 169076 100716 169082 100768
rect 175182 100648 175188 100700
rect 175240 100688 175246 100700
rect 190638 100688 190644 100700
rect 175240 100660 190644 100688
rect 175240 100648 175246 100660
rect 190638 100648 190644 100660
rect 190696 100648 190702 100700
rect 57790 99968 57796 100020
rect 57848 100008 57854 100020
rect 64782 100008 64788 100020
rect 57848 99980 64788 100008
rect 57848 99968 57854 99980
rect 64782 99968 64788 99980
rect 64840 100008 64846 100020
rect 66806 100008 66812 100020
rect 64840 99980 66812 100008
rect 64840 99968 64846 99980
rect 66806 99968 66812 99980
rect 66864 99968 66870 100020
rect 227530 99968 227536 100020
rect 227588 100008 227594 100020
rect 227990 100008 227996 100020
rect 227588 99980 227996 100008
rect 227588 99968 227594 99980
rect 227990 99968 227996 99980
rect 228048 100008 228054 100020
rect 247034 100008 247040 100020
rect 228048 99980 247040 100008
rect 228048 99968 228054 99980
rect 247034 99968 247040 99980
rect 247092 100008 247098 100020
rect 327718 100008 327724 100020
rect 247092 99980 327724 100008
rect 247092 99968 247098 99980
rect 327718 99968 327724 99980
rect 327776 99968 327782 100020
rect 97810 99424 97816 99476
rect 97868 99464 97874 99476
rect 128262 99464 128268 99476
rect 97868 99436 128268 99464
rect 97868 99424 97874 99436
rect 128262 99424 128268 99436
rect 128320 99424 128326 99476
rect 97902 99356 97908 99408
rect 97960 99396 97966 99408
rect 173342 99396 173348 99408
rect 97960 99368 173348 99396
rect 97960 99356 97966 99368
rect 173342 99356 173348 99368
rect 173400 99356 173406 99408
rect 61930 99288 61936 99340
rect 61988 99328 61994 99340
rect 66622 99328 66628 99340
rect 61988 99300 66628 99328
rect 61988 99288 61994 99300
rect 66622 99288 66628 99300
rect 66680 99288 66686 99340
rect 97810 99288 97816 99340
rect 97868 99328 97874 99340
rect 132586 99328 132592 99340
rect 97868 99300 132592 99328
rect 97868 99288 97874 99300
rect 132586 99288 132592 99300
rect 132644 99328 132650 99340
rect 133782 99328 133788 99340
rect 132644 99300 133788 99328
rect 132644 99288 132650 99300
rect 133782 99288 133788 99300
rect 133840 99288 133846 99340
rect 226150 99288 226156 99340
rect 226208 99328 226214 99340
rect 287054 99328 287060 99340
rect 226208 99300 287060 99328
rect 226208 99288 226214 99300
rect 287054 99288 287060 99300
rect 287112 99328 287118 99340
rect 288342 99328 288348 99340
rect 287112 99300 288348 99328
rect 287112 99288 287118 99300
rect 288342 99288 288348 99300
rect 288400 99288 288406 99340
rect 97534 99084 97540 99136
rect 97592 99124 97598 99136
rect 99282 99124 99288 99136
rect 97592 99096 99288 99124
rect 97592 99084 97598 99096
rect 99282 99084 99288 99096
rect 99340 99124 99346 99136
rect 100018 99124 100024 99136
rect 99340 99096 100024 99124
rect 99340 99084 99346 99096
rect 100018 99084 100024 99096
rect 100076 99084 100082 99136
rect 133782 98608 133788 98660
rect 133840 98648 133846 98660
rect 178770 98648 178776 98660
rect 133840 98620 178776 98648
rect 133840 98608 133846 98620
rect 178770 98608 178776 98620
rect 178828 98608 178834 98660
rect 288342 98608 288348 98660
rect 288400 98648 288406 98660
rect 331214 98648 331220 98660
rect 288400 98620 331220 98648
rect 288400 98608 288406 98620
rect 331214 98608 331220 98620
rect 331272 98608 331278 98660
rect 188522 98064 188528 98116
rect 188580 98104 188586 98116
rect 191742 98104 191748 98116
rect 188580 98076 191748 98104
rect 188580 98064 188586 98076
rect 191742 98064 191748 98076
rect 191800 98064 191806 98116
rect 225046 98064 225052 98116
rect 225104 98064 225110 98116
rect 101398 97996 101404 98048
rect 101456 98036 101462 98048
rect 190822 98036 190828 98048
rect 101456 98008 190828 98036
rect 101456 97996 101462 98008
rect 190822 97996 190828 98008
rect 190880 97996 190886 98048
rect 225064 97912 225092 98064
rect 226610 97928 226616 97980
rect 226668 97968 226674 97980
rect 232498 97968 232504 97980
rect 226668 97940 232504 97968
rect 226668 97928 226674 97940
rect 232498 97928 232504 97940
rect 232556 97928 232562 97980
rect 225046 97860 225052 97912
rect 225104 97860 225110 97912
rect 96614 97656 96620 97708
rect 96672 97696 96678 97708
rect 98638 97696 98644 97708
rect 96672 97668 98644 97696
rect 96672 97656 96678 97668
rect 98638 97656 98644 97668
rect 98696 97656 98702 97708
rect 57698 97248 57704 97300
rect 57756 97288 57762 97300
rect 66622 97288 66628 97300
rect 57756 97260 66628 97288
rect 57756 97248 57762 97260
rect 66622 97248 66628 97260
rect 66680 97248 66686 97300
rect 100018 97248 100024 97300
rect 100076 97288 100082 97300
rect 188430 97288 188436 97300
rect 100076 97260 188436 97288
rect 100076 97248 100082 97260
rect 188430 97248 188436 97260
rect 188488 97248 188494 97300
rect 226426 96704 226432 96756
rect 226484 96744 226490 96756
rect 226702 96744 226708 96756
rect 226484 96716 226708 96744
rect 226484 96704 226490 96716
rect 226702 96704 226708 96716
rect 226760 96704 226766 96756
rect 3050 96636 3056 96688
rect 3108 96676 3114 96688
rect 57238 96676 57244 96688
rect 3108 96648 57244 96676
rect 3108 96636 3114 96648
rect 57238 96636 57244 96648
rect 57296 96636 57302 96688
rect 97902 96636 97908 96688
rect 97960 96676 97966 96688
rect 184290 96676 184296 96688
rect 97960 96648 184296 96676
rect 97960 96636 97966 96648
rect 184290 96636 184296 96648
rect 184348 96636 184354 96688
rect 226426 96568 226432 96620
rect 226484 96608 226490 96620
rect 262214 96608 262220 96620
rect 226484 96580 262220 96608
rect 226484 96568 226490 96580
rect 262214 96568 262220 96580
rect 262272 96568 262278 96620
rect 226610 96500 226616 96552
rect 226668 96540 226674 96552
rect 240778 96540 240784 96552
rect 226668 96512 240784 96540
rect 226668 96500 226674 96512
rect 240778 96500 240784 96512
rect 240836 96500 240842 96552
rect 97442 95888 97448 95940
rect 97500 95928 97506 95940
rect 169662 95928 169668 95940
rect 97500 95900 169668 95928
rect 97500 95888 97506 95900
rect 169662 95888 169668 95900
rect 169720 95928 169726 95940
rect 186130 95928 186136 95940
rect 169720 95900 186136 95928
rect 169720 95888 169726 95900
rect 186130 95888 186136 95900
rect 186188 95928 186194 95940
rect 191558 95928 191564 95940
rect 186188 95900 191564 95928
rect 186188 95888 186194 95900
rect 191558 95888 191564 95900
rect 191616 95888 191622 95940
rect 264238 95888 264244 95940
rect 264296 95928 264302 95940
rect 280154 95928 280160 95940
rect 264296 95900 280160 95928
rect 264296 95888 264302 95900
rect 280154 95888 280160 95900
rect 280212 95888 280218 95940
rect 97902 95208 97908 95260
rect 97960 95248 97966 95260
rect 191834 95248 191840 95260
rect 97960 95220 191840 95248
rect 97960 95208 97966 95220
rect 191834 95208 191840 95220
rect 191892 95208 191898 95260
rect 97810 95140 97816 95192
rect 97868 95180 97874 95192
rect 114554 95180 114560 95192
rect 97868 95152 114560 95180
rect 97868 95140 97874 95152
rect 114554 95140 114560 95152
rect 114612 95140 114618 95192
rect 226702 94528 226708 94580
rect 226760 94568 226766 94580
rect 240778 94568 240784 94580
rect 226760 94540 240784 94568
rect 226760 94528 226766 94540
rect 240778 94528 240784 94540
rect 240836 94528 240842 94580
rect 106182 94460 106188 94512
rect 106240 94500 106246 94512
rect 188430 94500 188436 94512
rect 106240 94472 188436 94500
rect 106240 94460 106246 94472
rect 188430 94460 188436 94472
rect 188488 94460 188494 94512
rect 226242 94460 226248 94512
rect 226300 94500 226306 94512
rect 245746 94500 245752 94512
rect 226300 94472 245752 94500
rect 226300 94460 226306 94472
rect 245746 94460 245752 94472
rect 245804 94460 245810 94512
rect 166902 93848 166908 93900
rect 166960 93888 166966 93900
rect 184842 93888 184848 93900
rect 166960 93860 184848 93888
rect 166960 93848 166966 93860
rect 184842 93848 184848 93860
rect 184900 93888 184906 93900
rect 191650 93888 191656 93900
rect 184900 93860 191656 93888
rect 184900 93848 184906 93860
rect 191650 93848 191656 93860
rect 191708 93848 191714 93900
rect 63402 93780 63408 93832
rect 63460 93820 63466 93832
rect 67818 93820 67824 93832
rect 63460 93792 67824 93820
rect 63460 93780 63466 93792
rect 67818 93780 67824 93792
rect 67876 93780 67882 93832
rect 95142 93100 95148 93152
rect 95200 93140 95206 93152
rect 165522 93140 165528 93152
rect 95200 93112 165528 93140
rect 95200 93100 95206 93112
rect 165522 93100 165528 93112
rect 165580 93140 165586 93152
rect 178678 93140 178684 93152
rect 165580 93112 178684 93140
rect 165580 93100 165586 93112
rect 178678 93100 178684 93112
rect 178736 93100 178742 93152
rect 249150 93100 249156 93152
rect 249208 93140 249214 93152
rect 262858 93140 262864 93152
rect 249208 93112 262864 93140
rect 249208 93100 249214 93112
rect 262858 93100 262864 93112
rect 262916 93100 262922 93152
rect 68922 92692 68928 92744
rect 68980 92732 68986 92744
rect 69704 92732 69710 92744
rect 68980 92704 69710 92732
rect 68980 92692 68986 92704
rect 69704 92692 69710 92704
rect 69762 92692 69768 92744
rect 72832 92692 72838 92744
rect 72890 92732 72896 92744
rect 72970 92732 72976 92744
rect 72890 92704 72976 92732
rect 72890 92692 72896 92704
rect 72970 92692 72976 92704
rect 73028 92692 73034 92744
rect 94360 92692 94366 92744
rect 94418 92732 94424 92744
rect 95234 92732 95240 92744
rect 94418 92704 95240 92732
rect 94418 92692 94424 92704
rect 95234 92692 95240 92704
rect 95292 92692 95298 92744
rect 90128 92624 90134 92676
rect 90186 92664 90192 92676
rect 91002 92664 91008 92676
rect 90186 92636 91008 92664
rect 90186 92624 90192 92636
rect 91002 92624 91008 92636
rect 91060 92624 91066 92676
rect 74534 92556 74540 92608
rect 74592 92596 74598 92608
rect 75776 92596 75782 92608
rect 74592 92568 75782 92596
rect 74592 92556 74598 92568
rect 75776 92556 75782 92568
rect 75834 92556 75840 92608
rect 185670 92596 185676 92608
rect 113146 92568 185676 92596
rect 48038 92488 48044 92540
rect 48096 92528 48102 92540
rect 70302 92528 70308 92540
rect 48096 92500 70308 92528
rect 48096 92488 48102 92500
rect 70302 92488 70308 92500
rect 70360 92488 70366 92540
rect 107010 92488 107016 92540
rect 107068 92528 107074 92540
rect 107654 92528 107660 92540
rect 107068 92500 107660 92528
rect 107068 92488 107074 92500
rect 107654 92488 107660 92500
rect 107712 92528 107718 92540
rect 113146 92528 113174 92568
rect 185670 92556 185676 92568
rect 185728 92556 185734 92608
rect 107712 92500 113174 92528
rect 107712 92488 107718 92500
rect 179230 92488 179236 92540
rect 179288 92528 179294 92540
rect 195974 92528 195980 92540
rect 179288 92500 195980 92528
rect 179288 92488 179294 92500
rect 195974 92488 195980 92500
rect 196032 92488 196038 92540
rect 224862 92488 224868 92540
rect 224920 92528 224926 92540
rect 242894 92528 242900 92540
rect 224920 92500 242900 92528
rect 224920 92488 224926 92500
rect 242894 92488 242900 92500
rect 242952 92488 242958 92540
rect 67358 92420 67364 92472
rect 67416 92460 67422 92472
rect 188522 92460 188528 92472
rect 67416 92432 188528 92460
rect 67416 92420 67422 92432
rect 188522 92420 188528 92432
rect 188580 92420 188586 92472
rect 193030 92420 193036 92472
rect 193088 92460 193094 92472
rect 202598 92460 202604 92472
rect 193088 92432 202604 92460
rect 193088 92420 193094 92432
rect 202598 92420 202604 92432
rect 202656 92420 202662 92472
rect 204162 92420 204168 92472
rect 204220 92460 204226 92472
rect 206094 92460 206100 92472
rect 204220 92432 206100 92460
rect 204220 92420 204226 92432
rect 206094 92420 206100 92432
rect 206152 92420 206158 92472
rect 67542 92352 67548 92404
rect 67600 92392 67606 92404
rect 166902 92392 166908 92404
rect 67600 92364 166908 92392
rect 67600 92352 67606 92364
rect 166902 92352 166908 92364
rect 166960 92352 166966 92404
rect 166166 91740 166172 91792
rect 166224 91780 166230 91792
rect 223574 91780 223580 91792
rect 166224 91752 223580 91780
rect 166224 91740 166230 91752
rect 223574 91740 223580 91752
rect 223632 91740 223638 91792
rect 222378 91168 222384 91180
rect 222212 91140 222384 91168
rect 64506 90992 64512 91044
rect 64564 91032 64570 91044
rect 70762 91032 70768 91044
rect 64564 91004 70768 91032
rect 64564 90992 64570 91004
rect 70762 90992 70768 91004
rect 70820 90992 70826 91044
rect 84654 90992 84660 91044
rect 84712 91032 84718 91044
rect 100754 91032 100760 91044
rect 84712 91004 100760 91032
rect 84712 90992 84718 91004
rect 100754 90992 100760 91004
rect 100812 91032 100818 91044
rect 179322 91032 179328 91044
rect 100812 91004 179328 91032
rect 100812 90992 100818 91004
rect 179322 90992 179328 91004
rect 179380 91032 179386 91044
rect 211798 91032 211804 91044
rect 179380 91004 211804 91032
rect 179380 90992 179386 91004
rect 211798 90992 211804 91004
rect 211856 90992 211862 91044
rect 222212 91032 222240 91140
rect 222378 91128 222384 91140
rect 222436 91168 222442 91180
rect 227714 91168 227720 91180
rect 222436 91140 227720 91168
rect 222436 91128 222442 91140
rect 227714 91128 227720 91140
rect 227772 91128 227778 91180
rect 224218 91060 224224 91112
rect 224276 91100 224282 91112
rect 225138 91100 225144 91112
rect 224276 91072 225144 91100
rect 224276 91060 224282 91072
rect 225138 91060 225144 91072
rect 225196 91060 225202 91112
rect 219406 91004 222240 91032
rect 172422 90924 172428 90976
rect 172480 90964 172486 90976
rect 194594 90964 194600 90976
rect 172480 90936 194600 90964
rect 172480 90924 172486 90936
rect 194594 90924 194600 90936
rect 194652 90924 194658 90976
rect 217134 90856 217140 90908
rect 217192 90896 217198 90908
rect 219406 90896 219434 91004
rect 222470 90992 222476 91044
rect 222528 91032 222534 91044
rect 241606 91032 241612 91044
rect 222528 91004 241612 91032
rect 222528 90992 222534 91004
rect 241606 90992 241612 91004
rect 241664 91032 241670 91044
rect 242158 91032 242164 91044
rect 241664 91004 242164 91032
rect 241664 90992 241670 91004
rect 242158 90992 242164 91004
rect 242216 90992 242222 91044
rect 221366 90924 221372 90976
rect 221424 90964 221430 90976
rect 226242 90964 226248 90976
rect 221424 90936 226248 90964
rect 221424 90924 221430 90936
rect 226242 90924 226248 90936
rect 226300 90924 226306 90976
rect 217192 90868 219434 90896
rect 217192 90856 217198 90868
rect 46842 90312 46848 90364
rect 46900 90352 46906 90364
rect 67542 90352 67548 90364
rect 46900 90324 67548 90352
rect 46900 90312 46906 90324
rect 67542 90312 67548 90324
rect 67600 90352 67606 90364
rect 68462 90352 68468 90364
rect 67600 90324 68468 90352
rect 67600 90312 67606 90324
rect 68462 90312 68468 90324
rect 68520 90312 68526 90364
rect 93854 90244 93860 90296
rect 93912 90284 93918 90296
rect 95050 90284 95056 90296
rect 93912 90256 95056 90284
rect 93912 90244 93918 90256
rect 95050 90244 95056 90256
rect 95108 90284 95114 90296
rect 95878 90284 95884 90296
rect 95108 90256 95884 90284
rect 95108 90244 95114 90256
rect 95878 90244 95884 90256
rect 95936 90244 95942 90296
rect 206278 89700 206284 89752
rect 206336 89740 206342 89752
rect 207934 89740 207940 89752
rect 206336 89712 207940 89740
rect 206336 89700 206342 89712
rect 207934 89700 207940 89712
rect 207992 89700 207998 89752
rect 67174 89632 67180 89684
rect 67232 89672 67238 89684
rect 101398 89672 101404 89684
rect 67232 89644 101404 89672
rect 67232 89632 67238 89644
rect 101398 89632 101404 89644
rect 101456 89632 101462 89684
rect 111794 89632 111800 89684
rect 111852 89672 111858 89684
rect 112438 89672 112444 89684
rect 111852 89644 112444 89672
rect 111852 89632 111858 89644
rect 112438 89632 112444 89644
rect 112496 89672 112502 89684
rect 209222 89672 209228 89684
rect 112496 89644 209228 89672
rect 112496 89632 112502 89644
rect 209222 89632 209228 89644
rect 209280 89632 209286 89684
rect 214558 89632 214564 89684
rect 214616 89672 214622 89684
rect 258074 89672 258080 89684
rect 214616 89644 258080 89672
rect 214616 89632 214622 89644
rect 258074 89632 258080 89644
rect 258132 89632 258138 89684
rect 75454 89564 75460 89616
rect 75512 89604 75518 89616
rect 95970 89604 95976 89616
rect 75512 89576 95976 89604
rect 75512 89564 75518 89576
rect 95970 89564 95976 89576
rect 96028 89564 96034 89616
rect 239398 89604 239404 89616
rect 219406 89576 239404 89604
rect 215846 89496 215852 89548
rect 215904 89536 215910 89548
rect 219406 89536 219434 89576
rect 239398 89564 239404 89576
rect 239456 89564 239462 89616
rect 215904 89508 219434 89536
rect 215904 89496 215910 89508
rect 209866 88476 209872 88528
rect 209924 88516 209930 88528
rect 210694 88516 210700 88528
rect 209924 88488 210700 88516
rect 209924 88476 209930 88488
rect 210694 88476 210700 88488
rect 210752 88476 210758 88528
rect 69198 88272 69204 88324
rect 69256 88312 69262 88324
rect 158714 88312 158720 88324
rect 69256 88284 158720 88312
rect 69256 88272 69262 88284
rect 158714 88272 158720 88284
rect 158772 88312 158778 88324
rect 193858 88312 193864 88324
rect 158772 88284 193864 88312
rect 158772 88272 158778 88284
rect 193858 88272 193864 88284
rect 193916 88312 193922 88324
rect 194134 88312 194140 88324
rect 193916 88284 194140 88312
rect 193916 88272 193922 88284
rect 194134 88272 194140 88284
rect 194192 88272 194198 88324
rect 204438 88272 204444 88324
rect 204496 88312 204502 88324
rect 208394 88312 208400 88324
rect 204496 88284 208400 88312
rect 204496 88272 204502 88284
rect 208394 88272 208400 88284
rect 208452 88272 208458 88324
rect 211614 88272 211620 88324
rect 211672 88312 211678 88324
rect 263594 88312 263600 88324
rect 211672 88284 263600 88312
rect 211672 88272 211678 88284
rect 263594 88272 263600 88284
rect 263652 88272 263658 88324
rect 80054 88204 80060 88256
rect 80112 88244 80118 88256
rect 95142 88244 95148 88256
rect 80112 88216 95148 88244
rect 80112 88204 80118 88216
rect 95142 88204 95148 88216
rect 95200 88204 95206 88256
rect 178770 88204 178776 88256
rect 178828 88244 178834 88256
rect 224954 88244 224960 88256
rect 178828 88216 224960 88244
rect 178828 88204 178834 88216
rect 224954 88204 224960 88216
rect 225012 88204 225018 88256
rect 73798 86912 73804 86964
rect 73856 86952 73862 86964
rect 167730 86952 167736 86964
rect 73856 86924 167736 86952
rect 73856 86912 73862 86924
rect 167730 86912 167736 86924
rect 167788 86952 167794 86964
rect 167788 86924 171134 86952
rect 167788 86912 167794 86924
rect 62022 86844 62028 86896
rect 62080 86884 62086 86896
rect 100018 86884 100024 86896
rect 62080 86856 100024 86884
rect 62080 86844 62086 86856
rect 100018 86844 100024 86856
rect 100076 86844 100082 86896
rect 171106 86884 171134 86924
rect 188430 86912 188436 86964
rect 188488 86952 188494 86964
rect 226518 86952 226524 86964
rect 188488 86924 226524 86952
rect 188488 86912 188494 86924
rect 226518 86912 226524 86924
rect 226576 86912 226582 86964
rect 285766 86912 285772 86964
rect 285824 86952 285830 86964
rect 580166 86952 580172 86964
rect 285824 86924 580172 86952
rect 285824 86912 285830 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 199378 86884 199384 86896
rect 171106 86856 199384 86884
rect 199378 86844 199384 86856
rect 199436 86844 199442 86896
rect 220630 86844 220636 86896
rect 220688 86884 220694 86896
rect 253198 86884 253204 86896
rect 220688 86856 253204 86884
rect 220688 86844 220694 86856
rect 253198 86844 253204 86856
rect 253256 86844 253262 86896
rect 3418 85484 3424 85536
rect 3476 85524 3482 85536
rect 61378 85524 61384 85536
rect 3476 85496 61384 85524
rect 3476 85484 3482 85496
rect 61378 85484 61384 85496
rect 61436 85524 61442 85536
rect 116578 85524 116584 85536
rect 61436 85496 116584 85524
rect 61436 85484 61442 85496
rect 116578 85484 116584 85496
rect 116636 85484 116642 85536
rect 124030 85484 124036 85536
rect 124088 85524 124094 85536
rect 215294 85524 215300 85536
rect 124088 85496 215300 85524
rect 124088 85484 124094 85496
rect 215294 85484 215300 85496
rect 215352 85484 215358 85536
rect 67450 85416 67456 85468
rect 67508 85456 67514 85468
rect 97442 85456 97448 85468
rect 67508 85428 97448 85456
rect 67508 85416 67514 85428
rect 97442 85416 97448 85428
rect 97500 85416 97506 85468
rect 173250 85416 173256 85468
rect 173308 85456 173314 85468
rect 201402 85456 201408 85468
rect 173308 85428 201408 85456
rect 173308 85416 173314 85428
rect 201402 85416 201408 85428
rect 201460 85416 201466 85468
rect 201402 84804 201408 84856
rect 201460 84844 201466 84856
rect 214558 84844 214564 84856
rect 201460 84816 214564 84844
rect 201460 84804 201466 84816
rect 214558 84804 214564 84816
rect 214616 84804 214622 84856
rect 216582 84260 216588 84312
rect 216640 84300 216646 84312
rect 266354 84300 266360 84312
rect 216640 84272 266360 84300
rect 216640 84260 216646 84272
rect 266354 84260 266360 84272
rect 266412 84260 266418 84312
rect 222838 84192 222844 84244
rect 222896 84232 222902 84244
rect 342346 84232 342352 84244
rect 222896 84204 342352 84232
rect 222896 84192 222902 84204
rect 342346 84192 342352 84204
rect 342404 84192 342410 84244
rect 71774 84124 71780 84176
rect 71832 84164 71838 84176
rect 102134 84164 102140 84176
rect 71832 84136 102140 84164
rect 71832 84124 71838 84136
rect 102134 84124 102140 84136
rect 102192 84164 102198 84176
rect 196066 84164 196072 84176
rect 102192 84136 196072 84164
rect 102192 84124 102198 84136
rect 196066 84124 196072 84136
rect 196124 84124 196130 84176
rect 73154 84056 73160 84108
rect 73212 84096 73218 84108
rect 161474 84096 161480 84108
rect 73212 84068 161480 84096
rect 73212 84056 73218 84068
rect 161474 84056 161480 84068
rect 161532 84096 161538 84108
rect 162762 84096 162768 84108
rect 161532 84068 162768 84096
rect 161532 84056 161538 84068
rect 162762 84056 162768 84068
rect 162820 84056 162826 84108
rect 191742 82832 191748 82884
rect 191800 82872 191806 82884
rect 248414 82872 248420 82884
rect 191800 82844 248420 82872
rect 191800 82832 191806 82844
rect 248414 82832 248420 82844
rect 248472 82832 248478 82884
rect 75914 82764 75920 82816
rect 75972 82804 75978 82816
rect 107654 82804 107660 82816
rect 75972 82776 107660 82804
rect 75972 82764 75978 82776
rect 107654 82764 107660 82776
rect 107712 82764 107718 82816
rect 153838 82764 153844 82816
rect 153896 82804 153902 82816
rect 244458 82804 244464 82816
rect 153896 82776 244464 82804
rect 153896 82764 153902 82776
rect 244458 82764 244464 82776
rect 244516 82764 244522 82816
rect 92474 82696 92480 82748
rect 92532 82736 92538 82748
rect 122098 82736 122104 82748
rect 92532 82708 122104 82736
rect 92532 82696 92538 82708
rect 122098 82696 122104 82708
rect 122156 82696 122162 82748
rect 185670 82696 185676 82748
rect 185728 82736 185734 82748
rect 203518 82736 203524 82748
rect 185728 82708 203524 82736
rect 185728 82696 185734 82708
rect 203518 82696 203524 82708
rect 203576 82696 203582 82748
rect 203610 82696 203616 82748
rect 203668 82736 203674 82748
rect 284294 82736 284300 82748
rect 203668 82708 284300 82736
rect 203668 82696 203674 82708
rect 284294 82696 284300 82708
rect 284352 82696 284358 82748
rect 284294 82084 284300 82136
rect 284352 82124 284358 82136
rect 582742 82124 582748 82136
rect 284352 82096 582748 82124
rect 284352 82084 284358 82096
rect 582742 82084 582748 82096
rect 582800 82084 582806 82136
rect 244458 81404 244464 81456
rect 244516 81444 244522 81456
rect 244918 81444 244924 81456
rect 244516 81416 244924 81444
rect 244516 81404 244522 81416
rect 244918 81404 244924 81416
rect 244976 81404 244982 81456
rect 63310 81336 63316 81388
rect 63368 81376 63374 81388
rect 159450 81376 159456 81388
rect 63368 81348 159456 81376
rect 63368 81336 63374 81348
rect 159450 81336 159456 81348
rect 159508 81336 159514 81388
rect 173342 81336 173348 81388
rect 173400 81376 173406 81388
rect 227990 81376 227996 81388
rect 173400 81348 227996 81376
rect 173400 81336 173406 81348
rect 227990 81336 227996 81348
rect 228048 81336 228054 81388
rect 77294 81268 77300 81320
rect 77352 81308 77358 81320
rect 108390 81308 108396 81320
rect 77352 81280 108396 81308
rect 77352 81268 77358 81280
rect 108390 81268 108396 81280
rect 108448 81268 108454 81320
rect 191098 80656 191104 80708
rect 191156 80696 191162 80708
rect 280798 80696 280804 80708
rect 191156 80668 280804 80696
rect 191156 80656 191162 80668
rect 280798 80656 280804 80668
rect 280856 80656 280862 80708
rect 64782 79976 64788 80028
rect 64840 80016 64846 80028
rect 191742 80016 191748 80028
rect 64840 79988 191748 80016
rect 64840 79976 64846 79988
rect 191742 79976 191748 79988
rect 191800 79976 191806 80028
rect 85666 79908 85672 79960
rect 85724 79948 85730 79960
rect 104894 79948 104900 79960
rect 85724 79920 104900 79948
rect 85724 79908 85730 79920
rect 104894 79908 104900 79920
rect 104952 79908 104958 79960
rect 162762 79908 162768 79960
rect 162820 79948 162826 79960
rect 198826 79948 198832 79960
rect 162820 79920 198832 79948
rect 162820 79908 162826 79920
rect 198826 79908 198832 79920
rect 198884 79908 198890 79960
rect 198826 79364 198832 79416
rect 198884 79404 198890 79416
rect 240134 79404 240140 79416
rect 198884 79376 240140 79404
rect 198884 79364 198890 79376
rect 240134 79364 240140 79376
rect 240192 79364 240198 79416
rect 240778 79364 240784 79416
rect 240836 79404 240842 79416
rect 241514 79404 241520 79416
rect 240836 79376 241520 79404
rect 240836 79364 240842 79376
rect 241514 79364 241520 79376
rect 241572 79364 241578 79416
rect 211062 79296 211068 79348
rect 211120 79336 211126 79348
rect 582834 79336 582840 79348
rect 211120 79308 582840 79336
rect 211120 79296 211126 79308
rect 582834 79296 582840 79308
rect 582892 79296 582898 79348
rect 87046 78616 87052 78668
rect 87104 78656 87110 78668
rect 216582 78656 216588 78668
rect 87104 78628 216588 78656
rect 87104 78616 87110 78628
rect 216582 78616 216588 78628
rect 216640 78616 216646 78668
rect 80238 78548 80244 78600
rect 80296 78588 80302 78600
rect 177942 78588 177948 78600
rect 80296 78560 177948 78588
rect 80296 78548 80302 78560
rect 177942 78548 177948 78560
rect 178000 78588 178006 78600
rect 206278 78588 206284 78600
rect 178000 78560 206284 78588
rect 178000 78548 178006 78560
rect 206278 78548 206284 78560
rect 206336 78548 206342 78600
rect 207014 77256 207020 77308
rect 207072 77296 207078 77308
rect 208302 77296 208308 77308
rect 207072 77268 208308 77296
rect 207072 77256 207078 77268
rect 208302 77256 208308 77268
rect 208360 77296 208366 77308
rect 246298 77296 246304 77308
rect 208360 77268 246304 77296
rect 208360 77256 208366 77268
rect 246298 77256 246304 77268
rect 246356 77256 246362 77308
rect 95142 77188 95148 77240
rect 95200 77228 95206 77240
rect 222838 77228 222844 77240
rect 95200 77200 222844 77228
rect 95200 77188 95206 77200
rect 222838 77188 222844 77200
rect 222896 77188 222902 77240
rect 61838 77120 61844 77172
rect 61896 77160 61902 77172
rect 100110 77160 100116 77172
rect 61896 77132 100116 77160
rect 61896 77120 61902 77132
rect 100110 77120 100116 77132
rect 100168 77120 100174 77172
rect 109678 77120 109684 77172
rect 109736 77160 109742 77172
rect 227806 77160 227812 77172
rect 109736 77132 227812 77160
rect 109736 77120 109742 77132
rect 227806 77120 227812 77132
rect 227864 77120 227870 77172
rect 66070 75828 66076 75880
rect 66128 75868 66134 75880
rect 180242 75868 180248 75880
rect 66128 75840 180248 75868
rect 66128 75828 66134 75840
rect 180242 75828 180248 75840
rect 180300 75828 180306 75880
rect 177390 75760 177396 75812
rect 177448 75800 177454 75812
rect 229094 75800 229100 75812
rect 177448 75772 229100 75800
rect 177448 75760 177454 75772
rect 229094 75760 229100 75772
rect 229152 75760 229158 75812
rect 75822 75148 75828 75200
rect 75880 75188 75886 75200
rect 171778 75188 171784 75200
rect 75880 75160 171784 75188
rect 75880 75148 75886 75160
rect 171778 75148 171784 75160
rect 171836 75148 171842 75200
rect 190454 75148 190460 75200
rect 190512 75188 190518 75200
rect 207014 75188 207020 75200
rect 190512 75160 207020 75188
rect 190512 75148 190518 75160
rect 207014 75148 207020 75160
rect 207072 75148 207078 75200
rect 59078 74468 59084 74520
rect 59136 74508 59142 74520
rect 187050 74508 187056 74520
rect 59136 74480 187056 74508
rect 59136 74468 59142 74480
rect 187050 74468 187056 74480
rect 187108 74468 187114 74520
rect 180150 74400 180156 74452
rect 180208 74440 180214 74452
rect 230566 74440 230572 74452
rect 180208 74412 230572 74440
rect 180208 74400 180214 74412
rect 230566 74400 230572 74412
rect 230624 74400 230630 74452
rect 89622 73788 89628 73840
rect 89680 73828 89686 73840
rect 173158 73828 173164 73840
rect 89680 73800 173164 73828
rect 89680 73788 89686 73800
rect 173158 73788 173164 73800
rect 173216 73788 173222 73840
rect 58618 73176 58624 73228
rect 58676 73216 58682 73228
rect 59078 73216 59084 73228
rect 58676 73188 59084 73216
rect 58676 73176 58682 73188
rect 59078 73176 59084 73188
rect 59136 73176 59142 73228
rect 169018 73108 169024 73160
rect 169076 73148 169082 73160
rect 227898 73148 227904 73160
rect 169076 73120 227904 73148
rect 169076 73108 169082 73120
rect 227898 73108 227904 73120
rect 227956 73108 227962 73160
rect 178678 73040 178684 73092
rect 178736 73080 178742 73092
rect 205726 73080 205732 73092
rect 178736 73052 205732 73080
rect 178736 73040 178742 73052
rect 205726 73040 205732 73052
rect 205784 73040 205790 73092
rect 86862 72428 86868 72480
rect 86920 72468 86926 72480
rect 170398 72468 170404 72480
rect 86920 72440 170404 72468
rect 86920 72428 86926 72440
rect 170398 72428 170404 72440
rect 170456 72428 170462 72480
rect 211798 72428 211804 72480
rect 211856 72468 211862 72480
rect 356054 72468 356060 72480
rect 211856 72440 356060 72468
rect 211856 72428 211862 72440
rect 356054 72428 356060 72440
rect 356112 72428 356118 72480
rect 205726 71748 205732 71800
rect 205784 71788 205790 71800
rect 206370 71788 206376 71800
rect 205784 71760 206376 71788
rect 205784 71748 205790 71760
rect 206370 71748 206376 71760
rect 206428 71748 206434 71800
rect 227898 71748 227904 71800
rect 227956 71788 227962 71800
rect 228358 71788 228364 71800
rect 227956 71760 228364 71788
rect 227956 71748 227962 71760
rect 228358 71748 228364 71760
rect 228416 71748 228422 71800
rect 3418 71680 3424 71732
rect 3476 71720 3482 71732
rect 95326 71720 95332 71732
rect 3476 71692 95332 71720
rect 3476 71680 3482 71692
rect 95326 71680 95332 71692
rect 95384 71680 95390 71732
rect 128262 71680 128268 71732
rect 128320 71720 128326 71732
rect 226334 71720 226340 71732
rect 128320 71692 226340 71720
rect 128320 71680 128326 71692
rect 226334 71680 226340 71692
rect 226392 71680 226398 71732
rect 93762 71000 93768 71052
rect 93820 71040 93826 71052
rect 157978 71040 157984 71052
rect 93820 71012 157984 71040
rect 93820 71000 93826 71012
rect 157978 71000 157984 71012
rect 158036 71000 158042 71052
rect 183370 71000 183376 71052
rect 183428 71040 183434 71052
rect 191098 71040 191104 71052
rect 183428 71012 191104 71040
rect 183428 71000 183434 71012
rect 191098 71000 191104 71012
rect 191156 71000 191162 71052
rect 192938 71000 192944 71052
rect 192996 71040 193002 71052
rect 281534 71040 281540 71052
rect 192996 71012 281540 71040
rect 192996 71000 193002 71012
rect 281534 71000 281540 71012
rect 281592 71000 281598 71052
rect 226334 70388 226340 70440
rect 226392 70428 226398 70440
rect 226978 70428 226984 70440
rect 226392 70400 226984 70428
rect 226392 70388 226398 70400
rect 226978 70388 226984 70400
rect 227036 70388 227042 70440
rect 162118 70320 162124 70372
rect 162176 70360 162182 70372
rect 231854 70360 231860 70372
rect 162176 70332 231860 70360
rect 162176 70320 162182 70332
rect 231854 70320 231860 70332
rect 231912 70320 231918 70372
rect 96522 69640 96528 69692
rect 96580 69680 96586 69692
rect 164878 69680 164884 69692
rect 96580 69652 164884 69680
rect 96580 69640 96586 69652
rect 164878 69640 164884 69652
rect 164936 69640 164942 69692
rect 190362 69640 190368 69692
rect 190420 69680 190426 69692
rect 250438 69680 250444 69692
rect 190420 69652 250444 69680
rect 190420 69640 190426 69652
rect 250438 69640 250444 69652
rect 250496 69640 250502 69692
rect 89898 68960 89904 69012
rect 89956 69000 89962 69012
rect 220078 69000 220084 69012
rect 89956 68972 220084 69000
rect 89956 68960 89962 68972
rect 220078 68960 220084 68972
rect 220136 68960 220142 69012
rect 80146 68892 80152 68944
rect 80204 68932 80210 68944
rect 190454 68932 190460 68944
rect 80204 68904 190460 68932
rect 80204 68892 80210 68904
rect 190454 68892 190460 68904
rect 190512 68892 190518 68944
rect 193122 68280 193128 68332
rect 193180 68320 193186 68332
rect 327074 68320 327080 68332
rect 193180 68292 327080 68320
rect 193180 68280 193186 68292
rect 327074 68280 327080 68292
rect 327132 68280 327138 68332
rect 91002 67532 91008 67584
rect 91060 67572 91066 67584
rect 218054 67572 218060 67584
rect 91060 67544 218060 67572
rect 91060 67532 91066 67544
rect 218054 67532 218060 67544
rect 218112 67532 218118 67584
rect 67542 66852 67548 66904
rect 67600 66892 67606 66904
rect 99926 66892 99932 66904
rect 67600 66864 99932 66892
rect 67600 66852 67606 66864
rect 99926 66852 99932 66864
rect 99984 66852 99990 66904
rect 81434 66172 81440 66224
rect 81492 66212 81498 66224
rect 208486 66212 208492 66224
rect 81492 66184 208492 66212
rect 81492 66172 81498 66184
rect 208486 66172 208492 66184
rect 208544 66212 208550 66224
rect 209038 66212 209044 66224
rect 208544 66184 209044 66212
rect 208544 66172 208550 66184
rect 209038 66172 209044 66184
rect 209096 66172 209102 66224
rect 86954 66104 86960 66156
rect 87012 66144 87018 66156
rect 115934 66144 115940 66156
rect 87012 66116 115940 66144
rect 87012 66104 87018 66116
rect 115934 66104 115940 66116
rect 115992 66144 115998 66156
rect 215938 66144 215944 66156
rect 115992 66116 215944 66144
rect 115992 66104 115998 66116
rect 215938 66104 215944 66116
rect 215996 66104 216002 66156
rect 93670 64812 93676 64864
rect 93728 64852 93734 64864
rect 241606 64852 241612 64864
rect 93728 64824 241612 64852
rect 93728 64812 93734 64824
rect 241606 64812 241612 64824
rect 241664 64812 241670 64864
rect 74534 64744 74540 64796
rect 74592 64784 74598 64796
rect 201494 64784 201500 64796
rect 74592 64756 201500 64784
rect 74592 64744 74598 64756
rect 201494 64744 201500 64756
rect 201552 64744 201558 64796
rect 201494 63520 201500 63572
rect 201552 63560 201558 63572
rect 202138 63560 202144 63572
rect 201552 63532 202144 63560
rect 201552 63520 201558 63532
rect 202138 63520 202144 63532
rect 202196 63520 202202 63572
rect 241606 63520 241612 63572
rect 241664 63560 241670 63572
rect 242158 63560 242164 63572
rect 241664 63532 242164 63560
rect 241664 63520 241670 63532
rect 242158 63520 242164 63532
rect 242216 63520 242222 63572
rect 71866 63452 71872 63504
rect 71924 63492 71930 63504
rect 197998 63492 198004 63504
rect 71924 63464 198004 63492
rect 71924 63452 71930 63464
rect 197998 63452 198004 63464
rect 198056 63452 198062 63504
rect 218054 63452 218060 63504
rect 218112 63492 218118 63504
rect 277394 63492 277400 63504
rect 218112 63464 277400 63492
rect 218112 63452 218118 63464
rect 277394 63452 277400 63464
rect 277452 63492 277458 63504
rect 278682 63492 278688 63504
rect 277452 63464 278688 63492
rect 277452 63452 277458 63464
rect 278682 63452 278688 63464
rect 278740 63452 278746 63504
rect 278682 62772 278688 62824
rect 278740 62812 278746 62824
rect 351914 62812 351920 62824
rect 278740 62784 351920 62812
rect 278740 62772 278746 62784
rect 351914 62772 351920 62784
rect 351972 62772 351978 62824
rect 85574 62024 85580 62076
rect 85632 62064 85638 62076
rect 212626 62064 212632 62076
rect 85632 62036 212632 62064
rect 85632 62024 85638 62036
rect 212626 62024 212632 62036
rect 212684 62024 212690 62076
rect 212626 60732 212632 60784
rect 212684 60772 212690 60784
rect 213270 60772 213276 60784
rect 212684 60744 213276 60772
rect 212684 60732 212690 60744
rect 213270 60732 213276 60744
rect 213328 60732 213334 60784
rect 88334 60664 88340 60716
rect 88392 60704 88398 60716
rect 222378 60704 222384 60716
rect 88392 60676 222384 60704
rect 88392 60664 88398 60676
rect 222378 60664 222384 60676
rect 222436 60704 222442 60716
rect 222930 60704 222936 60716
rect 222436 60676 222936 60704
rect 222436 60664 222442 60676
rect 222930 60664 222936 60676
rect 222988 60664 222994 60716
rect 193858 59984 193864 60036
rect 193916 60024 193922 60036
rect 264974 60024 264980 60036
rect 193916 59996 264980 60024
rect 193916 59984 193922 59996
rect 264974 59984 264980 59996
rect 265032 59984 265038 60036
rect 99926 59304 99932 59356
rect 99984 59344 99990 59356
rect 193306 59344 193312 59356
rect 99984 59316 193312 59344
rect 99984 59304 99990 59316
rect 193306 59304 193312 59316
rect 193364 59344 193370 59356
rect 193858 59344 193864 59356
rect 193364 59316 193864 59344
rect 193364 59304 193370 59316
rect 193858 59304 193864 59316
rect 193916 59304 193922 59356
rect 57882 58624 57888 58676
rect 57940 58664 57946 58676
rect 181438 58664 181444 58676
rect 57940 58636 181444 58664
rect 57940 58624 57946 58636
rect 181438 58624 181444 58636
rect 181496 58624 181502 58676
rect 82078 57876 82084 57928
rect 82136 57916 82142 57928
rect 210418 57916 210424 57928
rect 82136 57888 210424 57916
rect 82136 57876 82142 57888
rect 210418 57876 210424 57888
rect 210476 57876 210482 57928
rect 84194 57808 84200 57860
rect 84252 57848 84258 57860
rect 118694 57848 118700 57860
rect 84252 57820 118700 57848
rect 84252 57808 84258 57820
rect 118694 57808 118700 57820
rect 118752 57848 118758 57860
rect 213178 57848 213184 57860
rect 118752 57820 213184 57848
rect 118752 57808 118758 57820
rect 213178 57808 213184 57820
rect 213236 57808 213242 57860
rect 73798 56516 73804 56568
rect 73856 56556 73862 56568
rect 200114 56556 200120 56568
rect 73856 56528 200120 56556
rect 73856 56516 73862 56528
rect 200114 56516 200120 56528
rect 200172 56556 200178 56568
rect 200758 56556 200764 56568
rect 200172 56528 200764 56556
rect 200172 56516 200178 56528
rect 200758 56516 200764 56528
rect 200816 56516 200822 56568
rect 77202 54476 77208 54528
rect 77260 54516 77266 54528
rect 152550 54516 152556 54528
rect 77260 54488 152556 54516
rect 77260 54476 77266 54488
rect 152550 54476 152556 54488
rect 152608 54476 152614 54528
rect 193858 54476 193864 54528
rect 193916 54516 193922 54528
rect 291194 54516 291200 54528
rect 193916 54488 291200 54516
rect 193916 54476 193922 54488
rect 291194 54476 291200 54488
rect 291252 54476 291258 54528
rect 101398 53048 101404 53100
rect 101456 53088 101462 53100
rect 137370 53088 137376 53100
rect 101456 53060 137376 53088
rect 101456 53048 101462 53060
rect 137370 53048 137376 53060
rect 137428 53048 137434 53100
rect 184842 53048 184848 53100
rect 184900 53088 184906 53100
rect 292666 53088 292672 53100
rect 184900 53060 292672 53088
rect 184900 53048 184906 53060
rect 292666 53048 292672 53060
rect 292724 53048 292730 53100
rect 186130 51688 186136 51740
rect 186188 51728 186194 51740
rect 328454 51728 328460 51740
rect 186188 51700 328460 51728
rect 186188 51688 186194 51700
rect 328454 51688 328460 51700
rect 328512 51688 328518 51740
rect 55122 50328 55128 50380
rect 55180 50368 55186 50380
rect 141510 50368 141516 50380
rect 55180 50340 141516 50368
rect 55180 50328 55186 50340
rect 141510 50328 141516 50340
rect 141568 50328 141574 50380
rect 180242 50328 180248 50380
rect 180300 50368 180306 50380
rect 269114 50368 269120 50380
rect 180300 50340 269120 50368
rect 180300 50328 180306 50340
rect 269114 50328 269120 50340
rect 269172 50328 269178 50380
rect 73062 48968 73068 49020
rect 73120 49008 73126 49020
rect 149698 49008 149704 49020
rect 73120 48980 149704 49008
rect 73120 48968 73126 48980
rect 149698 48968 149704 48980
rect 149756 48968 149762 49020
rect 188982 48968 188988 49020
rect 189040 49008 189046 49020
rect 251266 49008 251272 49020
rect 189040 48980 251272 49008
rect 189040 48968 189046 48980
rect 251266 48968 251272 48980
rect 251324 48968 251330 49020
rect 68922 47540 68928 47592
rect 68980 47580 68986 47592
rect 175918 47580 175924 47592
rect 68980 47552 175924 47580
rect 68980 47540 68986 47552
rect 175918 47540 175924 47552
rect 175976 47540 175982 47592
rect 204898 47540 204904 47592
rect 204956 47580 204962 47592
rect 343634 47580 343640 47592
rect 204956 47552 343640 47580
rect 204956 47540 204962 47552
rect 343634 47540 343640 47552
rect 343692 47540 343698 47592
rect 189718 46860 189724 46912
rect 189776 46900 189782 46912
rect 580166 46900 580172 46912
rect 189776 46872 580172 46900
rect 189776 46860 189782 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 3418 45500 3424 45552
rect 3476 45540 3482 45552
rect 57238 45540 57244 45552
rect 3476 45512 57244 45540
rect 3476 45500 3482 45512
rect 57238 45500 57244 45512
rect 57296 45500 57302 45552
rect 59262 44820 59268 44872
rect 59320 44860 59326 44872
rect 144178 44860 144184 44872
rect 59320 44832 144184 44860
rect 59320 44820 59326 44832
rect 144178 44820 144184 44832
rect 144236 44820 144242 44872
rect 171042 44820 171048 44872
rect 171100 44860 171106 44872
rect 332686 44860 332692 44872
rect 171100 44832 332692 44860
rect 171100 44820 171106 44832
rect 332686 44820 332692 44832
rect 332744 44820 332750 44872
rect 181530 43392 181536 43444
rect 181588 43432 181594 43444
rect 222838 43432 222844 43444
rect 181588 43404 222844 43432
rect 181588 43392 181594 43404
rect 222838 43392 222844 43404
rect 222896 43392 222902 43444
rect 226978 43392 226984 43444
rect 227036 43432 227042 43444
rect 277394 43432 277400 43444
rect 227036 43404 277400 43432
rect 227036 43392 227042 43404
rect 277394 43392 277400 43404
rect 277452 43392 277458 43444
rect 61930 42032 61936 42084
rect 61988 42072 61994 42084
rect 138658 42072 138664 42084
rect 61988 42044 138664 42072
rect 61988 42032 61994 42044
rect 138658 42032 138664 42044
rect 138716 42032 138722 42084
rect 222930 42032 222936 42084
rect 222988 42072 222994 42084
rect 290458 42072 290464 42084
rect 222988 42044 290464 42072
rect 222988 42032 222994 42044
rect 290458 42032 290464 42044
rect 290516 42032 290522 42084
rect 186958 40672 186964 40724
rect 187016 40712 187022 40724
rect 338114 40712 338120 40724
rect 187016 40684 338120 40712
rect 187016 40672 187022 40684
rect 338114 40672 338120 40684
rect 338172 40672 338178 40724
rect 46842 39312 46848 39364
rect 46900 39352 46906 39364
rect 163498 39352 163504 39364
rect 46900 39324 163504 39352
rect 46900 39312 46906 39324
rect 163498 39312 163504 39324
rect 163556 39312 163562 39364
rect 206370 38020 206376 38072
rect 206428 38060 206434 38072
rect 213362 38060 213368 38072
rect 206428 38032 213368 38060
rect 206428 38020 206434 38032
rect 213362 38020 213368 38032
rect 213420 38020 213426 38072
rect 213178 37884 213184 37936
rect 213236 37924 213242 37936
rect 333974 37924 333980 37936
rect 213236 37896 333980 37924
rect 213236 37884 213242 37896
rect 333974 37884 333980 37896
rect 334032 37884 334038 37936
rect 66162 36524 66168 36576
rect 66220 36564 66226 36576
rect 140038 36564 140044 36576
rect 66220 36536 140044 36564
rect 66220 36524 66226 36536
rect 140038 36524 140044 36536
rect 140096 36524 140102 36576
rect 203518 36524 203524 36576
rect 203576 36564 203582 36576
rect 324406 36564 324412 36576
rect 203576 36536 324412 36564
rect 203576 36524 203582 36536
rect 324406 36524 324412 36536
rect 324464 36524 324470 36576
rect 213270 35164 213276 35216
rect 213328 35204 213334 35216
rect 287054 35204 287060 35216
rect 213328 35176 287060 35204
rect 213328 35164 213334 35176
rect 287054 35164 287060 35176
rect 287112 35164 287118 35216
rect 67726 33736 67732 33788
rect 67784 33776 67790 33788
rect 125594 33776 125600 33788
rect 67784 33748 125600 33776
rect 67784 33736 67790 33748
rect 125594 33736 125600 33748
rect 125652 33736 125658 33788
rect 193030 33736 193036 33788
rect 193088 33776 193094 33788
rect 270494 33776 270500 33788
rect 193088 33748 270500 33776
rect 193088 33736 193094 33748
rect 270494 33736 270500 33748
rect 270552 33736 270558 33788
rect 2866 33056 2872 33108
rect 2924 33096 2930 33108
rect 54478 33096 54484 33108
rect 2924 33068 54484 33096
rect 2924 33056 2930 33068
rect 54478 33056 54484 33068
rect 54536 33056 54542 33108
rect 200758 32376 200764 32428
rect 200816 32416 200822 32428
rect 340966 32416 340972 32428
rect 200816 32388 340972 32416
rect 200816 32376 200822 32388
rect 340966 32376 340972 32388
rect 341024 32376 341030 32428
rect 79962 31016 79968 31068
rect 80020 31056 80026 31068
rect 151078 31056 151084 31068
rect 80020 31028 151084 31056
rect 80020 31016 80026 31028
rect 151078 31016 151084 31028
rect 151136 31016 151142 31068
rect 210418 31016 210424 31068
rect 210476 31056 210482 31068
rect 322934 31056 322940 31068
rect 210476 31028 322940 31056
rect 210476 31016 210482 31028
rect 322934 31016 322940 31028
rect 322992 31016 322998 31068
rect 53742 29588 53748 29640
rect 53800 29628 53806 29640
rect 145558 29628 145564 29640
rect 53800 29600 145564 29628
rect 53800 29588 53806 29600
rect 145558 29588 145564 29600
rect 145616 29588 145622 29640
rect 183462 29588 183468 29640
rect 183520 29628 183526 29640
rect 249794 29628 249800 29640
rect 183520 29600 249800 29628
rect 183520 29588 183526 29600
rect 249794 29588 249800 29600
rect 249852 29588 249858 29640
rect 70302 28228 70308 28280
rect 70360 28268 70366 28280
rect 142890 28268 142896 28280
rect 70360 28240 142896 28268
rect 70360 28228 70366 28240
rect 142890 28228 142896 28240
rect 142948 28228 142954 28280
rect 199378 28228 199384 28280
rect 199436 28268 199442 28280
rect 244274 28268 244280 28280
rect 199436 28240 244280 28268
rect 199436 28228 199442 28240
rect 244274 28228 244280 28240
rect 244332 28228 244338 28280
rect 250438 28228 250444 28280
rect 250496 28268 250502 28280
rect 288434 28268 288440 28280
rect 250496 28240 288440 28268
rect 250496 28228 250502 28240
rect 288434 28228 288440 28240
rect 288492 28228 288498 28280
rect 86770 26868 86776 26920
rect 86828 26908 86834 26920
rect 167638 26908 167644 26920
rect 86828 26880 167644 26908
rect 86828 26868 86834 26880
rect 167638 26868 167644 26880
rect 167696 26868 167702 26920
rect 243538 26868 243544 26920
rect 243596 26908 243602 26920
rect 259546 26908 259552 26920
rect 243596 26880 259552 26908
rect 243596 26868 243602 26880
rect 259546 26868 259552 26880
rect 259604 26868 259610 26920
rect 84102 25508 84108 25560
rect 84160 25548 84166 25560
rect 147030 25548 147036 25560
rect 84160 25520 147036 25548
rect 84160 25508 84166 25520
rect 147030 25508 147036 25520
rect 147088 25508 147094 25560
rect 39942 24080 39948 24132
rect 40000 24120 40006 24132
rect 170490 24120 170496 24132
rect 40000 24092 170496 24120
rect 40000 24080 40006 24092
rect 170490 24080 170496 24092
rect 170548 24080 170554 24132
rect 121362 22720 121368 22772
rect 121420 22760 121426 22772
rect 126238 22760 126244 22772
rect 121420 22732 126244 22760
rect 121420 22720 121426 22732
rect 126238 22720 126244 22732
rect 126296 22720 126302 22772
rect 202138 22720 202144 22772
rect 202196 22760 202202 22772
rect 321554 22760 321560 22772
rect 202196 22732 321560 22760
rect 202196 22720 202202 22732
rect 321554 22720 321560 22732
rect 321612 22720 321618 22772
rect 91002 21360 91008 21412
rect 91060 21400 91066 21412
rect 146938 21400 146944 21412
rect 91060 21372 146944 21400
rect 91060 21360 91066 21372
rect 146938 21360 146944 21372
rect 146996 21360 147002 21412
rect 191098 21360 191104 21412
rect 191156 21400 191162 21412
rect 307754 21400 307760 21412
rect 191156 21372 307760 21400
rect 191156 21360 191162 21372
rect 307754 21360 307760 21372
rect 307812 21360 307818 21412
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 69658 20652 69664 20664
rect 3476 20624 69664 20652
rect 3476 20612 3482 20624
rect 69658 20612 69664 20624
rect 69716 20612 69722 20664
rect 100662 19932 100668 19984
rect 100720 19972 100726 19984
rect 166258 19972 166264 19984
rect 100720 19944 166264 19972
rect 100720 19932 100726 19944
rect 166258 19932 166264 19944
rect 166316 19932 166322 19984
rect 204990 19932 204996 19984
rect 205048 19972 205054 19984
rect 320266 19972 320272 19984
rect 205048 19944 320272 19972
rect 205048 19932 205054 19944
rect 320266 19932 320272 19944
rect 320324 19932 320330 19984
rect 78582 18572 78588 18624
rect 78640 18612 78646 18624
rect 177298 18612 177304 18624
rect 78640 18584 177304 18612
rect 78640 18572 78646 18584
rect 177298 18572 177304 18584
rect 177356 18572 177362 18624
rect 215938 18572 215944 18624
rect 215996 18612 216002 18624
rect 284386 18612 284392 18624
rect 215996 18584 284392 18612
rect 215996 18572 216002 18584
rect 284386 18572 284392 18584
rect 284444 18572 284450 18624
rect 271138 16192 271144 16244
rect 271196 16232 271202 16244
rect 276106 16232 276112 16244
rect 271196 16204 276112 16232
rect 271196 16192 271202 16204
rect 276106 16192 276112 16204
rect 276164 16192 276170 16244
rect 244918 15852 244924 15904
rect 244976 15892 244982 15904
rect 261754 15892 261760 15904
rect 244976 15864 261760 15892
rect 244976 15852 244982 15864
rect 261754 15852 261760 15864
rect 261812 15852 261818 15904
rect 106182 13064 106188 13116
rect 106240 13104 106246 13116
rect 141418 13104 141424 13116
rect 106240 13076 141424 13104
rect 106240 13064 106246 13076
rect 141418 13064 141424 13076
rect 141476 13064 141482 13116
rect 206278 13064 206284 13116
rect 206336 13104 206342 13116
rect 274818 13104 274824 13116
rect 206336 13076 274824 13104
rect 206336 13064 206342 13076
rect 274818 13064 274824 13076
rect 274876 13064 274882 13116
rect 284938 13064 284944 13116
rect 284996 13104 285002 13116
rect 330386 13104 330392 13116
rect 284996 13076 330392 13104
rect 284996 13064 285002 13076
rect 330386 13064 330392 13076
rect 330444 13064 330450 13116
rect 95050 11704 95056 11756
rect 95108 11744 95114 11756
rect 134518 11744 134524 11756
rect 95108 11716 134524 11744
rect 95108 11704 95114 11716
rect 134518 11704 134524 11716
rect 134576 11704 134582 11756
rect 195238 11704 195244 11756
rect 195296 11744 195302 11756
rect 312170 11744 312176 11756
rect 195296 11716 312176 11744
rect 195296 11704 195302 11716
rect 312170 11704 312176 11716
rect 312228 11704 312234 11756
rect 332686 11704 332692 11756
rect 332744 11744 332750 11756
rect 333882 11744 333888 11756
rect 332744 11716 333888 11744
rect 332744 11704 332750 11716
rect 333882 11704 333888 11716
rect 333940 11704 333946 11756
rect 197998 10276 198004 10328
rect 198056 10316 198062 10328
rect 342254 10316 342260 10328
rect 198056 10288 342260 10316
rect 198056 10276 198062 10288
rect 342254 10276 342260 10288
rect 342312 10276 342318 10328
rect 278038 8984 278044 9036
rect 278096 9024 278102 9036
rect 315022 9024 315028 9036
rect 278096 8996 315028 9024
rect 278096 8984 278102 8996
rect 315022 8984 315028 8996
rect 315080 8984 315086 9036
rect 209038 8916 209044 8968
rect 209096 8956 209102 8968
rect 279510 8956 279516 8968
rect 209096 8928 279516 8956
rect 209096 8916 209102 8928
rect 279510 8916 279516 8928
rect 279568 8916 279574 8968
rect 141142 7624 141148 7676
rect 141200 7664 141206 7676
rect 180058 7664 180064 7676
rect 141200 7636 180064 7664
rect 141200 7624 141206 7636
rect 180058 7624 180064 7636
rect 180116 7624 180122 7676
rect 224862 7624 224868 7676
rect 224920 7664 224926 7676
rect 254670 7664 254676 7676
rect 224920 7636 254676 7664
rect 224920 7624 224926 7636
rect 254670 7624 254676 7636
rect 254728 7624 254734 7676
rect 566 7556 572 7608
rect 624 7596 630 7608
rect 97258 7596 97264 7608
rect 624 7568 97264 7596
rect 624 7556 630 7568
rect 97258 7556 97264 7568
rect 97316 7556 97322 7608
rect 97442 7556 97448 7608
rect 97500 7596 97506 7608
rect 142798 7596 142804 7608
rect 97500 7568 142804 7596
rect 97500 7556 97506 7568
rect 142798 7556 142804 7568
rect 142856 7556 142862 7608
rect 195974 7556 195980 7608
rect 196032 7596 196038 7608
rect 258258 7596 258264 7608
rect 196032 7568 258264 7596
rect 196032 7556 196038 7568
rect 258258 7556 258264 7568
rect 258316 7556 258322 7608
rect 269758 7556 269764 7608
rect 269816 7596 269822 7608
rect 317322 7596 317328 7608
rect 269816 7568 317328 7596
rect 269816 7556 269822 7568
rect 317322 7556 317328 7568
rect 317380 7556 317386 7608
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 58618 6848 58624 6860
rect 3476 6820 58624 6848
rect 3476 6808 3482 6820
rect 58618 6808 58624 6820
rect 58676 6808 58682 6860
rect 222838 6196 222844 6248
rect 222896 6236 222902 6248
rect 244090 6236 244096 6248
rect 222896 6208 244096 6236
rect 222896 6196 222902 6208
rect 244090 6196 244096 6208
rect 244148 6196 244154 6248
rect 298738 6196 298744 6248
rect 298796 6236 298802 6248
rect 310238 6236 310244 6248
rect 298796 6208 310244 6236
rect 298796 6196 298802 6208
rect 310238 6196 310244 6208
rect 310296 6196 310302 6248
rect 56042 6128 56048 6180
rect 56100 6168 56106 6180
rect 159358 6168 159364 6180
rect 56100 6140 159364 6168
rect 56100 6128 56106 6140
rect 159358 6128 159364 6140
rect 159416 6128 159422 6180
rect 242158 6128 242164 6180
rect 242216 6168 242222 6180
rect 303154 6168 303160 6180
rect 242216 6140 303160 6168
rect 242216 6128 242222 6140
rect 303154 6128 303160 6140
rect 303212 6128 303218 6180
rect 309778 5516 309784 5568
rect 309836 5556 309842 5568
rect 311434 5556 311440 5568
rect 309836 5528 311440 5556
rect 309836 5516 309842 5528
rect 311434 5516 311440 5528
rect 311492 5516 311498 5568
rect 348050 5516 348056 5568
rect 348108 5556 348114 5568
rect 349154 5556 349160 5568
rect 348108 5528 349160 5556
rect 348108 5516 348114 5528
rect 349154 5516 349160 5528
rect 349212 5516 349218 5568
rect 130378 4768 130384 4820
rect 130436 4808 130442 4820
rect 136450 4808 136456 4820
rect 130436 4780 136456 4808
rect 130436 4768 130442 4780
rect 136450 4768 136456 4780
rect 136508 4768 136514 4820
rect 228358 4768 228364 4820
rect 228416 4808 228422 4820
rect 239306 4808 239312 4820
rect 228416 4780 239312 4808
rect 228416 4768 228422 4780
rect 239306 4768 239312 4780
rect 239364 4768 239370 4820
rect 304258 4768 304264 4820
rect 304316 4808 304322 4820
rect 307938 4808 307944 4820
rect 304316 4780 307944 4808
rect 304316 4768 304322 4780
rect 307938 4768 307944 4780
rect 307996 4768 308002 4820
rect 323578 4768 323584 4820
rect 323636 4808 323642 4820
rect 337470 4808 337476 4820
rect 323636 4780 337476 4808
rect 323636 4768 323642 4780
rect 337470 4768 337476 4780
rect 337528 4768 337534 4820
rect 291838 4428 291844 4480
rect 291896 4468 291902 4480
rect 297266 4468 297272 4480
rect 291896 4440 297272 4468
rect 291896 4428 291902 4440
rect 297266 4428 297272 4440
rect 297324 4428 297330 4480
rect 346946 4156 346952 4208
rect 347004 4196 347010 4208
rect 353294 4196 353300 4208
rect 347004 4168 353300 4196
rect 347004 4156 347010 4168
rect 353294 4156 353300 4168
rect 353352 4156 353358 4208
rect 6822 4088 6828 4140
rect 6880 4128 6886 4140
rect 7650 4128 7656 4140
rect 6880 4100 7656 4128
rect 6880 4088 6886 4100
rect 7650 4088 7656 4100
rect 7708 4088 7714 4140
rect 351638 4088 351644 4140
rect 351696 4128 351702 4140
rect 356054 4128 356060 4140
rect 351696 4100 356060 4128
rect 351696 4088 351702 4100
rect 356054 4088 356060 4100
rect 356112 4088 356118 4140
rect 322198 3952 322204 4004
rect 322256 3992 322262 4004
rect 326798 3992 326804 4004
rect 322256 3964 326804 3992
rect 322256 3952 322262 3964
rect 326798 3952 326804 3964
rect 326856 3952 326862 4004
rect 1302 3544 1308 3596
rect 1360 3584 1366 3596
rect 2866 3584 2872 3596
rect 1360 3556 2872 3584
rect 1360 3544 1366 3556
rect 2866 3544 2872 3556
rect 2924 3544 2930 3596
rect 52546 3544 52552 3596
rect 52604 3584 52610 3596
rect 53650 3584 53656 3596
rect 52604 3556 53656 3584
rect 52604 3544 52610 3556
rect 53650 3544 53656 3556
rect 53708 3544 53714 3596
rect 60826 3544 60832 3596
rect 60884 3584 60890 3596
rect 61930 3584 61936 3596
rect 60884 3556 61936 3584
rect 60884 3544 60890 3556
rect 61930 3544 61936 3556
rect 61988 3544 61994 3596
rect 69106 3544 69112 3596
rect 69164 3584 69170 3596
rect 70210 3584 70216 3596
rect 69164 3556 70216 3584
rect 69164 3544 69170 3556
rect 70210 3544 70216 3556
rect 70268 3544 70274 3596
rect 80882 3544 80888 3596
rect 80940 3584 80946 3596
rect 83458 3584 83464 3596
rect 80940 3556 83464 3584
rect 80940 3544 80946 3556
rect 83458 3544 83464 3556
rect 83516 3544 83522 3596
rect 105722 3544 105728 3596
rect 105780 3584 105786 3596
rect 106182 3584 106188 3596
rect 105780 3556 106188 3584
rect 105780 3544 105786 3556
rect 106182 3544 106188 3556
rect 106240 3544 106246 3596
rect 122282 3544 122288 3596
rect 122340 3584 122346 3596
rect 122742 3584 122748 3596
rect 122340 3556 122748 3584
rect 122340 3544 122346 3556
rect 122742 3544 122748 3556
rect 122800 3544 122806 3596
rect 123478 3544 123484 3596
rect 123536 3584 123542 3596
rect 124122 3584 124128 3596
rect 123536 3556 124128 3584
rect 123536 3544 123542 3556
rect 124122 3544 124128 3556
rect 124180 3544 124186 3596
rect 124674 3544 124680 3596
rect 124732 3584 124738 3596
rect 125502 3584 125508 3596
rect 124732 3556 125508 3584
rect 124732 3544 124738 3556
rect 125502 3544 125508 3556
rect 125560 3544 125566 3596
rect 251174 3544 251180 3596
rect 251232 3584 251238 3596
rect 252370 3584 252376 3596
rect 251232 3556 252376 3584
rect 251232 3544 251238 3556
rect 252370 3544 252376 3556
rect 252428 3544 252434 3596
rect 276014 3544 276020 3596
rect 276072 3584 276078 3596
rect 277118 3584 277124 3596
rect 276072 3556 277124 3584
rect 276072 3544 276078 3556
rect 277118 3544 277124 3556
rect 277176 3544 277182 3596
rect 1670 3476 1676 3528
rect 1728 3516 1734 3528
rect 2682 3516 2688 3528
rect 1728 3488 2688 3516
rect 1728 3476 1734 3488
rect 2682 3476 2688 3488
rect 2740 3476 2746 3528
rect 9950 3476 9956 3528
rect 10008 3516 10014 3528
rect 10962 3516 10968 3528
rect 10008 3488 10968 3516
rect 10008 3476 10014 3488
rect 10962 3476 10968 3488
rect 11020 3476 11026 3528
rect 11146 3476 11152 3528
rect 11204 3516 11210 3528
rect 12250 3516 12256 3528
rect 11204 3488 12256 3516
rect 11204 3476 11210 3488
rect 12250 3476 12256 3488
rect 12308 3476 12314 3528
rect 17034 3476 17040 3528
rect 17092 3516 17098 3528
rect 17862 3516 17868 3528
rect 17092 3488 17868 3516
rect 17092 3476 17098 3488
rect 17862 3476 17868 3488
rect 17920 3476 17926 3528
rect 18230 3476 18236 3528
rect 18288 3516 18294 3528
rect 19242 3516 19248 3528
rect 18288 3488 19248 3516
rect 18288 3476 18294 3488
rect 19242 3476 19248 3488
rect 19300 3476 19306 3528
rect 20622 3476 20628 3528
rect 20680 3516 20686 3528
rect 21358 3516 21364 3528
rect 20680 3488 21364 3516
rect 20680 3476 20686 3488
rect 21358 3476 21364 3488
rect 21416 3476 21422 3528
rect 24210 3476 24216 3528
rect 24268 3516 24274 3528
rect 24762 3516 24768 3528
rect 24268 3488 24768 3516
rect 24268 3476 24274 3488
rect 24762 3476 24768 3488
rect 24820 3476 24826 3528
rect 26510 3476 26516 3528
rect 26568 3516 26574 3528
rect 27522 3516 27528 3528
rect 26568 3488 27528 3516
rect 26568 3476 26574 3488
rect 27522 3476 27528 3488
rect 27580 3476 27586 3528
rect 32398 3476 32404 3528
rect 32456 3516 32462 3528
rect 33042 3516 33048 3528
rect 32456 3488 33048 3516
rect 32456 3476 32462 3488
rect 33042 3476 33048 3488
rect 33100 3476 33106 3528
rect 33594 3476 33600 3528
rect 33652 3516 33658 3528
rect 34422 3516 34428 3528
rect 33652 3488 34428 3516
rect 33652 3476 33658 3488
rect 34422 3476 34428 3488
rect 34480 3476 34486 3528
rect 34790 3476 34796 3528
rect 34848 3516 34854 3528
rect 35802 3516 35808 3528
rect 34848 3488 35808 3516
rect 34848 3476 34854 3488
rect 35802 3476 35808 3488
rect 35860 3476 35866 3528
rect 35986 3476 35992 3528
rect 36044 3516 36050 3528
rect 37090 3516 37096 3528
rect 36044 3488 37096 3516
rect 36044 3476 36050 3488
rect 37090 3476 37096 3488
rect 37148 3476 37154 3528
rect 40678 3476 40684 3528
rect 40736 3516 40742 3528
rect 41322 3516 41328 3528
rect 40736 3488 41328 3516
rect 40736 3476 40742 3488
rect 41322 3476 41328 3488
rect 41380 3476 41386 3528
rect 41874 3476 41880 3528
rect 41932 3516 41938 3528
rect 42702 3516 42708 3528
rect 41932 3488 42708 3516
rect 41932 3476 41938 3488
rect 42702 3476 42708 3488
rect 42760 3476 42766 3528
rect 43070 3476 43076 3528
rect 43128 3516 43134 3528
rect 44082 3516 44088 3528
rect 43128 3488 44088 3516
rect 43128 3476 43134 3488
rect 44082 3476 44088 3488
rect 44140 3476 44146 3528
rect 44266 3476 44272 3528
rect 44324 3516 44330 3528
rect 45370 3516 45376 3528
rect 44324 3488 45376 3516
rect 44324 3476 44330 3488
rect 45370 3476 45376 3488
rect 45428 3476 45434 3528
rect 48958 3476 48964 3528
rect 49016 3516 49022 3528
rect 49510 3516 49516 3528
rect 49016 3488 49516 3516
rect 49016 3476 49022 3488
rect 49510 3476 49516 3488
rect 49568 3476 49574 3528
rect 50154 3476 50160 3528
rect 50212 3516 50218 3528
rect 50890 3516 50896 3528
rect 50212 3488 50896 3516
rect 50212 3476 50218 3488
rect 50890 3476 50896 3488
rect 50948 3476 50954 3528
rect 57238 3476 57244 3528
rect 57296 3516 57302 3528
rect 57882 3516 57888 3528
rect 57296 3488 57888 3516
rect 57296 3476 57302 3488
rect 57882 3476 57888 3488
rect 57940 3476 57946 3528
rect 58434 3476 58440 3528
rect 58492 3516 58498 3528
rect 59262 3516 59268 3528
rect 58492 3488 59268 3516
rect 58492 3476 58498 3488
rect 59262 3476 59268 3488
rect 59320 3476 59326 3528
rect 59630 3476 59636 3528
rect 59688 3516 59694 3528
rect 60642 3516 60648 3528
rect 59688 3488 60648 3516
rect 59688 3476 59694 3488
rect 60642 3476 60648 3488
rect 60700 3476 60706 3528
rect 64322 3476 64328 3528
rect 64380 3516 64386 3528
rect 64782 3516 64788 3528
rect 64380 3488 64788 3516
rect 64380 3476 64386 3488
rect 64782 3476 64788 3488
rect 64840 3476 64846 3528
rect 65518 3476 65524 3528
rect 65576 3516 65582 3528
rect 66162 3516 66168 3528
rect 65576 3488 66168 3516
rect 65576 3476 65582 3488
rect 66162 3476 66168 3488
rect 66220 3476 66226 3528
rect 67910 3476 67916 3528
rect 67968 3516 67974 3528
rect 68922 3516 68928 3528
rect 67968 3488 68928 3516
rect 67968 3476 67974 3488
rect 68922 3476 68928 3488
rect 68980 3476 68986 3528
rect 72602 3476 72608 3528
rect 72660 3516 72666 3528
rect 73062 3516 73068 3528
rect 72660 3488 73068 3516
rect 72660 3476 72666 3488
rect 73062 3476 73068 3488
rect 73120 3476 73126 3528
rect 74994 3476 75000 3528
rect 75052 3516 75058 3528
rect 75822 3516 75828 3528
rect 75052 3488 75828 3516
rect 75052 3476 75058 3488
rect 75822 3476 75828 3488
rect 75880 3476 75886 3528
rect 76190 3476 76196 3528
rect 76248 3516 76254 3528
rect 77202 3516 77208 3528
rect 76248 3488 77208 3516
rect 76248 3476 76254 3488
rect 77202 3476 77208 3488
rect 77260 3476 77266 3528
rect 83274 3476 83280 3528
rect 83332 3516 83338 3528
rect 84102 3516 84108 3528
rect 83332 3488 84108 3516
rect 83332 3476 83338 3488
rect 84102 3476 84108 3488
rect 84160 3476 84166 3528
rect 84470 3476 84476 3528
rect 84528 3516 84534 3528
rect 85482 3516 85488 3528
rect 84528 3488 85488 3516
rect 84528 3476 84534 3488
rect 85482 3476 85488 3488
rect 85540 3476 85546 3528
rect 85666 3476 85672 3528
rect 85724 3516 85730 3528
rect 86770 3516 86776 3528
rect 85724 3488 86776 3516
rect 85724 3476 85730 3488
rect 86770 3476 86776 3488
rect 86828 3476 86834 3528
rect 89162 3476 89168 3528
rect 89220 3516 89226 3528
rect 89622 3516 89628 3528
rect 89220 3488 89628 3516
rect 89220 3476 89226 3488
rect 89622 3476 89628 3488
rect 89680 3476 89686 3528
rect 90358 3476 90364 3528
rect 90416 3516 90422 3528
rect 91002 3516 91008 3528
rect 90416 3488 91008 3516
rect 90416 3476 90422 3488
rect 91002 3476 91008 3488
rect 91060 3476 91066 3528
rect 92750 3476 92756 3528
rect 92808 3516 92814 3528
rect 93762 3516 93768 3528
rect 92808 3488 93768 3516
rect 92808 3476 92814 3488
rect 93762 3476 93768 3488
rect 93820 3476 93826 3528
rect 93946 3476 93952 3528
rect 94004 3516 94010 3528
rect 95050 3516 95056 3528
rect 94004 3488 95056 3516
rect 94004 3476 94010 3488
rect 95050 3476 95056 3488
rect 95108 3476 95114 3528
rect 98638 3476 98644 3528
rect 98696 3516 98702 3528
rect 99282 3516 99288 3528
rect 98696 3488 99288 3516
rect 98696 3476 98702 3488
rect 99282 3476 99288 3488
rect 99340 3476 99346 3528
rect 99834 3476 99840 3528
rect 99892 3516 99898 3528
rect 100662 3516 100668 3528
rect 99892 3488 100668 3516
rect 99892 3476 99898 3488
rect 100662 3476 100668 3488
rect 100720 3476 100726 3528
rect 102226 3476 102232 3528
rect 102284 3516 102290 3528
rect 106826 3516 106832 3528
rect 102284 3488 106832 3516
rect 102284 3476 102290 3488
rect 106826 3476 106832 3488
rect 106884 3476 106890 3528
rect 106918 3476 106924 3528
rect 106976 3516 106982 3528
rect 107562 3516 107568 3528
rect 106976 3488 107568 3516
rect 106976 3476 106982 3488
rect 107562 3476 107568 3488
rect 107620 3476 107626 3528
rect 108298 3516 108304 3528
rect 107672 3488 108304 3516
rect 6454 3408 6460 3460
rect 6512 3448 6518 3460
rect 31018 3448 31024 3460
rect 6512 3420 31024 3448
rect 6512 3408 6518 3420
rect 31018 3408 31024 3420
rect 31076 3408 31082 3460
rect 31294 3408 31300 3460
rect 31352 3448 31358 3460
rect 39298 3448 39304 3460
rect 31352 3420 39304 3448
rect 31352 3408 31358 3420
rect 39298 3408 39304 3420
rect 39356 3408 39362 3460
rect 66714 3408 66720 3460
rect 66772 3448 66778 3460
rect 90266 3448 90272 3460
rect 66772 3420 90272 3448
rect 66772 3408 66778 3420
rect 90266 3408 90272 3420
rect 90324 3408 90330 3460
rect 91554 3408 91560 3460
rect 91612 3448 91618 3460
rect 107672 3448 107700 3488
rect 108298 3476 108304 3488
rect 108356 3476 108362 3528
rect 110506 3476 110512 3528
rect 110564 3516 110570 3528
rect 111702 3516 111708 3528
rect 110564 3488 111708 3516
rect 110564 3476 110570 3488
rect 111702 3476 111708 3488
rect 111760 3476 111766 3528
rect 137278 3516 137284 3528
rect 113146 3488 137284 3516
rect 91612 3420 107700 3448
rect 91612 3408 91618 3420
rect 108114 3408 108120 3460
rect 108172 3448 108178 3460
rect 113146 3448 113174 3488
rect 137278 3476 137284 3488
rect 137336 3476 137342 3528
rect 140038 3476 140044 3528
rect 140096 3516 140102 3528
rect 141142 3516 141148 3528
rect 140096 3488 141148 3516
rect 140096 3476 140102 3488
rect 141142 3476 141148 3488
rect 141200 3476 141206 3528
rect 143534 3476 143540 3528
rect 143592 3516 143598 3528
rect 144822 3516 144828 3528
rect 143592 3488 144828 3516
rect 143592 3476 143598 3488
rect 144822 3476 144828 3488
rect 144880 3476 144886 3528
rect 238018 3476 238024 3528
rect 238076 3516 238082 3528
rect 260650 3516 260656 3528
rect 238076 3488 260656 3516
rect 238076 3476 238082 3488
rect 260650 3476 260656 3488
rect 260708 3476 260714 3528
rect 287698 3476 287704 3528
rect 287756 3516 287762 3528
rect 290182 3516 290188 3528
rect 287756 3488 290188 3516
rect 287756 3476 287762 3488
rect 290182 3476 290188 3488
rect 290240 3476 290246 3528
rect 290458 3476 290464 3528
rect 290516 3516 290522 3528
rect 294874 3516 294880 3528
rect 290516 3488 294880 3516
rect 290516 3476 290522 3488
rect 294874 3476 294880 3488
rect 294932 3476 294938 3528
rect 299474 3476 299480 3528
rect 299532 3516 299538 3528
rect 300762 3516 300768 3528
rect 299532 3488 300768 3516
rect 299532 3476 299538 3488
rect 300762 3476 300768 3488
rect 300820 3476 300826 3528
rect 304902 3476 304908 3528
rect 304960 3516 304966 3528
rect 305546 3516 305552 3528
rect 304960 3488 305552 3516
rect 304960 3476 304966 3488
rect 305546 3476 305552 3488
rect 305604 3476 305610 3528
rect 307754 3476 307760 3528
rect 307812 3516 307818 3528
rect 309042 3516 309048 3528
rect 307812 3488 309048 3516
rect 307812 3476 307818 3488
rect 309042 3476 309048 3488
rect 309100 3476 309106 3528
rect 319714 3476 319720 3528
rect 319772 3516 319778 3528
rect 320174 3516 320180 3528
rect 319772 3488 320180 3516
rect 319772 3476 319778 3488
rect 320174 3476 320180 3488
rect 320232 3476 320238 3528
rect 324314 3476 324320 3528
rect 324372 3516 324378 3528
rect 325602 3516 325608 3528
rect 324372 3488 325608 3516
rect 324372 3476 324378 3488
rect 325602 3476 325608 3488
rect 325660 3476 325666 3528
rect 340138 3476 340144 3528
rect 340196 3516 340202 3528
rect 342162 3516 342168 3528
rect 340196 3488 342168 3516
rect 340196 3476 340202 3488
rect 342162 3476 342168 3488
rect 342220 3476 342226 3528
rect 108172 3420 113174 3448
rect 108172 3408 108178 3420
rect 114002 3408 114008 3460
rect 114060 3448 114066 3460
rect 114462 3448 114468 3460
rect 114060 3420 114468 3448
rect 114060 3408 114066 3420
rect 114462 3408 114468 3420
rect 114520 3408 114526 3460
rect 115198 3408 115204 3460
rect 115256 3448 115262 3460
rect 115842 3448 115848 3460
rect 115256 3420 115848 3448
rect 115256 3408 115262 3420
rect 115842 3408 115848 3420
rect 115900 3408 115906 3460
rect 116394 3408 116400 3460
rect 116452 3448 116458 3460
rect 117222 3448 117228 3460
rect 116452 3420 117228 3448
rect 116452 3408 116458 3420
rect 117222 3408 117228 3420
rect 117280 3408 117286 3460
rect 117590 3408 117596 3460
rect 117648 3448 117654 3460
rect 118602 3448 118608 3460
rect 117648 3420 118608 3448
rect 117648 3408 117654 3420
rect 118602 3408 118608 3420
rect 118660 3408 118666 3460
rect 118786 3408 118792 3460
rect 118844 3448 118850 3460
rect 155218 3448 155224 3460
rect 118844 3420 155224 3448
rect 118844 3408 118850 3420
rect 155218 3408 155224 3420
rect 155276 3408 155282 3460
rect 213362 3408 213368 3460
rect 213420 3448 213426 3460
rect 242894 3448 242900 3460
rect 213420 3420 242900 3448
rect 213420 3408 213426 3420
rect 242894 3408 242900 3420
rect 242952 3408 242958 3460
rect 246298 3408 246304 3460
rect 246356 3448 246362 3460
rect 247586 3448 247592 3460
rect 246356 3420 247592 3448
rect 246356 3408 246362 3420
rect 247586 3408 247592 3420
rect 247644 3408 247650 3460
rect 257062 3408 257068 3460
rect 257120 3448 257126 3460
rect 258166 3448 258172 3460
rect 257120 3420 258172 3448
rect 257120 3408 257126 3420
rect 258166 3408 258172 3420
rect 258224 3408 258230 3460
rect 260098 3408 260104 3460
rect 260156 3448 260162 3460
rect 272426 3448 272432 3460
rect 260156 3420 272432 3448
rect 260156 3408 260162 3420
rect 272426 3408 272432 3420
rect 272484 3408 272490 3460
rect 273898 3408 273904 3460
rect 273956 3448 273962 3460
rect 283098 3448 283104 3460
rect 273956 3420 283104 3448
rect 273956 3408 273962 3420
rect 283098 3408 283104 3420
rect 283156 3408 283162 3460
rect 295978 3408 295984 3460
rect 296036 3448 296042 3460
rect 301958 3448 301964 3460
rect 296036 3420 301964 3448
rect 296036 3408 296042 3420
rect 301958 3408 301964 3420
rect 302016 3408 302022 3460
rect 341518 3408 341524 3460
rect 341576 3448 341582 3460
rect 350442 3448 350448 3460
rect 341576 3420 350448 3448
rect 341576 3408 341582 3420
rect 350442 3408 350448 3420
rect 350500 3408 350506 3460
rect 262858 3272 262864 3324
rect 262916 3312 262922 3324
rect 267734 3312 267740 3324
rect 262916 3284 267740 3312
rect 262916 3272 262922 3284
rect 267734 3272 267740 3284
rect 267792 3272 267798 3324
rect 268470 3272 268476 3324
rect 268528 3312 268534 3324
rect 273622 3312 273628 3324
rect 268528 3284 273628 3312
rect 268528 3272 268534 3284
rect 273622 3272 273628 3284
rect 273680 3272 273686 3324
rect 280798 3272 280804 3324
rect 280856 3312 280862 3324
rect 284294 3312 284300 3324
rect 280856 3284 284300 3312
rect 280856 3272 280862 3284
rect 284294 3272 284300 3284
rect 284352 3272 284358 3324
rect 25314 3136 25320 3188
rect 25372 3176 25378 3188
rect 26142 3176 26148 3188
rect 25372 3148 26148 3176
rect 25372 3136 25378 3148
rect 26142 3136 26148 3148
rect 26200 3136 26206 3188
rect 349246 3136 349252 3188
rect 349304 3176 349310 3188
rect 351914 3176 351920 3188
rect 349304 3148 351920 3176
rect 349304 3136 349310 3148
rect 351914 3136 351920 3148
rect 351972 3136 351978 3188
rect 27706 3068 27712 3120
rect 27764 3108 27770 3120
rect 29638 3108 29644 3120
rect 27764 3080 29644 3108
rect 27764 3068 27770 3080
rect 29638 3068 29644 3080
rect 29696 3068 29702 3120
rect 299658 3068 299664 3120
rect 299716 3108 299722 3120
rect 302234 3108 302240 3120
rect 299716 3080 302240 3108
rect 299716 3068 299722 3080
rect 302234 3068 302240 3080
rect 302292 3068 302298 3120
rect 77386 3000 77392 3052
rect 77444 3040 77450 3052
rect 79318 3040 79324 3052
rect 77444 3012 79324 3040
rect 77444 3000 77450 3012
rect 79318 3000 79324 3012
rect 79376 3000 79382 3052
rect 289078 2932 289084 2984
rect 289136 2972 289142 2984
rect 292574 2972 292580 2984
rect 289136 2944 292580 2972
rect 289136 2932 289142 2944
rect 292574 2932 292580 2944
rect 292632 2932 292638 2984
rect 327718 2932 327724 2984
rect 327776 2972 327782 2984
rect 332686 2972 332692 2984
rect 327776 2944 332692 2972
rect 327776 2932 327782 2944
rect 332686 2932 332692 2944
rect 332744 2932 332750 2984
rect 339862 2932 339868 2984
rect 339920 2972 339926 2984
rect 342346 2972 342352 2984
rect 339920 2944 342352 2972
rect 339920 2932 339926 2944
rect 342346 2932 342352 2944
rect 342404 2932 342410 2984
rect 580994 2932 581000 2984
rect 581052 2972 581058 2984
rect 583110 2972 583116 2984
rect 581052 2944 583116 2972
rect 581052 2932 581058 2944
rect 583110 2932 583116 2944
rect 583168 2932 583174 2984
rect 15930 2864 15936 2916
rect 15988 2904 15994 2916
rect 16482 2904 16488 2916
rect 15988 2876 16488 2904
rect 15988 2864 15994 2876
rect 16482 2864 16488 2876
rect 16540 2864 16546 2916
rect 51350 2048 51356 2100
rect 51408 2088 51414 2100
rect 101398 2088 101404 2100
rect 51408 2060 101404 2088
rect 51408 2048 51414 2060
rect 101398 2048 101404 2060
rect 101456 2048 101462 2100
<< via1 >>
rect 264244 703332 264296 703384
rect 332508 703332 332560 703384
rect 70308 703264 70360 703316
rect 154120 703264 154172 703316
rect 282184 703264 282236 703316
rect 397460 703264 397512 703316
rect 90364 703196 90416 703248
rect 235172 703196 235224 703248
rect 273904 703196 273956 703248
rect 413652 703196 413704 703248
rect 119344 703128 119396 703180
rect 218980 703128 219032 703180
rect 280804 703128 280856 703180
rect 462320 703128 462372 703180
rect 102048 703060 102100 703112
rect 300124 703060 300176 703112
rect 67640 702992 67692 703044
rect 170312 702992 170364 703044
rect 287704 702992 287756 703044
rect 580172 702992 580224 703044
rect 71780 702924 71832 702976
rect 72976 702924 73028 702976
rect 84108 702924 84160 702976
rect 202788 702924 202840 702976
rect 286324 702924 286376 702976
rect 543464 702924 543516 702976
rect 61936 702856 61988 702908
rect 364984 702856 365036 702908
rect 97264 702788 97316 702840
rect 478512 702788 478564 702840
rect 24308 702720 24360 702772
rect 86224 702720 86276 702772
rect 116584 702720 116636 702772
rect 429844 702720 429896 702772
rect 77208 702652 77260 702704
rect 494796 702652 494848 702704
rect 8116 702584 8168 702636
rect 94688 702584 94740 702636
rect 105636 702584 105688 702636
rect 527180 702584 527232 702636
rect 57796 702516 57848 702568
rect 582380 702516 582432 702568
rect 66076 702448 66128 702500
rect 559656 702448 559708 702500
rect 71688 700272 71740 700324
rect 105452 700272 105504 700324
rect 277308 700272 277360 700324
rect 283840 700272 283892 700324
rect 87604 699660 87656 699712
rect 89168 699660 89220 699712
rect 3516 670692 3568 670744
rect 17224 670692 17276 670744
rect 3516 656888 3568 656940
rect 15844 656888 15896 656940
rect 3516 632068 3568 632120
rect 21364 632068 21416 632120
rect 3516 618264 3568 618316
rect 43444 618264 43496 618316
rect 2780 605888 2832 605940
rect 4804 605888 4856 605940
rect 67548 589908 67600 589960
rect 71688 589908 71740 589960
rect 124220 589908 124272 589960
rect 40040 588548 40092 588600
rect 95332 588548 95384 588600
rect 84108 587868 84160 587920
rect 101404 587868 101456 587920
rect 4804 587120 4856 587172
rect 96620 587120 96672 587172
rect 86500 586508 86552 586560
rect 140780 586508 140832 586560
rect 78588 585760 78640 585812
rect 87604 585760 87656 585812
rect 121736 585760 121788 585812
rect 582656 585760 582708 585812
rect 82728 585216 82780 585268
rect 98644 585216 98696 585268
rect 55128 585148 55180 585200
rect 77944 585148 77996 585200
rect 78588 585148 78640 585200
rect 87512 585148 87564 585200
rect 121460 585148 121512 585200
rect 121736 585148 121788 585200
rect 92112 583788 92164 583840
rect 73528 583720 73580 583772
rect 111064 583720 111116 583772
rect 122840 583720 122892 583772
rect 582840 583720 582892 583772
rect 81808 582564 81860 582616
rect 84108 582564 84160 582616
rect 62028 582428 62080 582480
rect 73804 582428 73856 582480
rect 93768 582428 93820 582480
rect 105544 582428 105596 582480
rect 52368 582360 52420 582412
rect 69940 582360 69992 582412
rect 76288 582360 76340 582412
rect 87880 582360 87932 582412
rect 90272 582360 90324 582412
rect 103520 582360 103572 582412
rect 87880 581612 87932 581664
rect 108304 581612 108356 581664
rect 69664 581068 69716 581120
rect 80244 581068 80296 581120
rect 50988 581000 51040 581052
rect 90548 581000 90600 581052
rect 57888 580252 57940 580304
rect 69664 580660 69716 580712
rect 85488 580660 85540 580712
rect 3332 579640 3384 579692
rect 57888 579640 57940 579692
rect 64788 579640 64840 579692
rect 66812 579640 66864 579692
rect 94688 580456 94740 580508
rect 94688 580252 94740 580304
rect 113456 579640 113508 579692
rect 96896 578212 96948 578264
rect 130384 578212 130436 578264
rect 102048 576920 102100 576972
rect 118700 576920 118752 576972
rect 97080 576852 97132 576904
rect 128360 576852 128412 576904
rect 97908 576716 97960 576768
rect 102048 576716 102100 576768
rect 21364 576104 21416 576156
rect 31760 576104 31812 576156
rect 31760 575492 31812 575544
rect 33048 575492 33100 575544
rect 66536 575492 66588 575544
rect 94780 574744 94832 574796
rect 120080 574744 120132 574796
rect 96252 574064 96304 574116
rect 105636 574064 105688 574116
rect 56508 571956 56560 572008
rect 66444 571956 66496 572008
rect 64696 571344 64748 571396
rect 66720 571344 66772 571396
rect 107568 570596 107620 570648
rect 582748 570596 582800 570648
rect 97908 569916 97960 569968
rect 107568 569916 107620 569968
rect 97908 569168 97960 569220
rect 133880 569168 133932 569220
rect 3424 568488 3476 568540
rect 4804 568488 4856 568540
rect 60648 567196 60700 567248
rect 66996 567196 67048 567248
rect 52276 565836 52328 565888
rect 67640 565836 67692 565888
rect 41328 564408 41380 564460
rect 66720 564408 66772 564460
rect 57796 564340 57848 564392
rect 66444 564340 66496 564392
rect 48136 563660 48188 563712
rect 57796 563660 57848 563712
rect 50896 560260 50948 560312
rect 66996 560260 67048 560312
rect 59176 558900 59228 558952
rect 66996 558900 67048 558952
rect 97264 558152 97316 558204
rect 115204 558152 115256 558204
rect 53748 557540 53800 557592
rect 66996 557540 67048 557592
rect 97356 555432 97408 555484
rect 121552 555432 121604 555484
rect 63316 554752 63368 554804
rect 66996 554752 67048 554804
rect 3516 553800 3568 553852
rect 7564 553800 7616 553852
rect 57796 553392 57848 553444
rect 66996 553392 67048 553444
rect 96988 552032 97040 552084
rect 109684 552032 109736 552084
rect 96804 551896 96856 551948
rect 96804 551692 96856 551744
rect 97908 550604 97960 550656
rect 115940 550604 115992 550656
rect 48044 549244 48096 549296
rect 66536 549244 66588 549296
rect 53472 546456 53524 546508
rect 66996 546456 67048 546508
rect 95148 546456 95200 546508
rect 96712 546456 96764 546508
rect 54944 544348 54996 544400
rect 61936 544348 61988 544400
rect 66720 544348 66772 544400
rect 97540 543736 97592 543788
rect 108396 543736 108448 543788
rect 3424 540200 3476 540252
rect 34520 540200 34572 540252
rect 67732 539792 67784 539844
rect 71780 539792 71832 539844
rect 93216 539792 93268 539844
rect 94688 539792 94740 539844
rect 70308 539656 70360 539708
rect 72332 539656 72384 539708
rect 34520 539588 34572 539640
rect 35716 539588 35768 539640
rect 61292 539588 61344 539640
rect 67824 539520 67876 539572
rect 68928 539520 68980 539572
rect 68928 538840 68980 538892
rect 82912 538840 82964 538892
rect 88248 538296 88300 538348
rect 95424 538296 95476 538348
rect 15844 538228 15896 538280
rect 93952 538228 94004 538280
rect 7564 538160 7616 538212
rect 70676 538160 70728 538212
rect 90364 538160 90416 538212
rect 136640 538160 136692 538212
rect 61844 537480 61896 537532
rect 96896 537480 96948 537532
rect 70676 536800 70728 536852
rect 71136 536800 71188 536852
rect 43444 536732 43496 536784
rect 73436 536732 73488 536784
rect 86868 536732 86920 536784
rect 119344 536732 119396 536784
rect 61292 536664 61344 536716
rect 69388 536664 69440 536716
rect 73436 535712 73488 535764
rect 76564 535712 76616 535764
rect 72792 535440 72844 535492
rect 73804 535440 73856 535492
rect 91008 535440 91060 535492
rect 92756 535440 92808 535492
rect 3424 534692 3476 534744
rect 94504 534692 94556 534744
rect 49516 533400 49568 533452
rect 84292 533400 84344 533452
rect 88340 533400 88392 533452
rect 88892 533400 88944 533452
rect 80060 533332 80112 533384
rect 80612 533332 80664 533384
rect 84016 533332 84068 533384
rect 136640 533332 136692 533384
rect 60004 531972 60056 532024
rect 98092 531972 98144 532024
rect 65984 529184 66036 529236
rect 117320 529184 117372 529236
rect 3516 527824 3568 527876
rect 128360 527824 128412 527876
rect 75184 526396 75236 526448
rect 96804 526396 96856 526448
rect 109684 521568 109736 521620
rect 111800 521568 111852 521620
rect 71044 520888 71096 520940
rect 91192 520888 91244 520940
rect 55036 518168 55088 518220
rect 98000 518168 98052 518220
rect 3516 514768 3568 514820
rect 40684 514768 40736 514820
rect 50896 511232 50948 511284
rect 580172 511232 580224 511284
rect 63316 490560 63368 490612
rect 128452 490560 128504 490612
rect 80152 487772 80204 487824
rect 129740 487772 129792 487824
rect 71136 485052 71188 485104
rect 122932 485052 122984 485104
rect 66076 482264 66128 482316
rect 118792 482264 118844 482316
rect 3424 478116 3476 478168
rect 15844 478116 15896 478168
rect 67732 478116 67784 478168
rect 98736 478116 98788 478168
rect 85488 475124 85540 475176
rect 93216 475124 93268 475176
rect 77208 473288 77260 473340
rect 77944 473288 77996 473340
rect 73804 472608 73856 472660
rect 116124 472608 116176 472660
rect 82820 467100 82872 467152
rect 109040 467100 109092 467152
rect 65984 466420 66036 466472
rect 70492 466420 70544 466472
rect 86316 464312 86368 464364
rect 95240 464312 95292 464364
rect 85580 462952 85632 463004
rect 120172 462952 120224 463004
rect 3516 462340 3568 462392
rect 14464 462340 14516 462392
rect 67732 460164 67784 460216
rect 96712 460164 96764 460216
rect 64788 458804 64840 458856
rect 92572 458804 92624 458856
rect 86868 457512 86920 457564
rect 104348 457512 104400 457564
rect 64604 457444 64656 457496
rect 86960 457444 87012 457496
rect 64696 454656 64748 454708
rect 106924 454656 106976 454708
rect 60648 453296 60700 453348
rect 123116 453296 123168 453348
rect 79324 451868 79376 451920
rect 90364 451868 90416 451920
rect 68928 449896 68980 449948
rect 80060 449896 80112 449948
rect 78680 449216 78732 449268
rect 101496 449216 101548 449268
rect 53748 449148 53800 449200
rect 85672 449148 85724 449200
rect 101404 449148 101456 449200
rect 117504 449148 117556 449200
rect 3148 448536 3200 448588
rect 36544 448536 36596 448588
rect 78036 447856 78088 447908
rect 91100 447856 91152 447908
rect 88340 447788 88392 447840
rect 113272 447788 113324 447840
rect 91008 446428 91060 446480
rect 118884 446428 118936 446480
rect 52368 446360 52420 446412
rect 95976 446360 96028 446412
rect 95884 444388 95936 444440
rect 96528 444388 96580 444440
rect 116032 444388 116084 444440
rect 81440 443708 81492 443760
rect 96528 443708 96580 443760
rect 48136 443640 48188 443692
rect 88432 443640 88484 443692
rect 100024 443640 100076 443692
rect 115296 443640 115348 443692
rect 93860 442960 93912 443012
rect 95148 442960 95200 443012
rect 124312 442960 124364 443012
rect 40684 442892 40736 442944
rect 103520 442892 103572 442944
rect 115204 442892 115256 442944
rect 120264 442892 120316 442944
rect 106280 442280 106332 442332
rect 106924 442280 106976 442332
rect 77300 442212 77352 442264
rect 113364 442212 113416 442264
rect 106280 441600 106332 441652
rect 131120 441600 131172 441652
rect 54944 440920 54996 440972
rect 78404 440920 78456 440972
rect 67640 440852 67692 440904
rect 114560 440852 114612 440904
rect 102600 438948 102652 439000
rect 102784 438948 102836 439000
rect 127072 438948 127124 439000
rect 108120 438880 108172 438932
rect 108396 438880 108448 438932
rect 137284 438880 137336 438932
rect 50896 438132 50948 438184
rect 74724 438132 74776 438184
rect 122196 438132 122248 438184
rect 583116 438132 583168 438184
rect 108304 437520 108356 437572
rect 125600 437520 125652 437572
rect 95976 437452 96028 437504
rect 122196 437452 122248 437504
rect 71136 437384 71188 437436
rect 75184 437384 75236 437436
rect 57704 436160 57756 436212
rect 73988 436160 74040 436212
rect 77944 436160 77996 436212
rect 82912 436160 82964 436212
rect 33784 436092 33836 436144
rect 71136 436092 71188 436144
rect 76840 436092 76892 436144
rect 79324 436092 79376 436144
rect 98736 436092 98788 436144
rect 99932 436092 99984 436144
rect 101496 436092 101548 436144
rect 103704 436092 103756 436144
rect 123024 436160 123076 436212
rect 111064 436092 111116 436144
rect 140872 436092 140924 436144
rect 68468 435344 68520 435396
rect 71780 435344 71832 435396
rect 72700 435344 72752 435396
rect 72608 434800 72660 434852
rect 132500 434800 132552 434852
rect 4804 434732 4856 434784
rect 111800 434732 111852 434784
rect 112444 434732 112496 434784
rect 117412 434732 117464 434784
rect 67364 433984 67416 434036
rect 74540 433984 74592 434036
rect 105912 433984 105964 434036
rect 118976 433984 119028 434036
rect 68376 433712 68428 433764
rect 71228 433712 71280 433764
rect 68652 433644 68704 433696
rect 69204 433644 69256 433696
rect 110880 433644 110932 433696
rect 61752 433304 61804 433356
rect 63408 433304 63460 433356
rect 66260 433304 66312 433356
rect 112720 433236 112772 433288
rect 112720 432012 112772 432064
rect 117596 432012 117648 432064
rect 59084 431944 59136 431996
rect 66444 431944 66496 431996
rect 115572 431944 115624 431996
rect 133972 431944 134024 431996
rect 60556 430584 60608 430636
rect 66720 430584 66772 430636
rect 115848 430584 115900 430636
rect 135904 430584 135956 430636
rect 115756 430516 115808 430568
rect 136640 430516 136692 430568
rect 142804 430516 142856 430568
rect 52368 429224 52420 429276
rect 66720 429224 66772 429276
rect 115848 429088 115900 429140
rect 118792 429088 118844 429140
rect 124864 429088 124916 429140
rect 60648 427796 60700 427848
rect 66720 427796 66772 427848
rect 53748 426436 53800 426488
rect 66720 426436 66772 426488
rect 118792 426368 118844 426420
rect 122840 426368 122892 426420
rect 50896 425688 50948 425740
rect 65984 425688 66036 425740
rect 66536 425688 66588 425740
rect 115848 425076 115900 425128
rect 118792 425076 118844 425128
rect 115848 424328 115900 424380
rect 144920 424328 144972 424380
rect 44088 423648 44140 423700
rect 66720 423648 66772 423700
rect 115756 423648 115808 423700
rect 126980 423648 127032 423700
rect 2780 423580 2832 423632
rect 4804 423580 4856 423632
rect 115848 423580 115900 423632
rect 122932 423580 122984 423632
rect 124128 423580 124180 423632
rect 60740 423444 60792 423496
rect 61844 423444 61896 423496
rect 66720 423444 66772 423496
rect 49608 422900 49660 422952
rect 60740 422900 60792 422952
rect 124128 422900 124180 422952
rect 148324 422900 148376 422952
rect 50988 422220 51040 422272
rect 66996 422220 67048 422272
rect 41236 421540 41288 421592
rect 50988 421540 51040 421592
rect 114560 421540 114612 421592
rect 146944 421540 146996 421592
rect 61844 419500 61896 419552
rect 66904 419500 66956 419552
rect 115756 419500 115808 419552
rect 129832 419500 129884 419552
rect 32956 418140 33008 418192
rect 66904 418208 66956 418260
rect 64788 418140 64840 418192
rect 66628 418140 66680 418192
rect 57796 417392 57848 417444
rect 66628 417392 66680 417444
rect 64144 416848 64196 416900
rect 66996 416848 67048 416900
rect 115848 416780 115900 416832
rect 143540 416780 143592 416832
rect 116216 416712 116268 416764
rect 118976 416712 119028 416764
rect 115848 415692 115900 415744
rect 116216 415692 116268 415744
rect 53564 415420 53616 415472
rect 60004 415420 60056 415472
rect 115848 414808 115900 414860
rect 117320 414808 117372 414860
rect 121644 414808 121696 414860
rect 60004 414740 60056 414792
rect 66904 414740 66956 414792
rect 56416 413992 56468 414044
rect 66720 413992 66772 414044
rect 115112 413992 115164 414044
rect 115296 413992 115348 414044
rect 147680 413992 147732 414044
rect 46848 413244 46900 413296
rect 59268 413244 59320 413296
rect 66904 413244 66956 413296
rect 115848 412632 115900 412684
rect 121552 412632 121604 412684
rect 122932 412632 122984 412684
rect 115204 411884 115256 411936
rect 116124 411884 116176 411936
rect 142160 411884 142212 411936
rect 59268 411272 59320 411324
rect 64604 411272 64656 411324
rect 66720 411272 66772 411324
rect 52276 411204 52328 411256
rect 66904 411204 66956 411256
rect 115848 411204 115900 411256
rect 123208 411204 123260 411256
rect 124128 411204 124180 411256
rect 124128 410524 124180 410576
rect 136640 410524 136692 410576
rect 50988 409912 51040 409964
rect 52276 409912 52328 409964
rect 2872 409844 2924 409896
rect 51724 409844 51776 409896
rect 53840 409776 53892 409828
rect 55036 409776 55088 409828
rect 66260 409776 66312 409828
rect 115848 409776 115900 409828
rect 120264 409776 120316 409828
rect 39948 409096 40000 409148
rect 53840 409096 53892 409148
rect 120264 409096 120316 409148
rect 139400 409096 139452 409148
rect 39856 408416 39908 408468
rect 66904 408416 66956 408468
rect 35808 407736 35860 407788
rect 39856 407736 39908 407788
rect 115020 407464 115072 407516
rect 121552 407464 121604 407516
rect 56508 407056 56560 407108
rect 57796 407056 57848 407108
rect 112720 407056 112772 407108
rect 117596 407056 117648 407108
rect 57796 405696 57848 405748
rect 66444 405696 66496 405748
rect 115848 405628 115900 405680
rect 140780 405628 140832 405680
rect 141424 405628 141476 405680
rect 117320 405560 117372 405612
rect 117504 405560 117556 405612
rect 115848 404540 115900 404592
rect 117320 404540 117372 404592
rect 63224 404336 63276 404388
rect 66904 404336 66956 404388
rect 141424 404336 141476 404388
rect 143632 404336 143684 404388
rect 115848 402976 115900 403028
rect 126336 402976 126388 403028
rect 115848 401956 115900 402008
rect 118976 401956 119028 402008
rect 120172 401956 120224 402008
rect 115848 401548 115900 401600
rect 128452 401548 128504 401600
rect 128452 400868 128504 400920
rect 146300 400868 146352 400920
rect 58900 400256 58952 400308
rect 66812 400256 66864 400308
rect 57612 400188 57664 400240
rect 66904 400188 66956 400240
rect 115388 399168 115440 399220
rect 117504 399168 117556 399220
rect 55036 398828 55088 398880
rect 66536 398828 66588 398880
rect 3516 397536 3568 397588
rect 21364 397536 21416 397588
rect 11704 397468 11756 397520
rect 67364 397536 67416 397588
rect 67732 397536 67784 397588
rect 115572 397468 115624 397520
rect 124220 397468 124272 397520
rect 66720 397400 66772 397452
rect 67732 397400 67784 397452
rect 128452 397400 128504 397452
rect 132592 397400 132644 397452
rect 42708 396788 42760 396840
rect 59176 396788 59228 396840
rect 66628 396788 66680 396840
rect 35716 396720 35768 396772
rect 117504 396720 117556 396772
rect 149060 396720 149112 396772
rect 67088 396652 67140 396704
rect 115848 396040 115900 396092
rect 128452 396040 128504 396092
rect 49516 395972 49568 396024
rect 66812 395972 66864 396024
rect 48228 395224 48280 395276
rect 49516 395224 49568 395276
rect 115848 394680 115900 394732
rect 190460 394680 190512 394732
rect 43996 393932 44048 393984
rect 49516 393932 49568 393984
rect 49516 393320 49568 393372
rect 66812 393320 66864 393372
rect 115848 393252 115900 393304
rect 128360 393252 128412 393304
rect 53656 392572 53708 392624
rect 66352 392572 66404 392624
rect 56508 391960 56560 392012
rect 66812 391960 66864 392012
rect 128360 391960 128412 392012
rect 134064 391960 134116 392012
rect 41328 391280 41380 391332
rect 3424 391212 3476 391264
rect 118884 391212 118936 391264
rect 138020 391212 138072 391264
rect 115020 391144 115072 391196
rect 120172 391144 120224 391196
rect 87696 390940 87748 390992
rect 108672 390940 108724 390992
rect 118884 390940 118936 390992
rect 93676 390872 93728 390924
rect 67640 390124 67692 390176
rect 68790 390124 68842 390176
rect 102048 389784 102100 389836
rect 113272 389784 113324 389836
rect 118700 389784 118752 389836
rect 128360 389784 128412 389836
rect 94596 389444 94648 389496
rect 62028 389240 62080 389292
rect 36544 389172 36596 389224
rect 100760 389376 100812 389428
rect 94596 389308 94648 389360
rect 98276 389308 98328 389360
rect 101680 389172 101732 389224
rect 118700 389172 118752 389224
rect 48044 389104 48096 389156
rect 83004 389104 83056 389156
rect 97264 389104 97316 389156
rect 110144 389036 110196 389088
rect 124772 389036 124824 389088
rect 46756 388696 46808 388748
rect 48044 388696 48096 388748
rect 102232 388492 102284 388544
rect 106372 388492 106424 388544
rect 84108 388424 84160 388476
rect 104164 388424 104216 388476
rect 105544 388424 105596 388476
rect 114744 388424 114796 388476
rect 71688 387812 71740 387864
rect 73252 387812 73304 387864
rect 79968 387812 80020 387864
rect 80704 387812 80756 387864
rect 84936 387812 84988 387864
rect 86224 387812 86276 387864
rect 90364 387812 90416 387864
rect 91376 387812 91428 387864
rect 93124 387812 93176 387864
rect 96988 387812 97040 387864
rect 100576 387812 100628 387864
rect 102508 387812 102560 387864
rect 57888 387744 57940 387796
rect 96620 387744 96672 387796
rect 120724 387744 120776 387796
rect 121460 387744 121512 387796
rect 101864 387132 101916 387184
rect 107660 387132 107712 387184
rect 52276 387064 52328 387116
rect 73988 387064 74040 387116
rect 86868 387064 86920 387116
rect 120724 387064 120776 387116
rect 84200 386996 84252 387048
rect 85028 386996 85080 387048
rect 111800 386996 111852 387048
rect 112260 386996 112312 387048
rect 96620 386384 96672 386436
rect 97356 386384 97408 386436
rect 65892 386316 65944 386368
rect 72424 386316 72476 386368
rect 75184 386316 75236 386368
rect 82268 386316 82320 386368
rect 80796 386248 80848 386300
rect 81256 386248 81308 386300
rect 115940 386316 115992 386368
rect 100392 386248 100444 386300
rect 129740 386248 129792 386300
rect 130292 386248 130344 386300
rect 54852 385636 54904 385688
rect 66812 385636 66864 385688
rect 130292 385024 130344 385076
rect 134156 385024 134208 385076
rect 55128 384956 55180 385008
rect 92480 384956 92532 385008
rect 133144 384956 133196 385008
rect 133880 384956 133932 385008
rect 91192 384344 91244 384396
rect 109132 384344 109184 384396
rect 105176 384276 105228 384328
rect 133144 384276 133196 384328
rect 88432 383596 88484 383648
rect 120080 383596 120132 383648
rect 101772 382916 101824 382968
rect 112720 382916 112772 382968
rect 120080 382236 120132 382288
rect 122840 382236 122892 382288
rect 45468 381488 45520 381540
rect 71780 381488 71832 381540
rect 84200 381488 84252 381540
rect 117320 381488 117372 381540
rect 21364 380808 21416 380860
rect 116216 380808 116268 380860
rect 94504 380128 94556 380180
rect 128544 380128 128596 380180
rect 115940 380060 115992 380112
rect 116216 380060 116268 380112
rect 79968 379516 80020 379568
rect 81440 379516 81492 379568
rect 88248 379448 88300 379500
rect 91376 379448 91428 379500
rect 43996 378768 44048 378820
rect 80060 378768 80112 378820
rect 100484 378768 100536 378820
rect 129740 378768 129792 378820
rect 97816 378224 97868 378276
rect 102324 378224 102376 378276
rect 92296 378088 92348 378140
rect 93124 378088 93176 378140
rect 87696 377476 87748 377528
rect 118700 377476 118752 377528
rect 33048 377408 33100 377460
rect 92296 377408 92348 377460
rect 41328 374620 41380 374672
rect 76012 374620 76064 374672
rect 86776 374620 86828 374672
rect 95332 374620 95384 374672
rect 101956 373260 102008 373312
rect 113180 373260 113232 373312
rect 3424 371220 3476 371272
rect 106188 371152 106240 371204
rect 118976 371152 119028 371204
rect 50804 369112 50856 369164
rect 75920 369112 75972 369164
rect 80704 369112 80756 369164
rect 102140 369112 102192 369164
rect 85580 367752 85632 367804
rect 106924 367752 106976 367804
rect 74540 366324 74592 366376
rect 108304 366324 108356 366376
rect 269764 364352 269816 364404
rect 580172 364352 580224 364404
rect 86224 363604 86276 363656
rect 112444 363604 112496 363656
rect 77300 360816 77352 360868
rect 110604 360816 110656 360868
rect 3332 358708 3384 358760
rect 11704 358708 11756 358760
rect 3424 355308 3476 355360
rect 33784 355308 33836 355360
rect 574744 351908 574796 351960
rect 580172 351908 580224 351960
rect 3332 345040 3384 345092
rect 18604 345040 18656 345092
rect 123484 343612 123536 343664
rect 124128 343612 124180 343664
rect 260840 343612 260892 343664
rect 97724 342252 97776 342304
rect 267832 342252 267884 342304
rect 124864 340892 124916 340944
rect 125508 340892 125560 340944
rect 263600 340892 263652 340944
rect 83556 339464 83608 339516
rect 259828 339464 259880 339516
rect 23388 338104 23440 338156
rect 222200 338104 222252 338156
rect 153844 336812 153896 336864
rect 233884 336812 233936 336864
rect 93124 336744 93176 336796
rect 93676 336744 93728 336796
rect 255964 336744 256016 336796
rect 87604 335792 87656 335844
rect 88248 335792 88300 335844
rect 88248 335316 88300 335368
rect 256700 335316 256752 335368
rect 100024 333956 100076 334008
rect 100576 333956 100628 334008
rect 246304 333956 246356 334008
rect 148416 332664 148468 332716
rect 266452 332664 266504 332716
rect 99288 332596 99340 332648
rect 244924 332596 244976 332648
rect 115204 331304 115256 331356
rect 115388 331304 115440 331356
rect 244188 331304 244240 331356
rect 57612 331236 57664 331288
rect 57888 331236 57940 331288
rect 266360 331236 266412 331288
rect 93676 331168 93728 331220
rect 94044 331168 94096 331220
rect 166356 329808 166408 329860
rect 227812 329808 227864 329860
rect 104808 328720 104860 328772
rect 110512 328720 110564 328772
rect 192484 328516 192536 328568
rect 250444 328516 250496 328568
rect 151084 328448 151136 328500
rect 212540 328448 212592 328500
rect 81440 327700 81492 327752
rect 91284 327700 91336 327752
rect 105728 327700 105780 327752
rect 129832 327700 129884 327752
rect 251824 327700 251876 327752
rect 162124 327088 162176 327140
rect 212632 327088 212684 327140
rect 85396 327020 85448 327072
rect 88340 327020 88392 327072
rect 103520 327020 103572 327072
rect 110696 327020 110748 327072
rect 114008 325728 114060 325780
rect 249064 325728 249116 325780
rect 61384 325660 61436 325712
rect 110696 325660 110748 325712
rect 270592 325660 270644 325712
rect 67732 325592 67784 325644
rect 108488 324980 108540 325032
rect 125600 324980 125652 325032
rect 259644 324980 259696 325032
rect 67732 324912 67784 324964
rect 252744 324912 252796 324964
rect 113824 323552 113876 323604
rect 121644 323552 121696 323604
rect 262220 323552 262272 323604
rect 53564 322872 53616 322924
rect 59360 322872 59412 322924
rect 256792 322940 256844 322992
rect 89444 322872 89496 322924
rect 93860 322872 93912 322924
rect 78496 322736 78548 322788
rect 84384 322736 84436 322788
rect 180064 321648 180116 321700
rect 245016 321648 245068 321700
rect 137376 321580 137428 321632
rect 254216 321580 254268 321632
rect 127072 321512 127124 321564
rect 264244 321512 264296 321564
rect 263784 321036 263836 321088
rect 264244 321036 264296 321088
rect 92204 320900 92256 320952
rect 123024 320900 123076 320952
rect 125324 320900 125376 320952
rect 64604 320832 64656 320884
rect 75184 320832 75236 320884
rect 89812 320832 89864 320884
rect 127072 320832 127124 320884
rect 53104 320152 53156 320204
rect 63500 320152 63552 320204
rect 64144 320152 64196 320204
rect 125324 320152 125376 320204
rect 261024 320152 261076 320204
rect 98368 319472 98420 319524
rect 106280 319472 106332 319524
rect 63500 319404 63552 319456
rect 251916 319404 251968 319456
rect 68468 318588 68520 318640
rect 69112 318588 69164 318640
rect 95884 317432 95936 317484
rect 116584 317432 116636 317484
rect 74540 316888 74592 316940
rect 81532 316888 81584 316940
rect 99288 316752 99340 316804
rect 117412 316752 117464 316804
rect 131028 316752 131080 316804
rect 82912 316684 82964 316736
rect 124312 316684 124364 316736
rect 125416 316684 125468 316736
rect 185584 316072 185636 316124
rect 267740 316072 267792 316124
rect 131028 316004 131080 316056
rect 250536 316004 250588 316056
rect 273352 315460 273404 315512
rect 273904 315460 273956 315512
rect 97908 315256 97960 315308
rect 273352 315256 273404 315308
rect 96620 314644 96672 314696
rect 97908 314644 97960 314696
rect 151268 314644 151320 314696
rect 247684 314644 247736 314696
rect 186320 313352 186372 313404
rect 265072 313352 265124 313404
rect 105636 313284 105688 313336
rect 106188 313284 106240 313336
rect 252836 313284 252888 313336
rect 3424 313216 3476 313268
rect 7564 313216 7616 313268
rect 67272 312536 67324 312588
rect 258172 312536 258224 312588
rect 187148 311856 187200 311908
rect 263876 311856 263928 311908
rect 278044 311856 278096 311908
rect 580172 311856 580224 311908
rect 109684 311108 109736 311160
rect 134064 311108 134116 311160
rect 259552 311108 259604 311160
rect 189816 310496 189868 310548
rect 261116 310496 261168 310548
rect 104164 310428 104216 310480
rect 108396 310428 108448 310480
rect 97724 309748 97776 309800
rect 117412 309748 117464 309800
rect 148324 309204 148376 309256
rect 238024 309204 238076 309256
rect 122748 309136 122800 309188
rect 220176 309136 220228 309188
rect 67364 309068 67416 309120
rect 186320 309068 186372 309120
rect 188436 307844 188488 307896
rect 254124 307844 254176 307896
rect 22008 307776 22060 307828
rect 202420 307776 202472 307828
rect 202512 307776 202564 307828
rect 262404 307776 262456 307828
rect 182916 306416 182968 306468
rect 210424 306416 210476 306468
rect 175924 306348 175976 306400
rect 241060 306348 241112 306400
rect 65892 305600 65944 305652
rect 151268 305600 151320 305652
rect 232504 305600 232556 305652
rect 269212 305600 269264 305652
rect 192576 305056 192628 305108
rect 255504 305056 255556 305108
rect 3240 304988 3292 305040
rect 32404 304988 32456 305040
rect 152464 304988 152516 305040
rect 216772 304988 216824 305040
rect 113916 304308 113968 304360
rect 123484 304308 123536 304360
rect 85580 304240 85632 304292
rect 95884 304240 95936 304292
rect 96436 304240 96488 304292
rect 108488 304240 108540 304292
rect 114100 304240 114152 304292
rect 125508 304240 125560 304292
rect 135996 304240 136048 304292
rect 246304 304240 246356 304292
rect 251272 304240 251324 304292
rect 250444 304036 250496 304088
rect 253940 304036 253992 304088
rect 142804 303764 142856 303816
rect 216128 303764 216180 303816
rect 170404 303696 170456 303748
rect 214196 303696 214248 303748
rect 215300 303696 215352 303748
rect 228916 303696 228968 303748
rect 213920 303628 213972 303680
rect 229560 303628 229612 303680
rect 233884 303628 233936 303680
rect 237840 303628 237892 303680
rect 240048 303628 240100 303680
rect 250628 303628 250680 303680
rect 149060 303560 149112 303612
rect 240692 303560 240744 303612
rect 247408 303560 247460 303612
rect 141608 302880 141660 302932
rect 149060 302880 149112 302932
rect 245016 302880 245068 302932
rect 252744 302880 252796 302932
rect 256884 302880 256936 302932
rect 274732 302880 274784 302932
rect 250536 302404 250588 302456
rect 256884 302404 256936 302456
rect 77300 302200 77352 302252
rect 78496 302200 78548 302252
rect 131856 302200 131908 302252
rect 191380 302200 191432 302252
rect 211068 302200 211120 302252
rect 255964 302132 256016 302184
rect 259736 302132 259788 302184
rect 249064 301860 249116 301912
rect 255688 301860 255740 301912
rect 79968 301452 80020 301504
rect 103612 301452 103664 301504
rect 189816 301452 189868 301504
rect 193312 301112 193364 301164
rect 195428 300976 195480 301028
rect 178684 300840 178736 300892
rect 190368 300772 190420 300824
rect 211988 300976 212040 301028
rect 208860 300908 208912 300960
rect 219440 300908 219492 300960
rect 244280 300908 244332 300960
rect 270500 300840 270552 300892
rect 179328 300160 179380 300212
rect 190460 300160 190512 300212
rect 126428 300092 126480 300144
rect 190552 300092 190604 300144
rect 252928 300092 252980 300144
rect 252836 299820 252888 299872
rect 253112 299820 253164 299872
rect 56508 299480 56560 299532
rect 159456 299480 159508 299532
rect 255412 299480 255464 299532
rect 287060 299480 287112 299532
rect 146944 299412 146996 299464
rect 191012 299412 191064 299464
rect 580908 299412 580960 299464
rect 583576 299412 583628 299464
rect 255320 298120 255372 298172
rect 288440 298120 288492 298172
rect 160100 298052 160152 298104
rect 161296 298052 161348 298104
rect 191104 298052 191156 298104
rect 255320 297984 255372 298036
rect 255504 297984 255556 298036
rect 255596 296760 255648 296812
rect 260932 296760 260984 296812
rect 82820 296692 82872 296744
rect 84016 296692 84068 296744
rect 184204 296692 184256 296744
rect 255504 296692 255556 296744
rect 282920 296692 282972 296744
rect 124128 295944 124180 295996
rect 192484 295944 192536 295996
rect 256056 295468 256108 295520
rect 258356 295468 258408 295520
rect 69664 295332 69716 295384
rect 156604 295332 156656 295384
rect 190460 295332 190512 295384
rect 255504 295332 255556 295384
rect 284392 295332 284444 295384
rect 120172 295264 120224 295316
rect 190552 295264 190604 295316
rect 180248 294584 180300 294636
rect 193312 294584 193364 294636
rect 117228 294040 117280 294092
rect 120172 294040 120224 294092
rect 255596 294040 255648 294092
rect 267924 294040 267976 294092
rect 69572 293972 69624 294024
rect 70216 293972 70268 294024
rect 126520 293972 126572 294024
rect 255504 293972 255556 294024
rect 273260 293972 273312 294024
rect 59176 293292 59228 293344
rect 87604 293292 87656 293344
rect 84568 293224 84620 293276
rect 93032 293224 93084 293276
rect 124128 293224 124180 293276
rect 169024 293224 169076 293276
rect 192576 293224 192628 293276
rect 255504 293224 255556 293276
rect 270592 293224 270644 293276
rect 71688 292612 71740 292664
rect 71964 292612 72016 292664
rect 3424 292544 3476 292596
rect 18696 292544 18748 292596
rect 36544 292544 36596 292596
rect 58992 292544 59044 292596
rect 59176 292544 59228 292596
rect 122104 292544 122156 292596
rect 193128 292544 193180 292596
rect 255596 292544 255648 292596
rect 280160 292544 280212 292596
rect 101404 292476 101456 292528
rect 193220 292476 193272 292528
rect 101496 291796 101548 291848
rect 114008 291796 114060 291848
rect 255688 291796 255740 291848
rect 269120 291796 269172 291848
rect 91468 291184 91520 291236
rect 97264 291184 97316 291236
rect 255504 291184 255556 291236
rect 262312 291184 262364 291236
rect 255504 290980 255556 291032
rect 259644 290980 259696 291032
rect 83004 289892 83056 289944
rect 84108 289892 84160 289944
rect 103520 289892 103572 289944
rect 94504 289824 94556 289876
rect 193220 289824 193272 289876
rect 255504 289756 255556 289808
rect 262220 289756 262272 289808
rect 82728 289076 82780 289128
rect 94504 289076 94556 289128
rect 45376 288464 45428 288516
rect 79324 288464 79376 288516
rect 79600 288464 79652 288516
rect 95608 288464 95660 288516
rect 96436 288464 96488 288516
rect 112536 288464 112588 288516
rect 142988 288464 143040 288516
rect 186228 288464 186280 288516
rect 191012 288464 191064 288516
rect 78588 288396 78640 288448
rect 168288 288396 168340 288448
rect 18604 288328 18656 288380
rect 71044 288328 71096 288380
rect 180064 288328 180116 288380
rect 255504 288328 255556 288380
rect 262404 288328 262456 288380
rect 127624 287648 127676 287700
rect 137376 287648 137428 287700
rect 159456 287648 159508 287700
rect 166908 287648 166960 287700
rect 95148 287104 95200 287156
rect 127624 287104 127676 287156
rect 60464 287036 60516 287088
rect 79416 287036 79468 287088
rect 96528 287036 96580 287088
rect 162860 287036 162912 287088
rect 166908 287036 166960 287088
rect 191748 287036 191800 287088
rect 255504 287036 255556 287088
rect 258356 287036 258408 287088
rect 259460 287036 259512 287088
rect 92388 286968 92440 287020
rect 93124 286968 93176 287020
rect 94688 286968 94740 287020
rect 255320 286968 255372 287020
rect 255596 286968 255648 287020
rect 261024 286968 261076 287020
rect 255504 286900 255556 286952
rect 176108 286356 176160 286408
rect 188712 286356 188764 286408
rect 71780 286288 71832 286340
rect 77024 286288 77076 286340
rect 188436 286288 188488 286340
rect 255412 286288 255464 286340
rect 267740 286288 267792 286340
rect 64512 285676 64564 285728
rect 80796 285676 80848 285728
rect 69480 284928 69532 284980
rect 69664 284928 69716 284980
rect 82912 284928 82964 284980
rect 83556 284928 83608 284980
rect 63132 284384 63184 284436
rect 72424 284384 72476 284436
rect 86868 284384 86920 284436
rect 98460 284384 98512 284436
rect 158720 284384 158772 284436
rect 191564 284384 191616 284436
rect 255504 284384 255556 284436
rect 266360 284384 266412 284436
rect 68560 284316 68612 284368
rect 164976 284316 165028 284368
rect 255412 284316 255464 284368
rect 269304 284316 269356 284368
rect 89950 283704 90002 283756
rect 91008 283704 91060 283756
rect 53472 283568 53524 283620
rect 57704 283568 57756 283620
rect 66812 283568 66864 283620
rect 68836 283568 68888 283620
rect 169024 283568 169076 283620
rect 66168 283024 66220 283076
rect 69664 282956 69716 283008
rect 81440 282956 81492 283008
rect 89628 282956 89680 283008
rect 63316 282820 63368 282872
rect 178040 282888 178092 282940
rect 179236 282888 179288 282940
rect 191012 282888 191064 282940
rect 255412 282888 255464 282940
rect 270684 282888 270736 282940
rect 192392 282820 192444 282872
rect 255504 282820 255556 282872
rect 262496 282820 262548 282872
rect 69020 282684 69072 282736
rect 255412 282684 255464 282736
rect 258264 282684 258316 282736
rect 98000 282208 98052 282260
rect 98736 282208 98788 282260
rect 100760 281528 100812 281580
rect 149704 281528 149756 281580
rect 107016 281460 107068 281512
rect 158720 281460 158772 281512
rect 162860 281460 162912 281512
rect 164148 281460 164200 281512
rect 255412 281460 255464 281512
rect 265072 281460 265124 281512
rect 100760 281392 100812 281444
rect 135904 281392 135956 281444
rect 164148 280780 164200 280832
rect 191748 280780 191800 280832
rect 10324 280168 10376 280220
rect 67272 280168 67324 280220
rect 68836 280168 68888 280220
rect 255412 280168 255464 280220
rect 262220 280168 262272 280220
rect 126980 280100 127032 280152
rect 127440 280100 127492 280152
rect 185584 280100 185636 280152
rect 100760 280032 100812 280084
rect 142896 280032 142948 280084
rect 7564 279420 7616 279472
rect 34336 279420 34388 279472
rect 65892 279420 65944 279472
rect 66536 279420 66588 279472
rect 102232 279420 102284 279472
rect 127440 279420 127492 279472
rect 255320 278740 255372 278792
rect 266544 278740 266596 278792
rect 47952 278672 48004 278724
rect 48136 278672 48188 278724
rect 99380 278672 99432 278724
rect 102048 278672 102100 278724
rect 122104 278672 122156 278724
rect 255504 278672 255556 278724
rect 263876 278672 263928 278724
rect 152648 278060 152700 278112
rect 188528 278060 188580 278112
rect 47952 277992 48004 278044
rect 66812 277992 66864 278044
rect 98460 277992 98512 278044
rect 177856 277992 177908 278044
rect 255412 277448 255464 277500
rect 259736 277448 259788 277500
rect 188620 277380 188672 277432
rect 191656 277380 191708 277432
rect 55128 277312 55180 277364
rect 66904 277312 66956 277364
rect 177948 277312 178000 277364
rect 187148 277312 187200 277364
rect 255412 277108 255464 277160
rect 259552 277108 259604 277160
rect 100760 276632 100812 276684
rect 118792 276632 118844 276684
rect 169208 276632 169260 276684
rect 190460 276632 190512 276684
rect 61936 276156 61988 276208
rect 66812 276156 66864 276208
rect 255504 276020 255556 276072
rect 273444 276020 273496 276072
rect 64696 275952 64748 276004
rect 66628 275952 66680 276004
rect 255412 275952 255464 276004
rect 267832 275952 267884 276004
rect 100852 275340 100904 275392
rect 148416 275340 148468 275392
rect 54944 275272 54996 275324
rect 61936 275272 61988 275324
rect 100116 275272 100168 275324
rect 181628 275272 181680 275324
rect 255412 274660 255464 274712
rect 281632 274660 281684 274712
rect 100760 274592 100812 274644
rect 146944 274592 146996 274644
rect 255504 274592 255556 274644
rect 269212 274592 269264 274644
rect 274640 274592 274692 274644
rect 255320 274524 255372 274576
rect 258080 274524 258132 274576
rect 134616 273912 134668 273964
rect 156696 273912 156748 273964
rect 180064 273232 180116 273284
rect 191656 273232 191708 273284
rect 100760 273164 100812 273216
rect 105728 273164 105780 273216
rect 255412 273164 255464 273216
rect 263692 273164 263744 273216
rect 106188 272552 106240 272604
rect 142988 272552 143040 272604
rect 146944 272552 146996 272604
rect 180156 272552 180208 272604
rect 46664 272484 46716 272536
rect 52368 272484 52420 272536
rect 66812 272484 66864 272536
rect 124128 272484 124180 272536
rect 175924 272484 175976 272536
rect 101128 272008 101180 272060
rect 101864 272008 101916 272060
rect 104900 272008 104952 272060
rect 106188 272008 106240 272060
rect 187148 271940 187200 271992
rect 191656 271940 191708 271992
rect 181536 271872 181588 271924
rect 191564 271872 191616 271924
rect 565084 271872 565136 271924
rect 580172 271872 580224 271924
rect 99288 271532 99340 271584
rect 105544 271532 105596 271584
rect 148416 271192 148468 271244
rect 188344 271192 188396 271244
rect 53748 271124 53800 271176
rect 66260 271124 66312 271176
rect 141516 271124 141568 271176
rect 187056 271124 187108 271176
rect 255964 271124 256016 271176
rect 266452 271124 266504 271176
rect 100300 270444 100352 270496
rect 106188 270444 106240 270496
rect 56324 269764 56376 269816
rect 66260 269764 66312 269816
rect 126520 269764 126572 269816
rect 159456 269764 159508 269816
rect 255504 269152 255556 269204
rect 261024 269152 261076 269204
rect 166264 269084 166316 269136
rect 191656 269084 191708 269136
rect 255412 269084 255464 269136
rect 268016 269084 268068 269136
rect 115940 268608 115992 268660
rect 116676 268608 116728 268660
rect 101220 268404 101272 268456
rect 113824 268404 113876 268456
rect 44088 268336 44140 268388
rect 53564 268336 53616 268388
rect 100760 268336 100812 268388
rect 115940 268336 115992 268388
rect 145564 268336 145616 268388
rect 166356 268336 166408 268388
rect 255412 267792 255464 267844
rect 267832 267792 267884 267844
rect 53564 267724 53616 267776
rect 66812 267724 66864 267776
rect 164884 267724 164936 267776
rect 191656 267724 191708 267776
rect 255320 267724 255372 267776
rect 273536 267724 273588 267776
rect 3516 267656 3568 267708
rect 36544 267656 36596 267708
rect 100760 267656 100812 267708
rect 122932 267656 122984 267708
rect 255504 267656 255556 267708
rect 277308 267656 277360 267708
rect 142896 266976 142948 267028
rect 173256 266976 173308 267028
rect 173164 266432 173216 266484
rect 191012 266432 191064 266484
rect 63316 266364 63368 266416
rect 66812 266364 66864 266416
rect 122932 266364 122984 266416
rect 131764 266364 131816 266416
rect 157984 266364 158036 266416
rect 191288 266364 191340 266416
rect 255412 266364 255464 266416
rect 265164 266364 265216 266416
rect 277308 266364 277360 266416
rect 277492 266364 277544 266416
rect 100852 266296 100904 266348
rect 142160 266296 142212 266348
rect 143448 266296 143500 266348
rect 254032 266296 254084 266348
rect 263784 266296 263836 266348
rect 143448 265684 143500 265736
rect 152556 265684 152608 265736
rect 41236 265616 41288 265668
rect 50528 265616 50580 265668
rect 105544 265616 105596 265668
rect 115296 265616 115348 265668
rect 140044 265616 140096 265668
rect 182916 265616 182968 265668
rect 61844 265140 61896 265192
rect 65708 265140 65760 265192
rect 255320 265004 255372 265056
rect 263692 265004 263744 265056
rect 167644 264936 167696 264988
rect 191564 264936 191616 264988
rect 100760 264868 100812 264920
rect 139400 264868 139452 264920
rect 144276 264868 144328 264920
rect 98276 264188 98328 264240
rect 115296 264188 115348 264240
rect 147128 264188 147180 264240
rect 176108 264188 176160 264240
rect 255320 263644 255372 263696
rect 271972 263644 272024 263696
rect 273352 263644 273404 263696
rect 3424 263576 3476 263628
rect 99288 263576 99340 263628
rect 101220 263576 101272 263628
rect 255504 263576 255556 263628
rect 278872 263576 278924 263628
rect 282184 263576 282236 263628
rect 53104 263508 53156 263560
rect 66904 263508 66956 263560
rect 101680 263508 101732 263560
rect 103428 263508 103480 263560
rect 117964 263508 118016 263560
rect 255412 263032 255464 263084
rect 258356 263032 258408 263084
rect 7564 262828 7616 262880
rect 32956 262828 33008 262880
rect 65892 262828 65944 262880
rect 66536 262828 66588 262880
rect 141424 262828 141476 262880
rect 153844 262828 153896 262880
rect 121368 262624 121420 262676
rect 121552 262624 121604 262676
rect 177304 262284 177356 262336
rect 191656 262284 191708 262336
rect 100760 262216 100812 262268
rect 121368 262216 121420 262268
rect 126336 262216 126388 262268
rect 191196 262216 191248 262268
rect 255412 262216 255464 262268
rect 265072 262216 265124 262268
rect 255504 262148 255556 262200
rect 285680 262148 285732 262200
rect 255320 262080 255372 262132
rect 263600 262080 263652 262132
rect 103428 261536 103480 261588
rect 109040 261536 109092 261588
rect 56416 261468 56468 261520
rect 66260 261468 66312 261520
rect 108212 261468 108264 261520
rect 143632 261468 143684 261520
rect 180248 261468 180300 261520
rect 171784 260856 171836 260908
rect 191656 260856 191708 260908
rect 100760 260788 100812 260840
rect 108212 260788 108264 260840
rect 255412 260788 255464 260840
rect 287704 260788 287756 260840
rect 55128 260176 55180 260228
rect 59360 260176 59412 260228
rect 66812 260176 66864 260228
rect 46756 260108 46808 260160
rect 55864 260108 55916 260160
rect 57520 260108 57572 260160
rect 66260 260108 66312 260160
rect 144184 260108 144236 260160
rect 178684 260108 178736 260160
rect 289728 260108 289780 260160
rect 582380 260108 582432 260160
rect 101220 259836 101272 259888
rect 102784 259836 102836 259888
rect 174544 259428 174596 259480
rect 191288 259428 191340 259480
rect 255412 259428 255464 259480
rect 288532 259428 288584 259480
rect 289728 259428 289780 259480
rect 59268 259360 59320 259412
rect 66444 259360 66496 259412
rect 100760 259360 100812 259412
rect 126336 259360 126388 259412
rect 50620 258680 50672 258732
rect 57612 258680 57664 258732
rect 66260 258680 66312 258732
rect 278688 258680 278740 258732
rect 582472 258680 582524 258732
rect 100760 258204 100812 258256
rect 105636 258204 105688 258256
rect 175924 258068 175976 258120
rect 190460 258068 190512 258120
rect 255504 258068 255556 258120
rect 277584 258068 277636 258120
rect 278688 258068 278740 258120
rect 190552 258000 190604 258052
rect 193404 258000 193456 258052
rect 268108 258000 268160 258052
rect 582840 258000 582892 258052
rect 100760 257388 100812 257440
rect 101128 257388 101180 257440
rect 105544 257388 105596 257440
rect 113824 257388 113876 257440
rect 138020 257388 138072 257440
rect 152556 257388 152608 257440
rect 178684 257388 178736 257440
rect 50988 257320 51040 257372
rect 59084 257320 59136 257372
rect 66812 257320 66864 257372
rect 137468 257320 137520 257372
rect 173256 257320 173308 257372
rect 255320 257320 255372 257372
rect 268108 257320 268160 257372
rect 185584 256708 185636 256760
rect 191656 256708 191708 256760
rect 255504 256708 255556 256760
rect 270776 256708 270828 256760
rect 101036 256640 101088 256692
rect 141608 256640 141660 256692
rect 255412 256640 255464 256692
rect 266636 256640 266688 256692
rect 39948 255960 40000 256012
rect 51080 255960 51132 256012
rect 137376 255960 137428 256012
rect 186964 255960 187016 256012
rect 273352 255960 273404 256012
rect 580264 255960 580316 256012
rect 51080 255280 51132 255332
rect 52000 255280 52052 255332
rect 66812 255280 66864 255332
rect 108948 255280 109000 255332
rect 111892 255280 111944 255332
rect 181444 255280 181496 255332
rect 190644 255280 190696 255332
rect 255504 255280 255556 255332
rect 272064 255280 272116 255332
rect 3148 255212 3200 255264
rect 10324 255212 10376 255264
rect 266728 255212 266780 255264
rect 583024 255212 583076 255264
rect 109040 255144 109092 255196
rect 113916 255144 113968 255196
rect 273628 255144 273680 255196
rect 583392 255144 583444 255196
rect 255504 254600 255556 254652
rect 266728 254600 266780 254652
rect 57796 254532 57848 254584
rect 59176 254532 59228 254584
rect 66812 254532 66864 254584
rect 100760 254532 100812 254584
rect 106648 254532 106700 254584
rect 121368 254532 121420 254584
rect 184388 254532 184440 254584
rect 255412 254532 255464 254584
rect 273628 254532 273680 254584
rect 100852 253920 100904 253972
rect 109040 253920 109092 253972
rect 110420 253920 110472 253972
rect 111064 253920 111116 253972
rect 151268 253920 151320 253972
rect 169116 253920 169168 253972
rect 191656 253920 191708 253972
rect 63224 253852 63276 253904
rect 66536 253852 66588 253904
rect 100760 253852 100812 253904
rect 140780 253852 140832 253904
rect 141056 253852 141108 253904
rect 255596 253852 255648 253904
rect 255964 253852 256016 253904
rect 583208 253852 583260 253904
rect 100852 253172 100904 253224
rect 126428 253172 126480 253224
rect 255412 253172 255464 253224
rect 269396 253172 269448 253224
rect 269764 253172 269816 253224
rect 186964 252560 187016 252612
rect 191656 252560 191708 252612
rect 103336 251880 103388 251932
rect 111800 251880 111852 251932
rect 256240 251880 256292 251932
rect 256976 251880 257028 251932
rect 278044 251880 278096 251932
rect 106188 251812 106240 251864
rect 115204 251812 115256 251864
rect 120080 251812 120132 251864
rect 263876 251812 263928 251864
rect 583576 251812 583628 251864
rect 64788 251336 64840 251388
rect 65984 251336 66036 251388
rect 66260 251336 66312 251388
rect 185676 251268 185728 251320
rect 190828 251268 190880 251320
rect 255412 251268 255464 251320
rect 263876 251268 263928 251320
rect 163504 251200 163556 251252
rect 191656 251200 191708 251252
rect 58900 251132 58952 251184
rect 61844 251132 61896 251184
rect 106280 251132 106332 251184
rect 109684 251132 109736 251184
rect 57888 251064 57940 251116
rect 66904 251064 66956 251116
rect 61016 250724 61068 250776
rect 61384 250724 61436 250776
rect 66812 250724 66864 250776
rect 262496 250520 262548 250572
rect 273352 250520 273404 250572
rect 101956 250452 102008 250504
rect 114560 250452 114612 250504
rect 153844 250452 153896 250504
rect 162124 250452 162176 250504
rect 164976 250452 165028 250504
rect 192576 250452 192628 250504
rect 265256 250452 265308 250504
rect 582380 250452 582432 250504
rect 255504 249840 255556 249892
rect 262496 249840 262548 249892
rect 57888 249772 57940 249824
rect 100760 249772 100812 249824
rect 106280 249772 106332 249824
rect 115388 249772 115440 249824
rect 159548 249772 159600 249824
rect 170496 249772 170548 249824
rect 191656 249772 191708 249824
rect 255412 249772 255464 249824
rect 265256 249772 265308 249824
rect 59268 249704 59320 249756
rect 100760 249636 100812 249688
rect 101128 249636 101180 249688
rect 101680 249024 101732 249076
rect 103336 249024 103388 249076
rect 140780 249024 140832 249076
rect 160836 249024 160888 249076
rect 169208 249024 169260 249076
rect 55036 248412 55088 248464
rect 57796 248412 57848 248464
rect 66812 248412 66864 248464
rect 106924 248412 106976 248464
rect 192484 248480 192536 248532
rect 255412 248480 255464 248532
rect 278044 248480 278096 248532
rect 188528 248412 188580 248464
rect 191656 248412 191708 248464
rect 255320 248412 255372 248464
rect 266636 248412 266688 248464
rect 582380 248412 582432 248464
rect 42708 248344 42760 248396
rect 61936 248344 61988 248396
rect 66904 248344 66956 248396
rect 99196 248344 99248 248396
rect 108948 248344 109000 248396
rect 108948 247732 109000 247784
rect 166356 247732 166408 247784
rect 105544 247664 105596 247716
rect 117320 247664 117372 247716
rect 177396 247664 177448 247716
rect 255412 247120 255464 247172
rect 272156 247120 272208 247172
rect 184296 247052 184348 247104
rect 191656 247052 191708 247104
rect 256424 247052 256476 247104
rect 256884 247052 256936 247104
rect 582380 247052 582432 247104
rect 101128 246984 101180 247036
rect 111064 246984 111116 247036
rect 56508 246304 56560 246356
rect 66812 246304 66864 246356
rect 101036 246304 101088 246356
rect 104808 246304 104860 246356
rect 128452 246304 128504 246356
rect 140780 246304 140832 246356
rect 193680 246304 193732 246356
rect 255412 245692 255464 245744
rect 287152 245692 287204 245744
rect 187240 245624 187292 245676
rect 190644 245624 190696 245676
rect 48228 244944 48280 244996
rect 57888 244944 57940 244996
rect 53656 244876 53708 244928
rect 67548 244876 67600 244928
rect 102232 244876 102284 244928
rect 113824 244876 113876 244928
rect 255504 244400 255556 244452
rect 258172 244400 258224 244452
rect 108396 244264 108448 244316
rect 165528 244264 165580 244316
rect 255412 244264 255464 244316
rect 285772 244264 285824 244316
rect 69020 243516 69072 243568
rect 169208 243516 169260 243568
rect 49516 242904 49568 242956
rect 55036 242904 55088 242956
rect 66260 242904 66312 242956
rect 67824 242904 67876 242956
rect 68468 242904 68520 242956
rect 108304 242904 108356 242956
rect 161480 242904 161532 242956
rect 169300 242224 169352 242276
rect 54852 242156 54904 242208
rect 62120 242156 62172 242208
rect 153936 242156 153988 242208
rect 96896 241748 96948 241800
rect 99564 241748 99616 241800
rect 101036 241680 101088 241732
rect 104164 241680 104216 241732
rect 107660 241680 107712 241732
rect 70952 241612 71004 241664
rect 127716 241612 127768 241664
rect 66168 241476 66220 241528
rect 69940 241476 69992 241528
rect 95332 241476 95384 241528
rect 96206 241476 96258 241528
rect 52184 241408 52236 241460
rect 76564 241408 76616 241460
rect 76886 241408 76938 241460
rect 81302 241408 81354 241460
rect 112444 241408 112496 241460
rect 154028 241544 154080 241596
rect 193588 241612 193640 241664
rect 193772 241612 193824 241664
rect 195244 241612 195296 241664
rect 195612 241612 195664 241664
rect 249064 241612 249116 241664
rect 256976 241612 257028 241664
rect 196624 241544 196676 241596
rect 255688 241476 255740 241528
rect 256148 241476 256200 241528
rect 582564 241476 582616 241528
rect 181628 241408 181680 241460
rect 252836 241408 252888 241460
rect 256056 241408 256108 241460
rect 565084 241408 565136 241460
rect 95884 241340 95936 241392
rect 100024 241340 100076 241392
rect 165528 241340 165580 241392
rect 199108 241340 199160 241392
rect 3516 241204 3568 241256
rect 7564 241204 7616 241256
rect 64512 240728 64564 240780
rect 77944 240728 77996 240780
rect 116676 240728 116728 240780
rect 155408 240728 155460 240780
rect 224132 240728 224184 240780
rect 256700 240728 256752 240780
rect 86224 240048 86276 240100
rect 87052 240048 87104 240100
rect 98276 240048 98328 240100
rect 197544 240048 197596 240100
rect 198004 240048 198056 240100
rect 242164 240048 242216 240100
rect 242900 240048 242952 240100
rect 243544 240048 243596 240100
rect 244556 240048 244608 240100
rect 251088 240048 251140 240100
rect 254124 240048 254176 240100
rect 254768 240048 254820 240100
rect 256700 240048 256752 240100
rect 45468 239980 45520 240032
rect 71780 239980 71832 240032
rect 72516 239980 72568 240032
rect 77392 239980 77444 240032
rect 83004 239980 83056 240032
rect 75920 239912 75972 239964
rect 77484 239912 77536 239964
rect 88524 239436 88576 239488
rect 98000 239436 98052 239488
rect 234804 239436 234856 239488
rect 237472 239436 237524 239488
rect 74264 239368 74316 239420
rect 167736 239368 167788 239420
rect 202420 239368 202472 239420
rect 41328 238688 41380 238740
rect 69664 238688 69716 238740
rect 74908 238824 74960 238876
rect 226984 238756 227036 238808
rect 231584 238756 231636 238808
rect 244924 238756 244976 238808
rect 253020 238756 253072 238808
rect 80336 238688 80388 238740
rect 108396 238688 108448 238740
rect 188436 238688 188488 238740
rect 221464 238688 221516 238740
rect 81532 238620 81584 238672
rect 106924 238620 106976 238672
rect 193036 238144 193088 238196
rect 198832 238144 198884 238196
rect 63132 238076 63184 238128
rect 72424 238076 72476 238128
rect 125508 238076 125560 238128
rect 188620 238076 188672 238128
rect 69848 238008 69900 238060
rect 79324 238008 79376 238060
rect 107568 238008 107620 238060
rect 187148 238008 187200 238060
rect 204904 238008 204956 238060
rect 253940 238008 253992 238060
rect 50804 237396 50856 237448
rect 52368 237396 52420 237448
rect 222108 237396 222160 237448
rect 227812 237396 227864 237448
rect 48044 237328 48096 237380
rect 75920 237328 75972 237380
rect 77208 237328 77260 237380
rect 184388 237328 184440 237380
rect 208860 237328 208912 237380
rect 55864 237260 55916 237312
rect 80060 237260 80112 237312
rect 98000 236716 98052 236768
rect 106188 236716 106240 236768
rect 121460 236716 121512 236768
rect 76840 236648 76892 236700
rect 95240 236648 95292 236700
rect 111708 236648 111760 236700
rect 181536 236648 181588 236700
rect 193220 236648 193272 236700
rect 206284 236648 206336 236700
rect 211068 236648 211120 236700
rect 256148 236648 256200 236700
rect 103428 236240 103480 236292
rect 103704 236240 103756 236292
rect 80060 235968 80112 236020
rect 80704 235968 80756 236020
rect 97816 235968 97868 236020
rect 99472 235968 99524 236020
rect 108948 235968 109000 236020
rect 109132 235968 109184 236020
rect 208400 235968 208452 236020
rect 208860 235968 208912 236020
rect 81440 235900 81492 235952
rect 105544 235900 105596 235952
rect 170588 235900 170640 235952
rect 179420 235900 179472 235952
rect 192576 235900 192628 235952
rect 200120 235900 200172 235952
rect 200764 235900 200816 235952
rect 83004 235832 83056 235884
rect 83924 235832 83976 235884
rect 102140 235832 102192 235884
rect 43996 235220 44048 235272
rect 56508 235220 56560 235272
rect 77576 235220 77628 235272
rect 186228 235220 186280 235272
rect 195152 235220 195204 235272
rect 200764 235220 200816 235272
rect 255964 235220 256016 235272
rect 105636 234608 105688 234660
rect 105820 234608 105872 234660
rect 115940 234608 115992 234660
rect 195244 234608 195296 234660
rect 224224 234608 224276 234660
rect 73160 234540 73212 234592
rect 108304 234540 108356 234592
rect 176016 234540 176068 234592
rect 267832 234540 267884 234592
rect 83924 234404 83976 234456
rect 84108 234404 84160 234456
rect 61660 233860 61712 233912
rect 75184 233860 75236 233912
rect 97908 233860 97960 233912
rect 98184 233860 98236 233912
rect 220728 233860 220780 233912
rect 229928 233860 229980 233912
rect 278044 233248 278096 233300
rect 580172 233248 580224 233300
rect 65892 233180 65944 233232
rect 67640 233180 67692 233232
rect 82912 233180 82964 233232
rect 118700 233180 118752 233232
rect 119344 233180 119396 233232
rect 124220 233180 124272 233232
rect 177396 233180 177448 233232
rect 177948 233180 178000 233232
rect 216956 233180 217008 233232
rect 58992 233112 59044 233164
rect 86224 233112 86276 233164
rect 217324 232568 217376 232620
rect 225052 232568 225104 232620
rect 234620 232568 234672 232620
rect 256976 232568 257028 232620
rect 91100 232500 91152 232552
rect 119344 232500 119396 232552
rect 206928 232500 206980 232552
rect 236460 232500 236512 232552
rect 240784 232500 240836 232552
rect 255320 232500 255372 232552
rect 76012 231752 76064 231804
rect 110696 231752 110748 231804
rect 180248 231752 180300 231804
rect 260840 231752 260892 231804
rect 261208 231752 261260 231804
rect 272064 231752 272116 231804
rect 272340 231752 272392 231804
rect 582748 231752 582800 231804
rect 154028 231684 154080 231736
rect 205640 231684 205692 231736
rect 77208 231072 77260 231124
rect 108396 231072 108448 231124
rect 110696 231072 110748 231124
rect 153200 231072 153252 231124
rect 208492 231072 208544 231124
rect 218612 231072 218664 231124
rect 255964 231072 256016 231124
rect 272340 231072 272392 231124
rect 205640 230936 205692 230988
rect 206376 230936 206428 230988
rect 191196 230392 191248 230444
rect 212080 230392 212132 230444
rect 221004 230392 221056 230444
rect 276204 230392 276256 230444
rect 60464 229780 60516 229832
rect 76748 229780 76800 229832
rect 48044 229712 48096 229764
rect 69480 229712 69532 229764
rect 72516 229712 72568 229764
rect 86868 229712 86920 229764
rect 224132 229712 224184 229764
rect 224224 229712 224276 229764
rect 238760 229712 238812 229764
rect 245016 229712 245068 229764
rect 256884 229712 256936 229764
rect 272156 229712 272208 229764
rect 580264 229712 580316 229764
rect 102784 229032 102836 229084
rect 273536 229032 273588 229084
rect 61844 228964 61896 229016
rect 160100 228964 160152 229016
rect 160836 228964 160888 229016
rect 202788 228352 202840 228404
rect 239680 228352 239732 228404
rect 258724 228352 258776 228404
rect 269396 228352 269448 228404
rect 128360 227672 128412 227724
rect 265164 227672 265216 227724
rect 270776 227672 270828 227724
rect 582656 227672 582708 227724
rect 159548 227604 159600 227656
rect 160008 227604 160060 227656
rect 249064 227604 249116 227656
rect 95148 226992 95200 227044
rect 122656 226992 122708 227044
rect 128360 226992 128412 227044
rect 256148 226992 256200 227044
rect 270776 226992 270828 227044
rect 59084 226244 59136 226296
rect 160928 226244 160980 226296
rect 173256 226244 173308 226296
rect 263876 226244 263928 226296
rect 95148 225564 95200 225616
rect 104900 225564 104952 225616
rect 113088 225564 113140 225616
rect 238852 225564 238904 225616
rect 173256 224952 173308 225004
rect 173808 224952 173860 225004
rect 174636 224884 174688 224936
rect 240784 224884 240836 224936
rect 252468 224884 252520 224936
rect 258264 224884 258316 224936
rect 264888 224408 264940 224460
rect 267924 224408 267976 224460
rect 138664 224272 138716 224324
rect 227812 224272 227864 224324
rect 63040 224204 63092 224256
rect 174728 224204 174780 224256
rect 256884 224204 256936 224256
rect 166356 223524 166408 223576
rect 266360 223524 266412 223576
rect 112536 222844 112588 222896
rect 117320 222844 117372 222896
rect 216036 222844 216088 222896
rect 254032 222844 254084 222896
rect 187056 221552 187108 221604
rect 224224 221552 224276 221604
rect 202144 221484 202196 221536
rect 252744 221484 252796 221536
rect 47952 221416 48004 221468
rect 202236 221416 202288 221468
rect 244280 221416 244332 221468
rect 254584 221416 254636 221468
rect 67364 220736 67416 220788
rect 273444 220736 273496 220788
rect 169208 220668 169260 220720
rect 169668 220668 169720 220720
rect 243544 220668 243596 220720
rect 82728 220056 82780 220108
rect 112444 220056 112496 220108
rect 224224 219376 224276 219428
rect 265256 219376 265308 219428
rect 84016 218696 84068 218748
rect 113272 218696 113324 218748
rect 149796 218696 149848 218748
rect 230388 218696 230440 218748
rect 113272 218016 113324 218068
rect 186320 218016 186372 218068
rect 229744 217948 229796 218000
rect 230388 217948 230440 218000
rect 251824 217948 251876 218000
rect 161388 217268 161440 217320
rect 266636 217268 266688 217320
rect 49608 216588 49660 216640
rect 161388 216588 161440 216640
rect 161572 216588 161624 216640
rect 198096 215976 198148 216028
rect 251180 215976 251232 216028
rect 160744 215908 160796 215960
rect 220820 215908 220872 215960
rect 258172 215908 258224 215960
rect 89720 215228 89772 215280
rect 117412 215228 117464 215280
rect 145656 215228 145708 215280
rect 251088 215228 251140 215280
rect 253940 215228 253992 215280
rect 117412 214752 117464 214804
rect 120172 214752 120224 214804
rect 174728 214548 174780 214600
rect 178684 214548 178736 214600
rect 251824 214548 251876 214600
rect 266544 214548 266596 214600
rect 98644 213868 98696 213920
rect 104164 213868 104216 213920
rect 262220 213868 262272 213920
rect 250444 213188 250496 213240
rect 274732 213188 274784 213240
rect 97264 211760 97316 211812
rect 114560 211760 114612 211812
rect 202236 211760 202288 211812
rect 249708 211760 249760 211812
rect 114560 211148 114612 211200
rect 262404 211148 262456 211200
rect 73068 211080 73120 211132
rect 249800 211080 249852 211132
rect 250996 211080 251048 211132
rect 186320 211012 186372 211064
rect 263600 211080 263652 211132
rect 264060 211080 264112 211132
rect 151268 209720 151320 209772
rect 247040 209720 247092 209772
rect 247776 209720 247828 209772
rect 191840 209652 191892 209704
rect 255964 209652 256016 209704
rect 33048 209040 33100 209092
rect 184296 209040 184348 209092
rect 44088 207612 44140 207664
rect 185676 207612 185728 207664
rect 246212 207612 246264 207664
rect 251824 207612 251876 207664
rect 255964 207612 256016 207664
rect 276204 207612 276256 207664
rect 94688 207000 94740 207052
rect 245752 207000 245804 207052
rect 246212 207000 246264 207052
rect 135076 206932 135128 206984
rect 270684 206932 270736 206984
rect 93124 206252 93176 206304
rect 103704 206252 103756 206304
rect 134156 206252 134208 206304
rect 135076 206252 135128 206304
rect 193128 206252 193180 206304
rect 226524 206252 226576 206304
rect 88248 204960 88300 205012
rect 104900 204960 104952 205012
rect 106096 204960 106148 205012
rect 96620 204892 96672 204944
rect 125600 204892 125652 204944
rect 133144 204892 133196 204944
rect 242900 204892 242952 204944
rect 281632 204892 281684 204944
rect 106096 204280 106148 204332
rect 258080 204280 258132 204332
rect 155408 204212 155460 204264
rect 259644 204212 259696 204264
rect 46848 203532 46900 203584
rect 67824 203532 67876 203584
rect 214564 203532 214616 203584
rect 253940 203532 253992 203584
rect 152556 202784 152608 202836
rect 155316 202784 155368 202836
rect 180156 202784 180208 202836
rect 180708 202784 180760 202836
rect 244924 202784 244976 202836
rect 3332 202172 3384 202224
rect 98092 202172 98144 202224
rect 108948 202172 109000 202224
rect 118700 202172 118752 202224
rect 138664 202172 138716 202224
rect 148416 202172 148468 202224
rect 37096 202104 37148 202156
rect 188528 202104 188580 202156
rect 253204 202104 253256 202156
rect 270684 202104 270736 202156
rect 126336 201628 126388 201680
rect 134616 201628 134668 201680
rect 171876 201424 171928 201476
rect 172336 201424 172388 201476
rect 277492 201424 277544 201476
rect 133236 201356 133288 201408
rect 231860 201356 231912 201408
rect 233148 201356 233200 201408
rect 75276 200744 75328 200796
rect 107660 200744 107712 200796
rect 112628 200744 112680 200796
rect 132592 200744 132644 200796
rect 149704 200064 149756 200116
rect 252652 200064 252704 200116
rect 170956 199996 171008 200048
rect 269304 199996 269356 200048
rect 45376 199384 45428 199436
rect 76656 199384 76708 199436
rect 86224 199384 86276 199436
rect 103612 199384 103664 199436
rect 106188 199384 106240 199436
rect 122840 199384 122892 199436
rect 147036 198704 147088 198756
rect 153844 198704 153896 198756
rect 38568 197956 38620 198008
rect 224960 197956 225012 198008
rect 256056 197956 256108 198008
rect 276020 197956 276072 198008
rect 217416 196596 217468 196648
rect 242164 196596 242216 196648
rect 249064 196596 249116 196648
rect 284392 196596 284444 196648
rect 193312 195304 193364 195356
rect 224960 195304 225012 195356
rect 79968 195236 80020 195288
rect 110420 195236 110472 195288
rect 222936 195236 222988 195288
rect 271972 195236 272024 195288
rect 246304 193808 246356 193860
rect 281540 193808 281592 193860
rect 84108 192516 84160 192568
rect 107016 192516 107068 192568
rect 2688 192448 2740 192500
rect 152648 192448 152700 192500
rect 166356 192448 166408 192500
rect 217324 192448 217376 192500
rect 240784 192448 240836 192500
rect 580172 192448 580224 192500
rect 178684 191768 178736 191820
rect 278044 191768 278096 191820
rect 187608 189728 187660 189780
rect 252928 189728 252980 189780
rect 3516 188980 3568 189032
rect 18604 188980 18656 189032
rect 195888 188300 195940 188352
rect 226984 188300 227036 188352
rect 254584 188300 254636 188352
rect 270592 188300 270644 188352
rect 27528 186940 27580 186992
rect 151176 186940 151228 186992
rect 242164 186940 242216 186992
rect 260932 186940 260984 186992
rect 6828 185580 6880 185632
rect 147128 185580 147180 185632
rect 198004 185580 198056 185632
rect 226432 185580 226484 185632
rect 232596 184152 232648 184204
rect 252652 184152 252704 184204
rect 10968 182792 11020 182844
rect 188344 182792 188396 182844
rect 192484 182792 192536 182844
rect 220176 182792 220228 182844
rect 93124 180820 93176 180872
rect 93768 180820 93820 180872
rect 218704 180820 218756 180872
rect 82084 180072 82136 180124
rect 109132 180072 109184 180124
rect 195244 180072 195296 180124
rect 226616 180072 226668 180124
rect 135904 179392 135956 179444
rect 218796 179392 218848 179444
rect 252468 178644 252520 178696
rect 580172 178644 580224 178696
rect 57612 178100 57664 178152
rect 156696 178100 156748 178152
rect 90364 178032 90416 178084
rect 91008 178032 91060 178084
rect 217324 178032 217376 178084
rect 251824 178032 251876 178084
rect 252468 178032 252520 178084
rect 82820 177284 82872 177336
rect 110512 177284 110564 177336
rect 214012 177284 214064 177336
rect 252468 177284 252520 177336
rect 262312 177284 262364 177336
rect 216128 176672 216180 176724
rect 251180 176672 251232 176724
rect 252468 176672 252520 176724
rect 195244 175312 195296 175364
rect 195888 175312 195940 175364
rect 295984 175312 296036 175364
rect 78864 175244 78916 175296
rect 207112 175244 207164 175296
rect 202880 174496 202932 174548
rect 226708 174496 226760 174548
rect 82912 173884 82964 173936
rect 211804 173884 211856 173936
rect 75920 173408 75972 173460
rect 76748 173408 76800 173460
rect 76748 173136 76800 173188
rect 202880 173136 202932 173188
rect 91744 172524 91796 172576
rect 220820 172524 220872 172576
rect 195980 172320 196032 172372
rect 196808 172320 196860 172372
rect 244924 171776 244976 171828
rect 246120 171776 246172 171828
rect 177856 171164 177908 171216
rect 188344 171164 188396 171216
rect 81440 171096 81492 171148
rect 196808 171096 196860 171148
rect 246396 171096 246448 171148
rect 249432 171096 249484 171148
rect 86224 170416 86276 170468
rect 177856 170416 177908 170468
rect 196716 170416 196768 170468
rect 273260 170416 273312 170468
rect 77944 170348 77996 170400
rect 204904 170348 204956 170400
rect 205640 170348 205692 170400
rect 217416 170348 217468 170400
rect 77392 169736 77444 169788
rect 77944 169736 77996 169788
rect 123668 169668 123720 169720
rect 224868 169668 224920 169720
rect 93860 168988 93912 169040
rect 122932 168988 122984 169040
rect 123668 168988 123720 169040
rect 182916 168988 182968 169040
rect 264980 168988 265032 169040
rect 224316 168376 224368 168428
rect 224868 168376 224920 168428
rect 193036 167696 193088 167748
rect 200120 167696 200172 167748
rect 53472 167628 53524 167680
rect 210424 167628 210476 167680
rect 221464 167016 221516 167068
rect 222108 167016 222160 167068
rect 285680 167016 285732 167068
rect 195060 166336 195112 166388
rect 222108 166336 222160 166388
rect 217416 166268 217468 166320
rect 259828 166268 259880 166320
rect 197360 166064 197412 166116
rect 198096 166064 198148 166116
rect 86316 165656 86368 165708
rect 197360 165656 197412 165708
rect 75276 165588 75328 165640
rect 194600 165588 194652 165640
rect 195060 165588 195112 165640
rect 91008 164908 91060 164960
rect 117320 164908 117372 164960
rect 220820 164908 220872 164960
rect 46664 164840 46716 164892
rect 192484 164840 192536 164892
rect 198740 164840 198792 164892
rect 259460 164840 259512 164892
rect 204168 163480 204220 163532
rect 237472 163480 237524 163532
rect 306380 163480 306432 163532
rect 131764 162936 131816 162988
rect 236092 162936 236144 162988
rect 3516 162868 3568 162920
rect 8944 162868 8996 162920
rect 73068 162868 73120 162920
rect 198740 162868 198792 162920
rect 97448 162800 97500 162852
rect 97908 162800 97960 162852
rect 213920 162800 213972 162852
rect 214564 162800 214616 162852
rect 245660 162800 245712 162852
rect 246396 162800 246448 162852
rect 97448 162120 97500 162172
rect 245660 162120 245712 162172
rect 180800 161440 180852 161492
rect 181996 161440 182048 161492
rect 213276 161440 213328 161492
rect 213920 161440 213972 161492
rect 582656 161440 582708 161492
rect 34336 160692 34388 160744
rect 60740 160692 60792 160744
rect 105544 160148 105596 160200
rect 230572 160148 230624 160200
rect 60740 160080 60792 160132
rect 61752 160080 61804 160132
rect 189816 160080 189868 160132
rect 188344 159400 188396 159452
rect 211160 159400 211212 159452
rect 87144 159332 87196 159384
rect 180800 159332 180852 159384
rect 208584 159332 208636 159384
rect 274640 159332 274692 159384
rect 83464 158720 83516 158772
rect 196072 158720 196124 158772
rect 190368 157972 190420 158024
rect 249708 157972 249760 158024
rect 580356 157972 580408 158024
rect 75184 157428 75236 157480
rect 189908 157428 189960 157480
rect 90456 157360 90508 157412
rect 208584 157360 208636 157412
rect 163596 156408 163648 156460
rect 164148 156408 164200 156460
rect 56324 156000 56376 156052
rect 160836 156000 160888 156052
rect 164148 156000 164200 156052
rect 220084 156000 220136 156052
rect 222292 156000 222344 156052
rect 260104 156000 260156 156052
rect 98736 155932 98788 155984
rect 99288 155932 99340 155984
rect 225144 155932 225196 155984
rect 211252 155864 211304 155916
rect 211804 155864 211856 155916
rect 288440 155864 288492 155916
rect 289728 155864 289780 155916
rect 177396 155184 177448 155236
rect 205088 155184 205140 155236
rect 289728 155184 289780 155236
rect 317420 155184 317472 155236
rect 60372 154572 60424 154624
rect 178776 154572 178828 154624
rect 251272 154504 251324 154556
rect 251824 154504 251876 154556
rect 39856 153824 39908 153876
rect 158076 153824 158128 153876
rect 175832 153280 175884 153332
rect 227904 153280 227956 153332
rect 155316 153212 155368 153264
rect 251272 153212 251324 153264
rect 130476 152600 130528 152652
rect 131028 152600 131080 152652
rect 86868 152532 86920 152584
rect 102140 152532 102192 152584
rect 88340 152464 88392 152516
rect 154212 152464 154264 152516
rect 209044 152464 209096 152516
rect 220728 152464 220780 152516
rect 302240 152464 302292 152516
rect 180248 151852 180300 151904
rect 208400 151852 208452 151904
rect 130476 151784 130528 151836
rect 223672 151784 223724 151836
rect 208400 151036 208452 151088
rect 225052 151036 225104 151088
rect 64696 150492 64748 150544
rect 118056 150492 118108 150544
rect 206376 150492 206428 150544
rect 305000 150492 305052 150544
rect 80520 150424 80572 150476
rect 208400 150424 208452 150476
rect 67732 149676 67784 149728
rect 159916 149676 159968 149728
rect 185492 149676 185544 149728
rect 196808 149676 196860 149728
rect 209780 149676 209832 149728
rect 210240 149132 210292 149184
rect 210424 149132 210476 149184
rect 243544 149132 243596 149184
rect 125416 149064 125468 149116
rect 216772 149064 216824 149116
rect 239404 148316 239456 148368
rect 256056 148316 256108 148368
rect 67548 147704 67600 147756
rect 112536 147704 112588 147756
rect 167828 147704 167880 147756
rect 168288 147704 168340 147756
rect 202144 147704 202196 147756
rect 206928 147704 206980 147756
rect 320180 147704 320232 147756
rect 100116 147636 100168 147688
rect 100668 147636 100720 147688
rect 227812 147636 227864 147688
rect 214012 147568 214064 147620
rect 256700 147568 256752 147620
rect 257436 147568 257488 147620
rect 210700 147160 210752 147212
rect 214012 147160 214064 147212
rect 3148 147024 3200 147076
rect 95516 147024 95568 147076
rect 96528 147024 96580 147076
rect 83556 146956 83608 147008
rect 90456 146956 90508 147008
rect 169024 146956 169076 147008
rect 184388 146956 184440 147008
rect 193496 146956 193548 147008
rect 207204 146956 207256 147008
rect 90916 146888 90968 146940
rect 127624 146888 127676 146940
rect 220820 146888 220872 146940
rect 257436 146888 257488 146940
rect 580264 146888 580316 146940
rect 213276 146208 213328 146260
rect 216588 146208 216640 146260
rect 244372 146208 244424 146260
rect 244924 146208 244976 146260
rect 197084 145596 197136 145648
rect 213736 145596 213788 145648
rect 8944 145528 8996 145580
rect 87512 145528 87564 145580
rect 114468 145528 114520 145580
rect 180064 145528 180116 145580
rect 218980 145528 219032 145580
rect 267832 145528 267884 145580
rect 282920 145528 282972 145580
rect 298744 145528 298796 145580
rect 160928 144984 160980 145036
rect 161296 144984 161348 145036
rect 193772 144984 193824 145036
rect 192576 144916 192628 144968
rect 244372 144916 244424 144968
rect 87512 144848 87564 144900
rect 125416 144848 125468 144900
rect 160836 144848 160888 144900
rect 184296 144848 184348 144900
rect 97540 144304 97592 144356
rect 99380 144304 99432 144356
rect 185492 144168 185544 144220
rect 193588 144168 193640 144220
rect 173348 144100 173400 144152
rect 180248 144100 180300 144152
rect 186964 143624 187016 143676
rect 226340 143624 226392 143676
rect 66076 143556 66128 143608
rect 91652 143556 91704 143608
rect 224132 143556 224184 143608
rect 224316 143556 224368 143608
rect 313280 143556 313332 143608
rect 208124 143488 208176 143540
rect 209044 143488 209096 143540
rect 69664 142808 69716 142860
rect 83464 142808 83516 142860
rect 86040 142808 86092 142860
rect 86776 142808 86828 142860
rect 215300 142808 215352 142860
rect 216128 142808 216180 142860
rect 217324 142400 217376 142452
rect 218244 142400 218296 142452
rect 220084 142196 220136 142248
rect 228364 142196 228416 142248
rect 78956 142128 79008 142180
rect 206376 142128 206428 142180
rect 213184 142128 213236 142180
rect 232596 142128 232648 142180
rect 80428 141448 80480 141500
rect 103520 141448 103572 141500
rect 104716 141448 104768 141500
rect 70308 141380 70360 141432
rect 105084 141380 105136 141432
rect 173808 141380 173860 141432
rect 200764 141380 200816 141432
rect 203432 140836 203484 140888
rect 289084 140836 289136 140888
rect 104716 140768 104768 140820
rect 207756 140768 207808 140820
rect 215024 140768 215076 140820
rect 255320 140768 255372 140820
rect 71320 140700 71372 140752
rect 73068 140700 73120 140752
rect 189080 140700 189132 140752
rect 218704 140700 218756 140752
rect 221832 140700 221884 140752
rect 64512 140020 64564 140072
rect 70400 140020 70452 140072
rect 184848 139544 184900 139596
rect 198648 140496 198700 140548
rect 67824 139408 67876 139460
rect 100208 139408 100260 139460
rect 210056 140496 210108 140548
rect 205916 140428 205968 140480
rect 206928 140428 206980 140480
rect 218520 140428 218572 140480
rect 222016 140428 222068 140480
rect 225236 140428 225288 140480
rect 264888 140088 264940 140140
rect 276020 140088 276072 140140
rect 287704 140020 287756 140072
rect 225236 139408 225288 139460
rect 264888 139408 264940 139460
rect 52184 138660 52236 138712
rect 72516 138660 72568 138712
rect 90824 138660 90876 138712
rect 163596 138660 163648 138712
rect 87052 138592 87104 138644
rect 278780 139340 278832 139392
rect 280068 139340 280120 139392
rect 280068 138660 280120 138712
rect 322204 138660 322256 138712
rect 78864 138048 78916 138100
rect 79508 138048 79560 138100
rect 3608 137980 3660 138032
rect 75828 137980 75880 138032
rect 3516 137912 3568 137964
rect 72976 137912 73028 137964
rect 78864 137912 78916 137964
rect 79324 137912 79376 137964
rect 77852 137844 77904 137896
rect 81348 137844 81400 137896
rect 69388 137776 69440 137828
rect 75276 137776 75328 137828
rect 79324 137708 79376 137760
rect 184848 137912 184900 137964
rect 101404 137844 101456 137896
rect 102048 137844 102100 137896
rect 192576 137844 192628 137896
rect 229744 137028 229796 137080
rect 237380 137028 237432 137080
rect 89352 136960 89404 137012
rect 90364 136960 90416 137012
rect 83372 136688 83424 136740
rect 86224 136688 86276 136740
rect 81348 136620 81400 136672
rect 83556 136620 83608 136672
rect 85948 136620 86000 136672
rect 87052 136620 87104 136672
rect 90272 136620 90324 136672
rect 91744 136620 91796 136672
rect 92388 136620 92440 136672
rect 93124 136620 93176 136672
rect 91652 136552 91704 136604
rect 166356 136552 166408 136604
rect 184388 136552 184440 136604
rect 191564 136552 191616 136604
rect 11704 135940 11756 135992
rect 91008 135940 91060 135992
rect 69572 135872 69624 135924
rect 160928 135872 160980 135924
rect 180064 135260 180116 135312
rect 191564 135260 191616 135312
rect 75644 135192 75696 135244
rect 94136 135192 94188 135244
rect 96712 135192 96764 135244
rect 145656 135192 145708 135244
rect 188436 135192 188488 135244
rect 192852 135192 192904 135244
rect 227076 135192 227128 135244
rect 227904 135192 227956 135244
rect 267740 135192 267792 135244
rect 68836 134580 68888 134632
rect 74540 134580 74592 134632
rect 75644 134580 75696 134632
rect 226708 134512 226760 134564
rect 278044 134512 278096 134564
rect 94688 133900 94740 133952
rect 130476 133968 130528 134020
rect 181536 133900 181588 133952
rect 193036 133900 193088 133952
rect 226340 133900 226392 133952
rect 127716 133832 127768 133884
rect 182916 133832 182968 133884
rect 226708 133832 226760 133884
rect 229284 133832 229336 133884
rect 269120 133832 269172 133884
rect 273904 133832 273956 133884
rect 96712 133288 96764 133340
rect 102784 133288 102836 133340
rect 53472 133152 53524 133204
rect 66352 133152 66404 133204
rect 153936 133152 153988 133204
rect 187148 133152 187200 133204
rect 50712 132404 50764 132456
rect 66260 132404 66312 132456
rect 96620 132404 96672 132456
rect 186964 132404 187016 132456
rect 226708 132404 226760 132456
rect 238760 132404 238812 132456
rect 142988 132336 143040 132388
rect 191656 132336 191708 132388
rect 104164 131044 104216 131096
rect 156604 131044 156656 131096
rect 188436 131044 188488 131096
rect 226708 131044 226760 131096
rect 230572 131044 230624 131096
rect 276112 131044 276164 131096
rect 96620 130976 96672 131028
rect 135904 130976 135956 131028
rect 97908 129684 97960 129736
rect 177396 129684 177448 129736
rect 226708 129684 226760 129736
rect 266452 129684 266504 129736
rect 267832 129684 267884 129736
rect 96712 129616 96764 129668
rect 115204 129616 115256 129668
rect 118056 129004 118108 129056
rect 169760 129004 169812 129056
rect 226708 129004 226760 129056
rect 299480 129004 299532 129056
rect 169760 128324 169812 128376
rect 171048 128324 171100 128376
rect 191656 128324 191708 128376
rect 61752 128256 61804 128308
rect 66812 128256 66864 128308
rect 100208 128256 100260 128308
rect 181536 128256 181588 128308
rect 226616 128256 226668 128308
rect 245660 128256 245712 128308
rect 97908 128188 97960 128240
rect 151176 128188 151228 128240
rect 245660 127576 245712 127628
rect 323584 127576 323636 127628
rect 54944 126896 54996 126948
rect 66812 126896 66864 126948
rect 94964 126896 95016 126948
rect 180156 126896 180208 126948
rect 188896 126896 188948 126948
rect 191656 126896 191708 126948
rect 226340 126896 226392 126948
rect 252560 126896 252612 126948
rect 253020 126896 253072 126948
rect 97172 126828 97224 126880
rect 105544 126828 105596 126880
rect 226708 126828 226760 126880
rect 234620 126828 234672 126880
rect 105636 126216 105688 126268
rect 155316 126216 155368 126268
rect 253020 126216 253072 126268
rect 349160 126216 349212 126268
rect 57612 125536 57664 125588
rect 66812 125536 66864 125588
rect 97448 125536 97500 125588
rect 173256 125536 173308 125588
rect 257344 125536 257396 125588
rect 280252 125536 280304 125588
rect 281448 125536 281500 125588
rect 156696 125468 156748 125520
rect 190368 125468 190420 125520
rect 226708 125468 226760 125520
rect 259460 125468 259512 125520
rect 64696 124924 64748 124976
rect 66904 124924 66956 124976
rect 281448 124856 281500 124908
rect 316040 124856 316092 124908
rect 61844 124108 61896 124160
rect 66628 124108 66680 124160
rect 94596 124108 94648 124160
rect 184204 124108 184256 124160
rect 226708 124108 226760 124160
rect 236092 124108 236144 124160
rect 287152 124108 287204 124160
rect 582748 124108 582800 124160
rect 178684 124040 178736 124092
rect 190644 124040 190696 124092
rect 232504 123428 232556 123480
rect 255964 123428 256016 123480
rect 187516 122816 187568 122868
rect 191656 122816 191708 122868
rect 46756 122748 46808 122800
rect 66812 122748 66864 122800
rect 97908 122748 97960 122800
rect 116676 122748 116728 122800
rect 226340 122748 226392 122800
rect 251272 122748 251324 122800
rect 182916 122068 182968 122120
rect 183468 122068 183520 122120
rect 191656 122068 191708 122120
rect 60464 121388 60516 121440
rect 66812 121388 66864 121440
rect 97172 121388 97224 121440
rect 153936 121388 153988 121440
rect 226708 121388 226760 121440
rect 233240 121388 233292 121440
rect 60556 121320 60608 121372
rect 66628 121320 66680 121372
rect 170956 120776 171008 120828
rect 184848 120776 184900 120828
rect 102876 120708 102928 120760
rect 183376 120708 183428 120760
rect 232596 120708 232648 120760
rect 295340 120708 295392 120760
rect 96068 120300 96120 120352
rect 98736 120300 98788 120352
rect 183376 120096 183428 120148
rect 188988 120096 189040 120148
rect 56416 120028 56468 120080
rect 66812 120028 66864 120080
rect 158076 120028 158128 120080
rect 187516 120028 187568 120080
rect 188344 120028 188396 120080
rect 191656 120028 191708 120080
rect 226524 119824 226576 119876
rect 229100 119824 229152 119876
rect 3424 119348 3476 119400
rect 53840 119348 53892 119400
rect 112536 119348 112588 119400
rect 184296 119348 184348 119400
rect 233240 119348 233292 119400
rect 260840 119348 260892 119400
rect 98736 118940 98788 118992
rect 103704 118940 103756 118992
rect 97264 118668 97316 118720
rect 100944 118668 100996 118720
rect 186964 118668 187016 118720
rect 187516 118668 187568 118720
rect 97908 118600 97960 118652
rect 108488 118600 108540 118652
rect 226616 118600 226668 118652
rect 231860 118600 231912 118652
rect 233148 118600 233200 118652
rect 53564 118532 53616 118584
rect 66260 118532 66312 118584
rect 97816 118192 97868 118244
rect 105636 118192 105688 118244
rect 233148 117920 233200 117972
rect 304264 117920 304316 117972
rect 63224 117240 63276 117292
rect 66260 117240 66312 117292
rect 97908 117240 97960 117292
rect 169300 117240 169352 117292
rect 184848 117240 184900 117292
rect 191656 117240 191708 117292
rect 63132 117172 63184 117224
rect 66904 117172 66956 117224
rect 97816 117172 97868 117224
rect 148416 117172 148468 117224
rect 226708 116628 226760 116680
rect 233240 116628 233292 116680
rect 226340 116560 226392 116612
rect 258172 116560 258224 116612
rect 188436 116016 188488 116068
rect 190644 116016 190696 116068
rect 50804 115880 50856 115932
rect 66812 115880 66864 115932
rect 97908 115880 97960 115932
rect 187056 115880 187108 115932
rect 97816 115812 97868 115864
rect 173348 115812 173400 115864
rect 226524 115200 226576 115252
rect 229100 115200 229152 115252
rect 273352 115200 273404 115252
rect 62028 114452 62080 114504
rect 66812 114452 66864 114504
rect 53840 113772 53892 113824
rect 62028 113772 62080 113824
rect 66904 113772 66956 113824
rect 228364 113772 228416 113824
rect 252560 113772 252612 113824
rect 97540 113160 97592 113212
rect 187148 113160 187200 113212
rect 188252 113160 188304 113212
rect 191012 113160 191064 113212
rect 227352 113160 227404 113212
rect 244464 113160 244516 113212
rect 157248 112412 157300 112464
rect 191748 112412 191800 112464
rect 97908 111868 97960 111920
rect 153844 111868 153896 111920
rect 156604 111868 156656 111920
rect 157248 111868 157300 111920
rect 97816 111800 97868 111852
rect 177396 111800 177448 111852
rect 238116 111800 238168 111852
rect 324320 111800 324372 111852
rect 3148 111732 3200 111784
rect 11704 111732 11756 111784
rect 225328 111732 225380 111784
rect 241520 111732 241572 111784
rect 57520 111052 57572 111104
rect 66168 111052 66220 111104
rect 66628 111052 66680 111104
rect 96804 111052 96856 111104
rect 100116 111052 100168 111104
rect 226524 111052 226576 111104
rect 240692 111052 240744 111104
rect 291844 111052 291896 111104
rect 184756 110848 184808 110900
rect 190368 110848 190420 110900
rect 187700 110440 187752 110492
rect 191748 110440 191800 110492
rect 97448 110236 97500 110288
rect 100760 110236 100812 110288
rect 55128 109692 55180 109744
rect 60740 109692 60792 109744
rect 116584 109692 116636 109744
rect 188252 109692 188304 109744
rect 226984 109692 227036 109744
rect 262404 109692 262456 109744
rect 60740 109012 60792 109064
rect 61384 109012 61436 109064
rect 66812 109012 66864 109064
rect 97172 109012 97224 109064
rect 160836 109012 160888 109064
rect 187056 109012 187108 109064
rect 191564 109012 191616 109064
rect 59084 108944 59136 108996
rect 66904 108944 66956 108996
rect 160744 108944 160796 108996
rect 187700 108944 187752 108996
rect 97908 108332 97960 108384
rect 109040 108332 109092 108384
rect 109684 108332 109736 108384
rect 225052 108332 225104 108384
rect 225236 108332 225288 108384
rect 230388 108332 230440 108384
rect 244280 108332 244332 108384
rect 95976 108264 96028 108316
rect 107660 108264 107712 108316
rect 173256 108264 173308 108316
rect 233148 108264 233200 108316
rect 288532 108264 288584 108316
rect 225052 108196 225104 108248
rect 225328 108196 225380 108248
rect 187608 107788 187660 107840
rect 189080 107788 189132 107840
rect 191748 107788 191800 107840
rect 226616 107720 226668 107772
rect 229192 107720 229244 107772
rect 230388 107720 230440 107772
rect 63316 107652 63368 107704
rect 66812 107652 66864 107704
rect 226708 107652 226760 107704
rect 231952 107652 232004 107704
rect 233148 107652 233200 107704
rect 52276 107584 52328 107636
rect 66904 107584 66956 107636
rect 162768 107584 162820 107636
rect 191564 107584 191616 107636
rect 50620 106904 50672 106956
rect 59084 106904 59136 106956
rect 97540 106360 97592 106412
rect 101496 106360 101548 106412
rect 59084 106292 59136 106344
rect 66812 106292 66864 106344
rect 97908 106292 97960 106344
rect 184204 106292 184256 106344
rect 226708 106292 226760 106344
rect 230572 106292 230624 106344
rect 353300 106292 353352 106344
rect 97540 106224 97592 106276
rect 120080 106224 120132 106276
rect 184296 105884 184348 105936
rect 191748 105884 191800 105936
rect 166356 105612 166408 105664
rect 190460 105612 190512 105664
rect 48136 105544 48188 105596
rect 65984 105544 66036 105596
rect 66536 105544 66588 105596
rect 97908 105544 97960 105596
rect 100852 105544 100904 105596
rect 180156 105544 180208 105596
rect 226340 105544 226392 105596
rect 270500 105544 270552 105596
rect 270500 105136 270552 105188
rect 271144 105136 271196 105188
rect 59176 104796 59228 104848
rect 66260 104796 66312 104848
rect 226524 104796 226576 104848
rect 244280 104796 244332 104848
rect 97908 104116 97960 104168
rect 106280 104116 106332 104168
rect 180248 104116 180300 104168
rect 191656 104116 191708 104168
rect 244280 104116 244332 104168
rect 284944 104116 284996 104168
rect 97908 103436 97960 103488
rect 134616 103436 134668 103488
rect 162124 103504 162176 103556
rect 97724 103368 97776 103420
rect 101404 103368 101456 103420
rect 64788 102348 64840 102400
rect 66076 102348 66128 102400
rect 66536 102348 66588 102400
rect 188344 102144 188396 102196
rect 191012 102144 191064 102196
rect 226616 102144 226668 102196
rect 231860 102144 231912 102196
rect 269764 102144 269816 102196
rect 226708 102076 226760 102128
rect 266360 102076 266412 102128
rect 98828 101396 98880 101448
rect 160100 101396 160152 101448
rect 187700 101396 187752 101448
rect 59268 101260 59320 101312
rect 61844 101260 61896 101312
rect 66444 101260 66496 101312
rect 187700 100988 187752 101040
rect 188988 100988 189040 101040
rect 190644 100988 190696 101040
rect 53748 100716 53800 100768
rect 57888 100716 57940 100768
rect 66812 100716 66864 100768
rect 97632 100716 97684 100768
rect 169024 100716 169076 100768
rect 175188 100648 175240 100700
rect 190644 100648 190696 100700
rect 57796 99968 57848 100020
rect 64788 99968 64840 100020
rect 66812 99968 66864 100020
rect 227536 99968 227588 100020
rect 227996 99968 228048 100020
rect 247040 99968 247092 100020
rect 327724 99968 327776 100020
rect 97816 99424 97868 99476
rect 128268 99424 128320 99476
rect 97908 99356 97960 99408
rect 173348 99356 173400 99408
rect 61936 99288 61988 99340
rect 66628 99288 66680 99340
rect 97816 99288 97868 99340
rect 132592 99288 132644 99340
rect 133788 99288 133840 99340
rect 226156 99288 226208 99340
rect 287060 99288 287112 99340
rect 288348 99288 288400 99340
rect 97540 99084 97592 99136
rect 99288 99084 99340 99136
rect 100024 99084 100076 99136
rect 133788 98608 133840 98660
rect 178776 98608 178828 98660
rect 288348 98608 288400 98660
rect 331220 98608 331272 98660
rect 188528 98064 188580 98116
rect 191748 98064 191800 98116
rect 225052 98064 225104 98116
rect 101404 97996 101456 98048
rect 190828 97996 190880 98048
rect 226616 97928 226668 97980
rect 232504 97928 232556 97980
rect 225052 97860 225104 97912
rect 96620 97656 96672 97708
rect 98644 97656 98696 97708
rect 57704 97248 57756 97300
rect 66628 97248 66680 97300
rect 100024 97248 100076 97300
rect 188436 97248 188488 97300
rect 226432 96704 226484 96756
rect 226708 96704 226760 96756
rect 3056 96636 3108 96688
rect 57244 96636 57296 96688
rect 97908 96636 97960 96688
rect 184296 96636 184348 96688
rect 226432 96568 226484 96620
rect 262220 96568 262272 96620
rect 226616 96500 226668 96552
rect 240784 96500 240836 96552
rect 97448 95888 97500 95940
rect 169668 95888 169720 95940
rect 186136 95888 186188 95940
rect 191564 95888 191616 95940
rect 264244 95888 264296 95940
rect 280160 95888 280212 95940
rect 97908 95208 97960 95260
rect 191840 95208 191892 95260
rect 97816 95140 97868 95192
rect 114560 95140 114612 95192
rect 226708 94528 226760 94580
rect 240784 94528 240836 94580
rect 106188 94460 106240 94512
rect 188436 94460 188488 94512
rect 226248 94460 226300 94512
rect 245752 94460 245804 94512
rect 166908 93848 166960 93900
rect 184848 93848 184900 93900
rect 191656 93848 191708 93900
rect 63408 93780 63460 93832
rect 67824 93780 67876 93832
rect 95148 93100 95200 93152
rect 165528 93100 165580 93152
rect 178684 93100 178736 93152
rect 249156 93100 249208 93152
rect 262864 93100 262916 93152
rect 68928 92692 68980 92744
rect 69710 92692 69762 92744
rect 72838 92692 72890 92744
rect 72976 92692 73028 92744
rect 94366 92692 94418 92744
rect 95240 92692 95292 92744
rect 90134 92624 90186 92676
rect 91008 92624 91060 92676
rect 74540 92556 74592 92608
rect 75782 92556 75834 92608
rect 48044 92488 48096 92540
rect 70308 92488 70360 92540
rect 107016 92488 107068 92540
rect 107660 92488 107712 92540
rect 185676 92556 185728 92608
rect 179236 92488 179288 92540
rect 195980 92488 196032 92540
rect 224868 92488 224920 92540
rect 242900 92488 242952 92540
rect 67364 92420 67416 92472
rect 188528 92420 188580 92472
rect 193036 92420 193088 92472
rect 202604 92420 202656 92472
rect 204168 92420 204220 92472
rect 206100 92420 206152 92472
rect 67548 92352 67600 92404
rect 166908 92352 166960 92404
rect 166172 91740 166224 91792
rect 223580 91740 223632 91792
rect 64512 90992 64564 91044
rect 70768 90992 70820 91044
rect 84660 90992 84712 91044
rect 100760 90992 100812 91044
rect 179328 90992 179380 91044
rect 211804 90992 211856 91044
rect 222384 91128 222436 91180
rect 227720 91128 227772 91180
rect 224224 91060 224276 91112
rect 225144 91060 225196 91112
rect 172428 90924 172480 90976
rect 194600 90924 194652 90976
rect 217140 90856 217192 90908
rect 222476 90992 222528 91044
rect 241612 90992 241664 91044
rect 242164 90992 242216 91044
rect 221372 90924 221424 90976
rect 226248 90924 226300 90976
rect 46848 90312 46900 90364
rect 67548 90312 67600 90364
rect 68468 90312 68520 90364
rect 93860 90244 93912 90296
rect 95056 90244 95108 90296
rect 95884 90244 95936 90296
rect 206284 89700 206336 89752
rect 207940 89700 207992 89752
rect 67180 89632 67232 89684
rect 101404 89632 101456 89684
rect 111800 89632 111852 89684
rect 112444 89632 112496 89684
rect 209228 89632 209280 89684
rect 214564 89632 214616 89684
rect 258080 89632 258132 89684
rect 75460 89564 75512 89616
rect 95976 89564 96028 89616
rect 215852 89496 215904 89548
rect 239404 89564 239456 89616
rect 209872 88476 209924 88528
rect 210700 88476 210752 88528
rect 69204 88272 69256 88324
rect 158720 88272 158772 88324
rect 193864 88272 193916 88324
rect 194140 88272 194192 88324
rect 204444 88272 204496 88324
rect 208400 88272 208452 88324
rect 211620 88272 211672 88324
rect 263600 88272 263652 88324
rect 80060 88204 80112 88256
rect 95148 88204 95200 88256
rect 178776 88204 178828 88256
rect 224960 88204 225012 88256
rect 73804 86912 73856 86964
rect 167736 86912 167788 86964
rect 62028 86844 62080 86896
rect 100024 86844 100076 86896
rect 188436 86912 188488 86964
rect 226524 86912 226576 86964
rect 285772 86912 285824 86964
rect 580172 86912 580224 86964
rect 199384 86844 199436 86896
rect 220636 86844 220688 86896
rect 253204 86844 253256 86896
rect 3424 85484 3476 85536
rect 61384 85484 61436 85536
rect 116584 85484 116636 85536
rect 124036 85484 124088 85536
rect 215300 85484 215352 85536
rect 67456 85416 67508 85468
rect 97448 85416 97500 85468
rect 173256 85416 173308 85468
rect 201408 85416 201460 85468
rect 201408 84804 201460 84856
rect 214564 84804 214616 84856
rect 216588 84260 216640 84312
rect 266360 84260 266412 84312
rect 222844 84192 222896 84244
rect 342352 84192 342404 84244
rect 71780 84124 71832 84176
rect 102140 84124 102192 84176
rect 196072 84124 196124 84176
rect 73160 84056 73212 84108
rect 161480 84056 161532 84108
rect 162768 84056 162820 84108
rect 191748 82832 191800 82884
rect 248420 82832 248472 82884
rect 75920 82764 75972 82816
rect 107660 82764 107712 82816
rect 153844 82764 153896 82816
rect 244464 82764 244516 82816
rect 92480 82696 92532 82748
rect 122104 82696 122156 82748
rect 185676 82696 185728 82748
rect 203524 82696 203576 82748
rect 203616 82696 203668 82748
rect 284300 82696 284352 82748
rect 284300 82084 284352 82136
rect 582748 82084 582800 82136
rect 244464 81404 244516 81456
rect 244924 81404 244976 81456
rect 63316 81336 63368 81388
rect 159456 81336 159508 81388
rect 173348 81336 173400 81388
rect 227996 81336 228048 81388
rect 77300 81268 77352 81320
rect 108396 81268 108448 81320
rect 191104 80656 191156 80708
rect 280804 80656 280856 80708
rect 64788 79976 64840 80028
rect 191748 79976 191800 80028
rect 85672 79908 85724 79960
rect 104900 79908 104952 79960
rect 162768 79908 162820 79960
rect 198832 79908 198884 79960
rect 198832 79364 198884 79416
rect 240140 79364 240192 79416
rect 240784 79364 240836 79416
rect 241520 79364 241572 79416
rect 211068 79296 211120 79348
rect 582840 79296 582892 79348
rect 87052 78616 87104 78668
rect 216588 78616 216640 78668
rect 80244 78548 80296 78600
rect 177948 78548 178000 78600
rect 206284 78548 206336 78600
rect 207020 77256 207072 77308
rect 208308 77256 208360 77308
rect 246304 77256 246356 77308
rect 95148 77188 95200 77240
rect 222844 77188 222896 77240
rect 61844 77120 61896 77172
rect 100116 77120 100168 77172
rect 109684 77120 109736 77172
rect 227812 77120 227864 77172
rect 66076 75828 66128 75880
rect 180248 75828 180300 75880
rect 177396 75760 177448 75812
rect 229100 75760 229152 75812
rect 75828 75148 75880 75200
rect 171784 75148 171836 75200
rect 190460 75148 190512 75200
rect 207020 75148 207072 75200
rect 59084 74468 59136 74520
rect 187056 74468 187108 74520
rect 180156 74400 180208 74452
rect 230572 74400 230624 74452
rect 89628 73788 89680 73840
rect 173164 73788 173216 73840
rect 58624 73176 58676 73228
rect 59084 73176 59136 73228
rect 169024 73108 169076 73160
rect 227904 73108 227956 73160
rect 178684 73040 178736 73092
rect 205732 73040 205784 73092
rect 86868 72428 86920 72480
rect 170404 72428 170456 72480
rect 211804 72428 211856 72480
rect 356060 72428 356112 72480
rect 205732 71748 205784 71800
rect 206376 71748 206428 71800
rect 227904 71748 227956 71800
rect 228364 71748 228416 71800
rect 3424 71680 3476 71732
rect 95332 71680 95384 71732
rect 128268 71680 128320 71732
rect 226340 71680 226392 71732
rect 93768 71000 93820 71052
rect 157984 71000 158036 71052
rect 183376 71000 183428 71052
rect 191104 71000 191156 71052
rect 192944 71000 192996 71052
rect 281540 71000 281592 71052
rect 226340 70388 226392 70440
rect 226984 70388 227036 70440
rect 162124 70320 162176 70372
rect 231860 70320 231912 70372
rect 96528 69640 96580 69692
rect 164884 69640 164936 69692
rect 190368 69640 190420 69692
rect 250444 69640 250496 69692
rect 89904 68960 89956 69012
rect 220084 68960 220136 69012
rect 80152 68892 80204 68944
rect 190460 68892 190512 68944
rect 193128 68280 193180 68332
rect 327080 68280 327132 68332
rect 91008 67532 91060 67584
rect 218060 67532 218112 67584
rect 67548 66852 67600 66904
rect 99932 66852 99984 66904
rect 81440 66172 81492 66224
rect 208492 66172 208544 66224
rect 209044 66172 209096 66224
rect 86960 66104 87012 66156
rect 115940 66104 115992 66156
rect 215944 66104 215996 66156
rect 93676 64812 93728 64864
rect 241612 64812 241664 64864
rect 74540 64744 74592 64796
rect 201500 64744 201552 64796
rect 201500 63520 201552 63572
rect 202144 63520 202196 63572
rect 241612 63520 241664 63572
rect 242164 63520 242216 63572
rect 71872 63452 71924 63504
rect 198004 63452 198056 63504
rect 218060 63452 218112 63504
rect 277400 63452 277452 63504
rect 278688 63452 278740 63504
rect 278688 62772 278740 62824
rect 351920 62772 351972 62824
rect 85580 62024 85632 62076
rect 212632 62024 212684 62076
rect 212632 60732 212684 60784
rect 213276 60732 213328 60784
rect 88340 60664 88392 60716
rect 222384 60664 222436 60716
rect 222936 60664 222988 60716
rect 193864 59984 193916 60036
rect 264980 59984 265032 60036
rect 99932 59304 99984 59356
rect 193312 59304 193364 59356
rect 193864 59304 193916 59356
rect 57888 58624 57940 58676
rect 181444 58624 181496 58676
rect 82084 57876 82136 57928
rect 210424 57876 210476 57928
rect 84200 57808 84252 57860
rect 118700 57808 118752 57860
rect 213184 57808 213236 57860
rect 73804 56516 73856 56568
rect 200120 56516 200172 56568
rect 200764 56516 200816 56568
rect 77208 54476 77260 54528
rect 152556 54476 152608 54528
rect 193864 54476 193916 54528
rect 291200 54476 291252 54528
rect 101404 53048 101456 53100
rect 137376 53048 137428 53100
rect 184848 53048 184900 53100
rect 292672 53048 292724 53100
rect 186136 51688 186188 51740
rect 328460 51688 328512 51740
rect 55128 50328 55180 50380
rect 141516 50328 141568 50380
rect 180248 50328 180300 50380
rect 269120 50328 269172 50380
rect 73068 48968 73120 49020
rect 149704 48968 149756 49020
rect 188988 48968 189040 49020
rect 251272 48968 251324 49020
rect 68928 47540 68980 47592
rect 175924 47540 175976 47592
rect 204904 47540 204956 47592
rect 343640 47540 343692 47592
rect 189724 46860 189776 46912
rect 580172 46860 580224 46912
rect 3424 45500 3476 45552
rect 57244 45500 57296 45552
rect 59268 44820 59320 44872
rect 144184 44820 144236 44872
rect 171048 44820 171100 44872
rect 332692 44820 332744 44872
rect 181536 43392 181588 43444
rect 222844 43392 222896 43444
rect 226984 43392 227036 43444
rect 277400 43392 277452 43444
rect 61936 42032 61988 42084
rect 138664 42032 138716 42084
rect 222936 42032 222988 42084
rect 290464 42032 290516 42084
rect 186964 40672 187016 40724
rect 338120 40672 338172 40724
rect 46848 39312 46900 39364
rect 163504 39312 163556 39364
rect 206376 38020 206428 38072
rect 213368 38020 213420 38072
rect 213184 37884 213236 37936
rect 333980 37884 334032 37936
rect 66168 36524 66220 36576
rect 140044 36524 140096 36576
rect 203524 36524 203576 36576
rect 324412 36524 324464 36576
rect 213276 35164 213328 35216
rect 287060 35164 287112 35216
rect 67732 33736 67784 33788
rect 125600 33736 125652 33788
rect 193036 33736 193088 33788
rect 270500 33736 270552 33788
rect 2872 33056 2924 33108
rect 54484 33056 54536 33108
rect 200764 32376 200816 32428
rect 340972 32376 341024 32428
rect 79968 31016 80020 31068
rect 151084 31016 151136 31068
rect 210424 31016 210476 31068
rect 322940 31016 322992 31068
rect 53748 29588 53800 29640
rect 145564 29588 145616 29640
rect 183468 29588 183520 29640
rect 249800 29588 249852 29640
rect 70308 28228 70360 28280
rect 142896 28228 142948 28280
rect 199384 28228 199436 28280
rect 244280 28228 244332 28280
rect 250444 28228 250496 28280
rect 288440 28228 288492 28280
rect 86776 26868 86828 26920
rect 167644 26868 167696 26920
rect 243544 26868 243596 26920
rect 259552 26868 259604 26920
rect 84108 25508 84160 25560
rect 147036 25508 147088 25560
rect 39948 24080 40000 24132
rect 170496 24080 170548 24132
rect 121368 22720 121420 22772
rect 126244 22720 126296 22772
rect 202144 22720 202196 22772
rect 321560 22720 321612 22772
rect 91008 21360 91060 21412
rect 146944 21360 146996 21412
rect 191104 21360 191156 21412
rect 307760 21360 307812 21412
rect 3424 20612 3476 20664
rect 69664 20612 69716 20664
rect 100668 19932 100720 19984
rect 166264 19932 166316 19984
rect 204996 19932 205048 19984
rect 320272 19932 320324 19984
rect 78588 18572 78640 18624
rect 177304 18572 177356 18624
rect 215944 18572 215996 18624
rect 284392 18572 284444 18624
rect 271144 16192 271196 16244
rect 276112 16192 276164 16244
rect 244924 15852 244976 15904
rect 261760 15852 261812 15904
rect 106188 13064 106240 13116
rect 141424 13064 141476 13116
rect 206284 13064 206336 13116
rect 274824 13064 274876 13116
rect 284944 13064 284996 13116
rect 330392 13064 330444 13116
rect 95056 11704 95108 11756
rect 134524 11704 134576 11756
rect 195244 11704 195296 11756
rect 312176 11704 312228 11756
rect 332692 11704 332744 11756
rect 333888 11704 333940 11756
rect 198004 10276 198056 10328
rect 342260 10276 342312 10328
rect 278044 8984 278096 9036
rect 315028 8984 315080 9036
rect 209044 8916 209096 8968
rect 279516 8916 279568 8968
rect 141148 7624 141200 7676
rect 180064 7624 180116 7676
rect 224868 7624 224920 7676
rect 254676 7624 254728 7676
rect 572 7556 624 7608
rect 97264 7556 97316 7608
rect 97448 7556 97500 7608
rect 142804 7556 142856 7608
rect 195980 7556 196032 7608
rect 258264 7556 258316 7608
rect 269764 7556 269816 7608
rect 317328 7556 317380 7608
rect 3424 6808 3476 6860
rect 58624 6808 58676 6860
rect 222844 6196 222896 6248
rect 244096 6196 244148 6248
rect 298744 6196 298796 6248
rect 310244 6196 310296 6248
rect 56048 6128 56100 6180
rect 159364 6128 159416 6180
rect 242164 6128 242216 6180
rect 303160 6128 303212 6180
rect 309784 5516 309836 5568
rect 311440 5516 311492 5568
rect 348056 5516 348108 5568
rect 349160 5516 349212 5568
rect 130384 4768 130436 4820
rect 136456 4768 136508 4820
rect 228364 4768 228416 4820
rect 239312 4768 239364 4820
rect 304264 4768 304316 4820
rect 307944 4768 307996 4820
rect 323584 4768 323636 4820
rect 337476 4768 337528 4820
rect 291844 4428 291896 4480
rect 297272 4428 297324 4480
rect 346952 4156 347004 4208
rect 353300 4156 353352 4208
rect 6828 4088 6880 4140
rect 7656 4088 7708 4140
rect 351644 4088 351696 4140
rect 356060 4088 356112 4140
rect 322204 3952 322256 4004
rect 326804 3952 326856 4004
rect 1308 3544 1360 3596
rect 2872 3544 2924 3596
rect 52552 3544 52604 3596
rect 53656 3544 53708 3596
rect 60832 3544 60884 3596
rect 61936 3544 61988 3596
rect 69112 3544 69164 3596
rect 70216 3544 70268 3596
rect 80888 3544 80940 3596
rect 83464 3544 83516 3596
rect 105728 3544 105780 3596
rect 106188 3544 106240 3596
rect 122288 3544 122340 3596
rect 122748 3544 122800 3596
rect 123484 3544 123536 3596
rect 124128 3544 124180 3596
rect 124680 3544 124732 3596
rect 125508 3544 125560 3596
rect 251180 3544 251232 3596
rect 252376 3544 252428 3596
rect 276020 3544 276072 3596
rect 277124 3544 277176 3596
rect 1676 3476 1728 3528
rect 2688 3476 2740 3528
rect 9956 3476 10008 3528
rect 10968 3476 11020 3528
rect 11152 3476 11204 3528
rect 12256 3476 12308 3528
rect 17040 3476 17092 3528
rect 17868 3476 17920 3528
rect 18236 3476 18288 3528
rect 19248 3476 19300 3528
rect 20628 3476 20680 3528
rect 21364 3476 21416 3528
rect 24216 3476 24268 3528
rect 24768 3476 24820 3528
rect 26516 3476 26568 3528
rect 27528 3476 27580 3528
rect 32404 3476 32456 3528
rect 33048 3476 33100 3528
rect 33600 3476 33652 3528
rect 34428 3476 34480 3528
rect 34796 3476 34848 3528
rect 35808 3476 35860 3528
rect 35992 3476 36044 3528
rect 37096 3476 37148 3528
rect 40684 3476 40736 3528
rect 41328 3476 41380 3528
rect 41880 3476 41932 3528
rect 42708 3476 42760 3528
rect 43076 3476 43128 3528
rect 44088 3476 44140 3528
rect 44272 3476 44324 3528
rect 45376 3476 45428 3528
rect 48964 3476 49016 3528
rect 49516 3476 49568 3528
rect 50160 3476 50212 3528
rect 50896 3476 50948 3528
rect 57244 3476 57296 3528
rect 57888 3476 57940 3528
rect 58440 3476 58492 3528
rect 59268 3476 59320 3528
rect 59636 3476 59688 3528
rect 60648 3476 60700 3528
rect 64328 3476 64380 3528
rect 64788 3476 64840 3528
rect 65524 3476 65576 3528
rect 66168 3476 66220 3528
rect 67916 3476 67968 3528
rect 68928 3476 68980 3528
rect 72608 3476 72660 3528
rect 73068 3476 73120 3528
rect 75000 3476 75052 3528
rect 75828 3476 75880 3528
rect 76196 3476 76248 3528
rect 77208 3476 77260 3528
rect 83280 3476 83332 3528
rect 84108 3476 84160 3528
rect 84476 3476 84528 3528
rect 85488 3476 85540 3528
rect 85672 3476 85724 3528
rect 86776 3476 86828 3528
rect 89168 3476 89220 3528
rect 89628 3476 89680 3528
rect 90364 3476 90416 3528
rect 91008 3476 91060 3528
rect 92756 3476 92808 3528
rect 93768 3476 93820 3528
rect 93952 3476 94004 3528
rect 95056 3476 95108 3528
rect 98644 3476 98696 3528
rect 99288 3476 99340 3528
rect 99840 3476 99892 3528
rect 100668 3476 100720 3528
rect 102232 3476 102284 3528
rect 106832 3476 106884 3528
rect 106924 3476 106976 3528
rect 107568 3476 107620 3528
rect 6460 3408 6512 3460
rect 31024 3408 31076 3460
rect 31300 3408 31352 3460
rect 39304 3408 39356 3460
rect 66720 3408 66772 3460
rect 90272 3408 90324 3460
rect 91560 3408 91612 3460
rect 108304 3476 108356 3528
rect 110512 3476 110564 3528
rect 111708 3476 111760 3528
rect 108120 3408 108172 3460
rect 137284 3476 137336 3528
rect 140044 3476 140096 3528
rect 141148 3476 141200 3528
rect 143540 3476 143592 3528
rect 144828 3476 144880 3528
rect 238024 3476 238076 3528
rect 260656 3476 260708 3528
rect 287704 3476 287756 3528
rect 290188 3476 290240 3528
rect 290464 3476 290516 3528
rect 294880 3476 294932 3528
rect 299480 3476 299532 3528
rect 300768 3476 300820 3528
rect 304908 3476 304960 3528
rect 305552 3476 305604 3528
rect 307760 3476 307812 3528
rect 309048 3476 309100 3528
rect 319720 3476 319772 3528
rect 320180 3476 320232 3528
rect 324320 3476 324372 3528
rect 325608 3476 325660 3528
rect 340144 3476 340196 3528
rect 342168 3476 342220 3528
rect 114008 3408 114060 3460
rect 114468 3408 114520 3460
rect 115204 3408 115256 3460
rect 115848 3408 115900 3460
rect 116400 3408 116452 3460
rect 117228 3408 117280 3460
rect 117596 3408 117648 3460
rect 118608 3408 118660 3460
rect 118792 3408 118844 3460
rect 155224 3408 155276 3460
rect 213368 3408 213420 3460
rect 242900 3408 242952 3460
rect 246304 3408 246356 3460
rect 247592 3408 247644 3460
rect 257068 3408 257120 3460
rect 258172 3408 258224 3460
rect 260104 3408 260156 3460
rect 272432 3408 272484 3460
rect 273904 3408 273956 3460
rect 283104 3408 283156 3460
rect 295984 3408 296036 3460
rect 301964 3408 302016 3460
rect 341524 3408 341576 3460
rect 350448 3408 350500 3460
rect 262864 3272 262916 3324
rect 267740 3272 267792 3324
rect 268476 3272 268528 3324
rect 273628 3272 273680 3324
rect 280804 3272 280856 3324
rect 284300 3272 284352 3324
rect 25320 3136 25372 3188
rect 26148 3136 26200 3188
rect 349252 3136 349304 3188
rect 351920 3136 351972 3188
rect 27712 3068 27764 3120
rect 29644 3068 29696 3120
rect 299664 3068 299716 3120
rect 302240 3068 302292 3120
rect 77392 3000 77444 3052
rect 79324 3000 79376 3052
rect 289084 2932 289136 2984
rect 292580 2932 292632 2984
rect 327724 2932 327776 2984
rect 332692 2932 332744 2984
rect 339868 2932 339920 2984
rect 342352 2932 342404 2984
rect 581000 2932 581052 2984
rect 583116 2932 583168 2984
rect 15936 2864 15988 2916
rect 16488 2864 16540 2916
rect 51356 2048 51408 2100
rect 101404 2048 101456 2100
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 8128 702642 8156 703520
rect 24320 702778 24348 703520
rect 24308 702772 24360 702778
rect 24308 702714 24360 702720
rect 8116 702636 8168 702642
rect 8116 702578 8168 702584
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 2778 606112 2834 606121
rect 2778 606047 2834 606056
rect 2792 605946 2820 606047
rect 2780 605940 2832 605946
rect 2780 605882 2832 605888
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 3436 568546 3464 684247
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 17224 670744 17276 670750
rect 17224 670686 17276 670692
rect 3514 658200 3570 658209
rect 3514 658135 3570 658144
rect 3528 656946 3556 658135
rect 3516 656940 3568 656946
rect 3516 656882 3568 656888
rect 15844 656940 15896 656946
rect 15844 656882 15896 656888
rect 3516 632120 3568 632126
rect 3514 632088 3516 632097
rect 3568 632088 3570 632097
rect 3514 632023 3570 632032
rect 15856 621625 15884 656882
rect 15842 621616 15898 621625
rect 15842 621551 15898 621560
rect 3514 619168 3570 619177
rect 3514 619103 3570 619112
rect 3528 618322 3556 619103
rect 3516 618316 3568 618322
rect 3516 618258 3568 618264
rect 4804 605940 4856 605946
rect 4804 605882 4856 605888
rect 4816 587178 4844 605882
rect 4804 587172 4856 587178
rect 4804 587114 4856 587120
rect 3424 568540 3476 568546
rect 3424 568482 3476 568488
rect 4804 568540 4856 568546
rect 4804 568482 4856 568488
rect 3422 566944 3478 566953
rect 3422 566879 3478 566888
rect 3436 540258 3464 566879
rect 3514 553888 3570 553897
rect 3514 553823 3516 553832
rect 3568 553823 3570 553832
rect 3516 553794 3568 553800
rect 4816 542473 4844 568482
rect 7564 553852 7616 553858
rect 7564 553794 7616 553800
rect 4802 542464 4858 542473
rect 4802 542399 4858 542408
rect 3424 540252 3476 540258
rect 3424 540194 3476 540200
rect 7576 538218 7604 553794
rect 17236 541113 17264 670686
rect 21364 632120 21416 632126
rect 21364 632062 21416 632068
rect 21376 576162 21404 632062
rect 40052 588606 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 136652 703582 137692 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 70308 703316 70360 703322
rect 70308 703258 70360 703264
rect 67640 703044 67692 703050
rect 67640 702986 67692 702992
rect 61936 702908 61988 702914
rect 61936 702850 61988 702856
rect 57796 702568 57848 702574
rect 57796 702510 57848 702516
rect 43444 618316 43496 618322
rect 43444 618258 43496 618264
rect 40040 588600 40092 588606
rect 40040 588542 40092 588548
rect 21364 576156 21416 576162
rect 21364 576098 21416 576104
rect 31760 576156 31812 576162
rect 31760 576098 31812 576104
rect 31772 575550 31800 576098
rect 31760 575544 31812 575550
rect 31760 575486 31812 575492
rect 33048 575544 33100 575550
rect 33048 575486 33100 575492
rect 17222 541104 17278 541113
rect 17222 541039 17278 541048
rect 15844 538280 15896 538286
rect 15844 538222 15896 538228
rect 7564 538212 7616 538218
rect 7564 538154 7616 538160
rect 3424 534744 3476 534750
rect 3424 534686 3476 534692
rect 3436 501809 3464 534686
rect 3514 527912 3570 527921
rect 3514 527847 3516 527856
rect 3568 527847 3570 527856
rect 3516 527818 3568 527824
rect 3514 514856 3570 514865
rect 3514 514791 3516 514800
rect 3568 514791 3570 514800
rect 3516 514762 3568 514768
rect 3422 501800 3478 501809
rect 3422 501735 3478 501744
rect 15856 478174 15884 538222
rect 3424 478168 3476 478174
rect 3424 478110 3476 478116
rect 15844 478168 15896 478174
rect 15844 478110 15896 478116
rect 3436 475697 3464 478110
rect 3422 475688 3478 475697
rect 3422 475623 3478 475632
rect 3146 449576 3202 449585
rect 3146 449511 3202 449520
rect 3160 448594 3188 449511
rect 3148 448588 3200 448594
rect 3148 448530 3200 448536
rect 2780 423632 2832 423638
rect 2778 423600 2780 423609
rect 2832 423600 2834 423609
rect 2778 423535 2834 423544
rect 2870 410544 2926 410553
rect 2870 410479 2926 410488
rect 2884 409902 2912 410479
rect 2872 409896 2924 409902
rect 2872 409838 2924 409844
rect 3436 391270 3464 475623
rect 3514 462632 3570 462641
rect 3514 462567 3570 462576
rect 3528 462398 3556 462567
rect 3516 462392 3568 462398
rect 3516 462334 3568 462340
rect 14464 462392 14516 462398
rect 14464 462334 14516 462340
rect 4804 434784 4856 434790
rect 4804 434726 4856 434732
rect 4816 423638 4844 434726
rect 4804 423632 4856 423638
rect 4804 423574 4856 423580
rect 3516 397588 3568 397594
rect 3516 397530 3568 397536
rect 3528 397497 3556 397530
rect 11704 397520 11756 397526
rect 3514 397488 3570 397497
rect 11704 397462 11756 397468
rect 3514 397423 3570 397432
rect 3424 391264 3476 391270
rect 3424 391206 3476 391212
rect 3422 371376 3478 371385
rect 3422 371311 3478 371320
rect 3436 371278 3464 371311
rect 3424 371272 3476 371278
rect 3424 371214 3476 371220
rect 11716 358766 11744 397462
rect 14476 388793 14504 462334
rect 32956 418192 33008 418198
rect 32956 418134 33008 418140
rect 21364 397588 21416 397594
rect 21364 397530 21416 397536
rect 14462 388784 14518 388793
rect 14462 388719 14518 388728
rect 21376 380866 21404 397530
rect 21364 380860 21416 380866
rect 21364 380802 21416 380808
rect 3332 358760 3384 358766
rect 3332 358702 3384 358708
rect 11704 358760 11756 358766
rect 11704 358702 11756 358708
rect 3344 358465 3372 358702
rect 3330 358456 3386 358465
rect 3330 358391 3386 358400
rect 3424 355360 3476 355366
rect 3424 355302 3476 355308
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 3344 345098 3372 345335
rect 3332 345092 3384 345098
rect 3332 345034 3384 345040
rect 3436 319297 3464 355302
rect 18604 345092 18656 345098
rect 18604 345034 18656 345040
rect 12346 328536 12402 328545
rect 12346 328471 12402 328480
rect 3422 319288 3478 319297
rect 3422 319223 3478 319232
rect 3436 313274 3464 319223
rect 3424 313268 3476 313274
rect 3424 313210 3476 313216
rect 7564 313268 7616 313274
rect 7564 313210 7616 313216
rect 1306 306776 1362 306785
rect 1306 306711 1362 306720
rect 572 7608 624 7614
rect 572 7550 624 7556
rect 584 480 612 7550
rect 1320 3602 1348 306711
rect 3238 306232 3294 306241
rect 3238 306167 3294 306176
rect 3252 305046 3280 306167
rect 3240 305040 3292 305046
rect 3240 304982 3292 304988
rect 4066 297392 4122 297401
rect 4066 297327 4122 297336
rect 3422 293176 3478 293185
rect 3422 293111 3478 293120
rect 3436 292602 3464 293111
rect 3424 292596 3476 292602
rect 3424 292538 3476 292544
rect 3516 267708 3568 267714
rect 3516 267650 3568 267656
rect 3528 267209 3556 267650
rect 3514 267200 3570 267209
rect 3514 267135 3570 267144
rect 3424 263628 3476 263634
rect 3424 263570 3476 263576
rect 3148 255264 3200 255270
rect 3148 255206 3200 255212
rect 3160 254153 3188 255206
rect 3146 254144 3202 254153
rect 3146 254079 3202 254088
rect 3436 214985 3464 263570
rect 3516 241256 3568 241262
rect 3516 241198 3568 241204
rect 3528 241097 3556 241198
rect 3514 241088 3570 241097
rect 3514 241023 3570 241032
rect 3422 214976 3478 214985
rect 3422 214911 3478 214920
rect 3332 202224 3384 202230
rect 3332 202166 3384 202172
rect 3344 201929 3372 202166
rect 3330 201920 3386 201929
rect 3330 201855 3386 201864
rect 2688 192500 2740 192506
rect 2688 192442 2740 192448
rect 1308 3596 1360 3602
rect 1308 3538 1360 3544
rect 2700 3534 2728 192442
rect 3146 149832 3202 149841
rect 3146 149767 3202 149776
rect 3160 147082 3188 149767
rect 3148 147076 3200 147082
rect 3148 147018 3200 147024
rect 3436 119406 3464 214911
rect 3516 189032 3568 189038
rect 3516 188974 3568 188980
rect 3528 188873 3556 188974
rect 3514 188864 3570 188873
rect 3514 188799 3570 188808
rect 3516 162920 3568 162926
rect 3514 162888 3516 162897
rect 3568 162888 3570 162897
rect 3514 162823 3570 162832
rect 3608 138032 3660 138038
rect 3608 137974 3660 137980
rect 3516 137964 3568 137970
rect 3516 137906 3568 137912
rect 3528 136785 3556 137906
rect 3514 136776 3570 136785
rect 3514 136711 3570 136720
rect 3620 122834 3648 137974
rect 3528 122806 3648 122834
rect 3424 119400 3476 119406
rect 3424 119342 3476 119348
rect 3148 111784 3200 111790
rect 3148 111726 3200 111732
rect 3160 110673 3188 111726
rect 3146 110664 3202 110673
rect 3146 110599 3202 110608
rect 3054 97608 3110 97617
rect 3054 97543 3110 97552
rect 3068 96694 3096 97543
rect 3056 96688 3108 96694
rect 3056 96630 3108 96636
rect 3424 85536 3476 85542
rect 3424 85478 3476 85484
rect 3436 84697 3464 85478
rect 3422 84688 3478 84697
rect 3422 84623 3478 84632
rect 3424 71732 3476 71738
rect 3424 71674 3476 71680
rect 3436 71641 3464 71674
rect 3422 71632 3478 71641
rect 3422 71567 3478 71576
rect 3528 58585 3556 122806
rect 3514 58576 3570 58585
rect 3514 58511 3570 58520
rect 3424 45552 3476 45558
rect 3422 45520 3424 45529
rect 3476 45520 3478 45529
rect 3422 45455 3478 45464
rect 2872 33108 2924 33114
rect 2872 33050 2924 33056
rect 2884 32473 2912 33050
rect 2870 32464 2926 32473
rect 2870 32399 2926 32408
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 2872 3596 2924 3602
rect 2872 3538 2924 3544
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 2688 3528 2740 3534
rect 2688 3470 2740 3476
rect 1688 480 1716 3470
rect 2884 480 2912 3538
rect 4080 480 4108 297327
rect 7576 279478 7604 313210
rect 12254 298888 12310 298897
rect 12254 298823 12310 298832
rect 10324 280220 10376 280226
rect 10324 280162 10376 280168
rect 7564 279472 7616 279478
rect 7564 279414 7616 279420
rect 7564 262880 7616 262886
rect 7564 262822 7616 262828
rect 7576 241262 7604 262822
rect 10336 255270 10364 280162
rect 10324 255264 10376 255270
rect 10324 255206 10376 255212
rect 7564 241256 7616 241262
rect 7564 241198 7616 241204
rect 5446 196616 5502 196625
rect 5446 196551 5502 196560
rect 5460 6914 5488 196551
rect 6828 185632 6880 185638
rect 6828 185574 6880 185580
rect 5276 6886 5488 6914
rect 5276 480 5304 6886
rect 6840 4146 6868 185574
rect 10968 182844 11020 182850
rect 10968 182786 11020 182792
rect 8944 162920 8996 162926
rect 8944 162862 8996 162868
rect 8956 145586 8984 162862
rect 8944 145580 8996 145586
rect 8944 145522 8996 145528
rect 6828 4140 6880 4146
rect 6828 4082 6880 4088
rect 7656 4140 7708 4146
rect 7656 4082 7708 4088
rect 6460 3460 6512 3466
rect 6460 3402 6512 3408
rect 6472 480 6500 3402
rect 7668 480 7696 4082
rect 10980 3534 11008 182786
rect 11704 135992 11756 135998
rect 11704 135934 11756 135940
rect 11716 111790 11744 135934
rect 11704 111784 11756 111790
rect 11704 111726 11756 111732
rect 12268 3534 12296 298823
rect 9956 3528 10008 3534
rect 9956 3470 10008 3476
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 11152 3528 11204 3534
rect 11152 3470 11204 3476
rect 12256 3528 12308 3534
rect 12256 3470 12308 3476
rect 8758 3360 8814 3369
rect 8758 3295 8814 3304
rect 8772 480 8800 3295
rect 9968 480 9996 3470
rect 11164 480 11192 3470
rect 12360 480 12388 328471
rect 17866 309224 17922 309233
rect 17866 309159 17922 309168
rect 16486 301336 16542 301345
rect 16486 301271 16542 301280
rect 15106 235240 15162 235249
rect 15106 235175 15162 235184
rect 13726 226944 13782 226953
rect 13726 226879 13782 226888
rect 13740 6914 13768 226879
rect 15120 6914 15148 235175
rect 13556 6886 13768 6914
rect 14752 6886 15148 6914
rect 13556 480 13584 6886
rect 14752 480 14780 6886
rect 16500 2922 16528 301271
rect 17880 3534 17908 309159
rect 18616 288386 18644 345034
rect 23388 338156 23440 338162
rect 23388 338098 23440 338104
rect 22008 307828 22060 307834
rect 22008 307770 22060 307776
rect 18696 292596 18748 292602
rect 18696 292538 18748 292544
rect 18604 288380 18656 288386
rect 18604 288322 18656 288328
rect 18708 241233 18736 292538
rect 18694 241224 18750 241233
rect 18694 241159 18750 241168
rect 21362 236056 21418 236065
rect 21362 235991 21418 236000
rect 18602 233472 18658 233481
rect 18602 233407 18658 233416
rect 18616 189038 18644 233407
rect 19246 211848 19302 211857
rect 19246 211783 19302 211792
rect 18604 189032 18656 189038
rect 18604 188974 18656 188980
rect 19260 3534 19288 211783
rect 19430 4856 19486 4865
rect 19430 4791 19486 4800
rect 17040 3528 17092 3534
rect 17040 3470 17092 3476
rect 17868 3528 17920 3534
rect 17868 3470 17920 3476
rect 18236 3528 18288 3534
rect 18236 3470 18288 3476
rect 19248 3528 19300 3534
rect 19248 3470 19300 3476
rect 15936 2916 15988 2922
rect 15936 2858 15988 2864
rect 16488 2916 16540 2922
rect 16488 2858 16540 2864
rect 15948 480 15976 2858
rect 17052 480 17080 3470
rect 18248 480 18276 3470
rect 19444 480 19472 4791
rect 21376 3534 21404 235991
rect 22020 6914 22048 307770
rect 23400 6914 23428 338098
rect 30286 311944 30342 311953
rect 30286 311879 30342 311888
rect 26146 294536 26202 294545
rect 26146 294471 26202 294480
rect 24766 221504 24822 221513
rect 24766 221439 24822 221448
rect 21836 6886 22048 6914
rect 23032 6886 23428 6914
rect 20628 3528 20680 3534
rect 20628 3470 20680 3476
rect 21364 3528 21416 3534
rect 21364 3470 21416 3476
rect 20640 480 20668 3470
rect 21836 480 21864 6886
rect 23032 480 23060 6886
rect 24780 3534 24808 221439
rect 24216 3528 24268 3534
rect 24216 3470 24268 3476
rect 24768 3528 24820 3534
rect 24768 3470 24820 3476
rect 24228 480 24256 3470
rect 26160 3194 26188 294471
rect 28906 232520 28962 232529
rect 28906 232455 28962 232464
rect 27528 186992 27580 186998
rect 27528 186934 27580 186940
rect 27540 3534 27568 186934
rect 26516 3528 26568 3534
rect 26516 3470 26568 3476
rect 27528 3528 27580 3534
rect 27528 3470 27580 3476
rect 25320 3188 25372 3194
rect 25320 3130 25372 3136
rect 26148 3188 26200 3194
rect 26148 3130 26200 3136
rect 25332 480 25360 3130
rect 26528 480 26556 3470
rect 27712 3120 27764 3126
rect 27712 3062 27764 3068
rect 27724 480 27752 3062
rect 28920 480 28948 232455
rect 29642 224224 29698 224233
rect 29642 224159 29698 224168
rect 29656 3126 29684 224159
rect 30300 6914 30328 311879
rect 32404 305040 32456 305046
rect 32404 304982 32456 304988
rect 31022 302832 31078 302841
rect 31022 302767 31078 302776
rect 30116 6886 30328 6914
rect 29644 3120 29696 3126
rect 29644 3062 29696 3068
rect 30116 480 30144 6886
rect 31036 3466 31064 302767
rect 32416 253881 32444 304982
rect 32968 262886 32996 418134
rect 33060 377466 33088 575486
rect 41328 564460 41380 564466
rect 41328 564402 41380 564408
rect 34520 540252 34572 540258
rect 34520 540194 34572 540200
rect 34532 539646 34560 540194
rect 34520 539640 34572 539646
rect 34520 539582 34572 539588
rect 35716 539640 35768 539646
rect 35716 539582 35768 539588
rect 33784 436144 33836 436150
rect 33784 436086 33836 436092
rect 33048 377460 33100 377466
rect 33048 377402 33100 377408
rect 33796 355366 33824 436086
rect 35728 396778 35756 539582
rect 39854 531992 39910 532001
rect 39854 531927 39910 531936
rect 36544 448588 36596 448594
rect 36544 448530 36596 448536
rect 35808 407788 35860 407794
rect 35808 407730 35860 407736
rect 35716 396772 35768 396778
rect 35716 396714 35768 396720
rect 33784 355360 33836 355366
rect 33784 355302 33836 355308
rect 35162 313440 35218 313449
rect 35162 313375 35218 313384
rect 34426 310584 34482 310593
rect 34426 310519 34482 310528
rect 34336 279472 34388 279478
rect 34336 279414 34388 279420
rect 32956 262880 33008 262886
rect 32956 262822 33008 262828
rect 32402 253872 32458 253881
rect 32402 253807 32458 253816
rect 33048 209092 33100 209098
rect 33048 209034 33100 209040
rect 33060 3534 33088 209034
rect 34348 160750 34376 279414
rect 34336 160744 34388 160750
rect 34336 160686 34388 160692
rect 34440 3534 34468 310519
rect 32404 3528 32456 3534
rect 32404 3470 32456 3476
rect 33048 3528 33100 3534
rect 33048 3470 33100 3476
rect 33600 3528 33652 3534
rect 33600 3470 33652 3476
rect 34428 3528 34480 3534
rect 34428 3470 34480 3476
rect 34796 3528 34848 3534
rect 34796 3470 34848 3476
rect 31024 3460 31076 3466
rect 31024 3402 31076 3408
rect 31300 3460 31352 3466
rect 31300 3402 31352 3408
rect 31312 480 31340 3402
rect 32416 480 32444 3470
rect 33612 480 33640 3470
rect 34808 480 34836 3470
rect 35176 3369 35204 313375
rect 35820 254561 35848 407730
rect 36556 389230 36584 448530
rect 39868 408474 39896 531927
rect 40684 514820 40736 514826
rect 40684 514762 40736 514768
rect 40696 442950 40724 514762
rect 40684 442944 40736 442950
rect 40684 442886 40736 442892
rect 41236 421592 41288 421598
rect 41236 421534 41288 421540
rect 39948 409148 40000 409154
rect 39948 409090 40000 409096
rect 39856 408468 39908 408474
rect 39856 408410 39908 408416
rect 39868 407794 39896 408410
rect 39856 407788 39908 407794
rect 39856 407730 39908 407736
rect 36544 389224 36596 389230
rect 36544 389166 36596 389172
rect 39302 314800 39358 314809
rect 39302 314735 39358 314744
rect 37186 310720 37242 310729
rect 37186 310655 37242 310664
rect 36544 292596 36596 292602
rect 36544 292538 36596 292544
rect 36556 267714 36584 292538
rect 36544 267708 36596 267714
rect 36544 267650 36596 267656
rect 35806 254552 35862 254561
rect 35806 254487 35862 254496
rect 35806 222864 35862 222873
rect 35806 222799 35862 222808
rect 35820 3534 35848 222799
rect 37096 202156 37148 202162
rect 37096 202098 37148 202104
rect 37108 3534 37136 202098
rect 35808 3528 35860 3534
rect 35808 3470 35860 3476
rect 35992 3528 36044 3534
rect 35992 3470 36044 3476
rect 37096 3528 37148 3534
rect 37096 3470 37148 3476
rect 35162 3360 35218 3369
rect 35162 3295 35218 3304
rect 36004 480 36032 3470
rect 37200 480 37228 310655
rect 38568 198008 38620 198014
rect 38568 197950 38620 197956
rect 38580 6914 38608 197950
rect 38396 6886 38608 6914
rect 38396 480 38424 6886
rect 39316 3466 39344 314735
rect 39854 269784 39910 269793
rect 39854 269719 39910 269728
rect 39868 153882 39896 269719
rect 39960 256018 39988 409090
rect 41248 265674 41276 421534
rect 41340 391338 41368 564402
rect 43456 536790 43484 618258
rect 55128 585200 55180 585206
rect 55128 585142 55180 585148
rect 52368 582412 52420 582418
rect 52368 582354 52420 582360
rect 50988 581052 51040 581058
rect 50988 580994 51040 581000
rect 48136 563712 48188 563718
rect 48136 563654 48188 563660
rect 48044 549296 48096 549302
rect 48044 549238 48096 549244
rect 43444 536784 43496 536790
rect 43444 536726 43496 536732
rect 43994 530632 44050 530641
rect 43994 530567 44050 530576
rect 42708 396840 42760 396846
rect 42708 396782 42760 396788
rect 41328 391332 41380 391338
rect 41328 391274 41380 391280
rect 41328 374672 41380 374678
rect 41328 374614 41380 374620
rect 41236 265668 41288 265674
rect 41236 265610 41288 265616
rect 39948 256012 40000 256018
rect 39948 255954 40000 255960
rect 41234 242992 41290 243001
rect 41234 242927 41290 242936
rect 39856 153876 39908 153882
rect 39856 153818 39908 153824
rect 39868 151814 39896 153818
rect 39868 151786 39988 151814
rect 39960 120737 39988 151786
rect 39946 120728 40002 120737
rect 39946 120663 40002 120672
rect 41248 91769 41276 242927
rect 41340 238746 41368 374614
rect 42720 248402 42748 396782
rect 44008 393990 44036 530567
rect 44088 423700 44140 423706
rect 44088 423642 44140 423648
rect 43996 393984 44048 393990
rect 43996 393926 44048 393932
rect 43996 378820 44048 378826
rect 43996 378762 44048 378768
rect 42708 248396 42760 248402
rect 42708 248338 42760 248344
rect 41328 238740 41380 238746
rect 41328 238682 41380 238688
rect 44008 235278 44036 378762
rect 44100 268394 44128 423642
rect 46848 413296 46900 413302
rect 46848 413238 46900 413244
rect 46756 388748 46808 388754
rect 46756 388690 46808 388696
rect 45468 381540 45520 381546
rect 45468 381482 45520 381488
rect 45376 288516 45428 288522
rect 45376 288458 45428 288464
rect 44088 268388 44140 268394
rect 44088 268330 44140 268336
rect 43996 235272 44048 235278
rect 43996 235214 44048 235220
rect 42706 218648 42762 218657
rect 42706 218583 42762 218592
rect 41326 204912 41382 204921
rect 41326 204847 41382 204856
rect 41234 91760 41290 91769
rect 41234 91695 41290 91704
rect 39948 24132 40000 24138
rect 39948 24074 40000 24080
rect 39960 6914 39988 24074
rect 39592 6886 39988 6914
rect 39304 3460 39356 3466
rect 39304 3402 39356 3408
rect 39592 480 39620 6886
rect 41340 3534 41368 204847
rect 42720 3534 42748 218583
rect 44088 207664 44140 207670
rect 44088 207606 44140 207612
rect 44100 3534 44128 207606
rect 45388 199442 45416 288458
rect 45480 240038 45508 381482
rect 46664 272536 46716 272542
rect 46664 272478 46716 272484
rect 45468 240032 45520 240038
rect 45468 239974 45520 239980
rect 45466 210352 45522 210361
rect 45466 210287 45522 210296
rect 45376 199436 45428 199442
rect 45376 199378 45428 199384
rect 45374 199336 45430 199345
rect 45374 199271 45430 199280
rect 45388 3534 45416 199271
rect 40684 3528 40736 3534
rect 40684 3470 40736 3476
rect 41328 3528 41380 3534
rect 41328 3470 41380 3476
rect 41880 3528 41932 3534
rect 41880 3470 41932 3476
rect 42708 3528 42760 3534
rect 42708 3470 42760 3476
rect 43076 3528 43128 3534
rect 43076 3470 43128 3476
rect 44088 3528 44140 3534
rect 44088 3470 44140 3476
rect 44272 3528 44324 3534
rect 44272 3470 44324 3476
rect 45376 3528 45428 3534
rect 45376 3470 45428 3476
rect 40696 480 40724 3470
rect 41892 480 41920 3470
rect 43088 480 43116 3470
rect 44284 480 44312 3470
rect 45480 480 45508 210287
rect 46676 164898 46704 272478
rect 46768 260166 46796 388690
rect 46756 260160 46808 260166
rect 46756 260102 46808 260108
rect 46860 258777 46888 413238
rect 48056 389162 48084 549238
rect 48148 443698 48176 563654
rect 50896 560312 50948 560318
rect 50896 560254 50948 560260
rect 49516 533452 49568 533458
rect 49516 533394 49568 533400
rect 48136 443692 48188 443698
rect 48136 443634 48188 443640
rect 48134 436112 48190 436121
rect 48134 436047 48190 436056
rect 48044 389156 48096 389162
rect 48044 389098 48096 389104
rect 48056 388754 48084 389098
rect 48044 388748 48096 388754
rect 48044 388690 48096 388696
rect 48042 385656 48098 385665
rect 48042 385591 48098 385600
rect 47952 278724 48004 278730
rect 47952 278666 48004 278672
rect 47964 278050 47992 278666
rect 47952 278044 48004 278050
rect 47952 277986 48004 277992
rect 46846 258768 46902 258777
rect 46846 258703 46902 258712
rect 47964 221474 47992 277986
rect 48056 237386 48084 385591
rect 48148 278730 48176 436047
rect 49528 396030 49556 533394
rect 50908 511290 50936 560254
rect 50896 511284 50948 511290
rect 50896 511226 50948 511232
rect 50908 438190 50936 511226
rect 50896 438184 50948 438190
rect 50896 438126 50948 438132
rect 50896 425740 50948 425746
rect 50896 425682 50948 425688
rect 49608 422952 49660 422958
rect 49608 422894 49660 422900
rect 49516 396024 49568 396030
rect 49516 395966 49568 395972
rect 49528 395282 49556 395966
rect 48228 395276 48280 395282
rect 48228 395218 48280 395224
rect 49516 395276 49568 395282
rect 49516 395218 49568 395224
rect 48136 278724 48188 278730
rect 48136 278666 48188 278672
rect 48134 254144 48190 254153
rect 48134 254079 48190 254088
rect 48044 237380 48096 237386
rect 48044 237322 48096 237328
rect 48044 229764 48096 229770
rect 48044 229706 48096 229712
rect 47952 221468 48004 221474
rect 47952 221410 48004 221416
rect 46848 203584 46900 203590
rect 46848 203526 46900 203532
rect 46664 164892 46716 164898
rect 46664 164834 46716 164840
rect 46676 161474 46704 164834
rect 46676 161446 46796 161474
rect 46768 122806 46796 161446
rect 46756 122800 46808 122806
rect 46756 122742 46808 122748
rect 46860 90370 46888 203526
rect 48056 92546 48084 229706
rect 48148 105602 48176 254079
rect 48240 245002 48268 395218
rect 49516 393984 49568 393990
rect 49516 393926 49568 393932
rect 49528 393378 49556 393926
rect 49516 393372 49568 393378
rect 49516 393314 49568 393320
rect 48228 244996 48280 245002
rect 48228 244938 48280 244944
rect 49528 242962 49556 393314
rect 49620 266529 49648 422894
rect 50804 369164 50856 369170
rect 50804 369106 50856 369112
rect 49606 266520 49662 266529
rect 49606 266455 49662 266464
rect 49516 242956 49568 242962
rect 49516 242898 49568 242904
rect 49514 217288 49570 217297
rect 49514 217223 49570 217232
rect 48226 206272 48282 206281
rect 48226 206207 48282 206216
rect 48136 105596 48188 105602
rect 48136 105538 48188 105544
rect 48044 92540 48096 92546
rect 48044 92482 48096 92488
rect 46848 90364 46900 90370
rect 46848 90306 46900 90312
rect 46848 39364 46900 39370
rect 46848 39306 46900 39312
rect 46860 6914 46888 39306
rect 48240 6914 48268 206207
rect 46676 6886 46888 6914
rect 47872 6886 48268 6914
rect 46676 480 46704 6886
rect 47872 480 47900 6886
rect 49528 3534 49556 217223
rect 49620 216646 49648 266455
rect 50528 265668 50580 265674
rect 50528 265610 50580 265616
rect 50540 265033 50568 265610
rect 50526 265024 50582 265033
rect 50526 264959 50582 264968
rect 50620 258732 50672 258738
rect 50620 258674 50672 258680
rect 49608 216640 49660 216646
rect 49608 216582 49660 216588
rect 50632 106962 50660 258674
rect 50816 237454 50844 369106
rect 50908 268433 50936 425682
rect 51000 422278 51028 580994
rect 52276 565888 52328 565894
rect 52276 565830 52328 565836
rect 50988 422272 51040 422278
rect 50988 422214 51040 422220
rect 51000 421598 51028 422214
rect 50988 421592 51040 421598
rect 50988 421534 51040 421540
rect 52288 411262 52316 565830
rect 52380 446418 52408 582354
rect 53748 557592 53800 557598
rect 53748 557534 53800 557540
rect 53472 546508 53524 546514
rect 53472 546450 53524 546456
rect 52368 446412 52420 446418
rect 52368 446354 52420 446360
rect 52368 429276 52420 429282
rect 52368 429218 52420 429224
rect 52276 411256 52328 411262
rect 52276 411198 52328 411204
rect 52288 409970 52316 411198
rect 50988 409964 51040 409970
rect 50988 409906 51040 409912
rect 52276 409964 52328 409970
rect 52276 409906 52328 409912
rect 50894 268424 50950 268433
rect 50894 268359 50950 268368
rect 50894 265024 50950 265033
rect 50894 264959 50950 264968
rect 50804 237448 50856 237454
rect 50804 237390 50856 237396
rect 50908 231849 50936 264959
rect 51000 257378 51028 409906
rect 51724 409896 51776 409902
rect 51724 409838 51776 409844
rect 51736 389201 51764 409838
rect 51722 389192 51778 389201
rect 51722 389127 51778 389136
rect 52276 387116 52328 387122
rect 52276 387058 52328 387064
rect 52182 384296 52238 384305
rect 52182 384231 52238 384240
rect 52090 285968 52146 285977
rect 52090 285903 52146 285912
rect 50988 257372 51040 257378
rect 50988 257314 51040 257320
rect 51080 256012 51132 256018
rect 51080 255954 51132 255960
rect 51092 255338 51120 255954
rect 51080 255332 51132 255338
rect 51080 255274 51132 255280
rect 52000 255332 52052 255338
rect 52000 255274 52052 255280
rect 50894 231840 50950 231849
rect 50894 231775 50950 231784
rect 50710 153096 50766 153105
rect 50710 153031 50766 153040
rect 50724 151881 50752 153031
rect 50710 151872 50766 151881
rect 50710 151807 50766 151816
rect 50908 151814 50936 231775
rect 52012 223553 52040 255274
rect 51998 223544 52054 223553
rect 51998 223479 52054 223488
rect 52104 175409 52132 285903
rect 52196 241466 52224 384231
rect 52184 241460 52236 241466
rect 52184 241402 52236 241408
rect 52288 239873 52316 387058
rect 52380 272542 52408 429218
rect 53484 391513 53512 546450
rect 53760 449206 53788 557534
rect 54944 544400 54996 544406
rect 54944 544342 54996 544348
rect 53748 449200 53800 449206
rect 53748 449142 53800 449148
rect 54956 440978 54984 544342
rect 55036 518220 55088 518226
rect 55036 518162 55088 518168
rect 54944 440972 54996 440978
rect 54944 440914 54996 440920
rect 54942 433528 54998 433537
rect 54942 433463 54998 433472
rect 53748 426488 53800 426494
rect 53748 426430 53800 426436
rect 53564 415472 53616 415478
rect 53564 415414 53616 415420
rect 53470 391504 53526 391513
rect 53470 391439 53526 391448
rect 53576 322930 53604 415414
rect 53656 392624 53708 392630
rect 53656 392566 53708 392572
rect 53564 322924 53616 322930
rect 53564 322866 53616 322872
rect 53104 320204 53156 320210
rect 53104 320146 53156 320152
rect 52368 272536 52420 272542
rect 52368 272478 52420 272484
rect 53116 263566 53144 320146
rect 53472 283620 53524 283626
rect 53472 283562 53524 283568
rect 53104 263560 53156 263566
rect 53104 263502 53156 263508
rect 52274 239864 52330 239873
rect 52274 239799 52330 239808
rect 52366 238096 52422 238105
rect 52366 238031 52422 238040
rect 52380 237454 52408 238031
rect 52368 237448 52420 237454
rect 52368 237390 52420 237396
rect 52274 223544 52330 223553
rect 52274 223479 52330 223488
rect 52288 222329 52316 223479
rect 52274 222320 52330 222329
rect 52274 222255 52330 222264
rect 52090 175400 52146 175409
rect 52090 175335 52146 175344
rect 52104 171134 52132 175335
rect 52104 171106 52224 171134
rect 50724 132462 50752 151807
rect 50816 151786 50936 151814
rect 50816 150793 50844 151786
rect 50802 150784 50858 150793
rect 50802 150719 50858 150728
rect 50712 132456 50764 132462
rect 50712 132398 50764 132404
rect 50816 115938 50844 150719
rect 50894 148336 50950 148345
rect 50894 148271 50950 148280
rect 50804 115932 50856 115938
rect 50804 115874 50856 115880
rect 50620 106956 50672 106962
rect 50620 106898 50672 106904
rect 50908 3534 50936 148271
rect 52196 138718 52224 171106
rect 52184 138712 52236 138718
rect 52184 138654 52236 138660
rect 52288 107642 52316 222255
rect 52276 107636 52328 107642
rect 52276 107578 52328 107584
rect 52380 90953 52408 237390
rect 53484 167686 53512 283562
rect 53564 268388 53616 268394
rect 53564 268330 53616 268336
rect 53576 267782 53604 268330
rect 53564 267776 53616 267782
rect 53564 267718 53616 267724
rect 53472 167680 53524 167686
rect 53472 167622 53524 167628
rect 53484 133210 53512 167622
rect 53576 149161 53604 267718
rect 53668 244934 53696 392566
rect 53760 271182 53788 426430
rect 53840 409828 53892 409834
rect 53840 409770 53892 409776
rect 53852 409154 53880 409770
rect 53840 409148 53892 409154
rect 53840 409090 53892 409096
rect 54852 385688 54904 385694
rect 54852 385630 54904 385636
rect 53748 271176 53800 271182
rect 53748 271118 53800 271124
rect 53746 251288 53802 251297
rect 53746 251223 53802 251232
rect 53656 244928 53708 244934
rect 53656 244870 53708 244876
rect 53654 149696 53710 149705
rect 53654 149631 53710 149640
rect 53562 149152 53618 149161
rect 53562 149087 53618 149096
rect 53472 133204 53524 133210
rect 53472 133146 53524 133152
rect 53576 118590 53604 149087
rect 53564 118584 53616 118590
rect 53564 118526 53616 118532
rect 52366 90944 52422 90953
rect 52366 90879 52422 90888
rect 53668 16574 53696 149631
rect 53760 100774 53788 251223
rect 54864 242214 54892 385630
rect 54956 289785 54984 433463
rect 55048 409834 55076 518162
rect 55036 409828 55088 409834
rect 55036 409770 55088 409776
rect 55036 398880 55088 398886
rect 55036 398822 55088 398828
rect 54942 289776 54998 289785
rect 54942 289711 54998 289720
rect 54944 275324 54996 275330
rect 54944 275266 54996 275272
rect 54852 242208 54904 242214
rect 54852 242150 54904 242156
rect 54956 157457 54984 275266
rect 55048 248470 55076 398822
rect 55140 385014 55168 585142
rect 56508 572008 56560 572014
rect 56508 571950 56560 571956
rect 56416 414044 56468 414050
rect 56416 413986 56468 413992
rect 55128 385008 55180 385014
rect 55128 384950 55180 384956
rect 55126 289776 55182 289785
rect 55126 289711 55182 289720
rect 55140 277370 55168 289711
rect 55128 277364 55180 277370
rect 55128 277306 55180 277312
rect 56324 269816 56376 269822
rect 56324 269758 56376 269764
rect 55128 260228 55180 260234
rect 55128 260170 55180 260176
rect 55036 248464 55088 248470
rect 55036 248406 55088 248412
rect 55036 242956 55088 242962
rect 55036 242898 55088 242904
rect 55048 211177 55076 242898
rect 55034 211168 55090 211177
rect 55034 211103 55090 211112
rect 54942 157448 54998 157457
rect 54942 157383 54998 157392
rect 54482 136096 54538 136105
rect 54482 136031 54538 136040
rect 53840 119400 53892 119406
rect 53840 119342 53892 119348
rect 53852 113830 53880 119342
rect 53840 113824 53892 113830
rect 53840 113766 53892 113772
rect 53748 100768 53800 100774
rect 53748 100710 53800 100716
rect 54496 33114 54524 136031
rect 54956 126954 54984 157383
rect 54944 126948 54996 126954
rect 54944 126890 54996 126896
rect 55048 95849 55076 211103
rect 55140 109750 55168 260170
rect 55864 260160 55916 260166
rect 55864 260102 55916 260108
rect 55876 237318 55904 260102
rect 55864 237312 55916 237318
rect 55864 237254 55916 237260
rect 56336 156058 56364 269758
rect 56428 261526 56456 413986
rect 56520 407114 56548 571950
rect 57808 564398 57836 702510
rect 59266 581224 59322 581233
rect 59266 581159 59322 581168
rect 57888 580304 57940 580310
rect 57888 580246 57940 580252
rect 57900 579698 57928 580246
rect 57888 579692 57940 579698
rect 57888 579634 57940 579640
rect 57796 564392 57848 564398
rect 57796 564334 57848 564340
rect 57808 563718 57836 564334
rect 57796 563712 57848 563718
rect 57796 563654 57848 563660
rect 57796 553444 57848 553450
rect 57796 553386 57848 553392
rect 57704 436212 57756 436218
rect 57704 436154 57756 436160
rect 56508 407108 56560 407114
rect 56508 407050 56560 407056
rect 57612 400240 57664 400246
rect 57612 400182 57664 400188
rect 56508 392012 56560 392018
rect 56508 391954 56560 391960
rect 56520 299538 56548 391954
rect 57624 331294 57652 400182
rect 57612 331288 57664 331294
rect 57612 331230 57664 331236
rect 56508 299532 56560 299538
rect 56508 299474 56560 299480
rect 56416 261520 56468 261526
rect 56416 261462 56468 261468
rect 56520 246362 56548 299474
rect 57610 290456 57666 290465
rect 57610 290391 57666 290400
rect 57520 260160 57572 260166
rect 57520 260102 57572 260108
rect 56508 246356 56560 246362
rect 56508 246298 56560 246304
rect 56508 235272 56560 235278
rect 56508 235214 56560 235220
rect 56324 156052 56376 156058
rect 56324 155994 56376 156000
rect 56336 151814 56364 155994
rect 56336 151786 56456 151814
rect 56428 120086 56456 151786
rect 56416 120080 56468 120086
rect 56416 120022 56468 120028
rect 55128 109744 55180 109750
rect 55128 109686 55180 109692
rect 55034 95840 55090 95849
rect 55034 95775 55090 95784
rect 56520 89729 56548 235214
rect 57532 111110 57560 260102
rect 57624 258738 57652 290391
rect 57716 283626 57744 436154
rect 57808 417450 57836 553386
rect 57796 417444 57848 417450
rect 57796 417386 57848 417392
rect 57796 407108 57848 407114
rect 57796 407050 57848 407056
rect 57808 405754 57836 407050
rect 57796 405748 57848 405754
rect 57796 405690 57848 405696
rect 57704 283620 57756 283626
rect 57704 283562 57756 283568
rect 57612 258732 57664 258738
rect 57612 258674 57664 258680
rect 57808 254590 57836 405690
rect 57900 387802 57928 579634
rect 59176 558952 59228 558958
rect 59176 558894 59228 558900
rect 59084 431996 59136 432002
rect 59084 431938 59136 431944
rect 58900 400308 58952 400314
rect 58900 400250 58952 400256
rect 57888 387796 57940 387802
rect 57888 387738 57940 387744
rect 57888 331288 57940 331294
rect 57888 331230 57940 331236
rect 57796 254584 57848 254590
rect 57796 254526 57848 254532
rect 57900 251122 57928 331230
rect 58912 251190 58940 400250
rect 58992 292596 59044 292602
rect 58992 292538 59044 292544
rect 58900 251184 58952 251190
rect 58900 251126 58952 251132
rect 57888 251116 57940 251122
rect 57888 251058 57940 251064
rect 57900 249830 57928 251058
rect 57888 249824 57940 249830
rect 57888 249766 57940 249772
rect 57796 248464 57848 248470
rect 57796 248406 57848 248412
rect 57702 244488 57758 244497
rect 57702 244423 57758 244432
rect 57716 212673 57744 244423
rect 57702 212664 57758 212673
rect 57702 212599 57758 212608
rect 57612 178152 57664 178158
rect 57612 178094 57664 178100
rect 57624 125594 57652 178094
rect 57612 125588 57664 125594
rect 57612 125530 57664 125536
rect 57520 111104 57572 111110
rect 57520 111046 57572 111052
rect 57716 97306 57744 212599
rect 57808 100026 57836 248406
rect 57888 244996 57940 245002
rect 57888 244938 57940 244944
rect 57900 244497 57928 244938
rect 57886 244488 57942 244497
rect 57886 244423 57942 244432
rect 59004 233170 59032 292538
rect 59096 277681 59124 431938
rect 59188 396846 59216 558894
rect 59280 413302 59308 581159
rect 60648 567248 60700 567254
rect 60648 567190 60700 567196
rect 60004 532024 60056 532030
rect 60004 531966 60056 531972
rect 60016 415478 60044 531966
rect 60660 453354 60688 567190
rect 61948 544406 61976 702850
rect 66076 702500 66128 702506
rect 66076 702442 66128 702448
rect 62028 582480 62080 582486
rect 62028 582422 62080 582428
rect 61936 544400 61988 544406
rect 61936 544342 61988 544348
rect 61292 539640 61344 539646
rect 61292 539582 61344 539588
rect 61304 536722 61332 539582
rect 61844 537532 61896 537538
rect 61844 537474 61896 537480
rect 61292 536716 61344 536722
rect 61292 536658 61344 536664
rect 60648 453348 60700 453354
rect 60648 453290 60700 453296
rect 61752 433356 61804 433362
rect 61752 433298 61804 433304
rect 60556 430636 60608 430642
rect 60556 430578 60608 430584
rect 60004 415472 60056 415478
rect 60004 415414 60056 415420
rect 60016 414798 60044 415414
rect 60004 414792 60056 414798
rect 60004 414734 60056 414740
rect 59268 413296 59320 413302
rect 59268 413238 59320 413244
rect 59268 411324 59320 411330
rect 59268 411266 59320 411272
rect 59176 396840 59228 396846
rect 59176 396782 59228 396788
rect 59176 293344 59228 293350
rect 59176 293286 59228 293292
rect 59188 292602 59216 293286
rect 59176 292596 59228 292602
rect 59176 292538 59228 292544
rect 59082 277672 59138 277681
rect 59082 277607 59138 277616
rect 59280 259418 59308 411266
rect 59360 322924 59412 322930
rect 59360 322866 59412 322872
rect 59372 260234 59400 322866
rect 60464 287088 60516 287094
rect 60464 287030 60516 287036
rect 60370 271960 60426 271969
rect 60370 271895 60426 271904
rect 59360 260228 59412 260234
rect 59360 260170 59412 260176
rect 59268 259412 59320 259418
rect 59268 259354 59320 259360
rect 59084 257372 59136 257378
rect 59084 257314 59136 257320
rect 58992 233164 59044 233170
rect 58992 233106 59044 233112
rect 59096 226302 59124 257314
rect 59176 254584 59228 254590
rect 59176 254526 59228 254532
rect 59188 228993 59216 254526
rect 59268 249756 59320 249762
rect 59268 249698 59320 249704
rect 59174 228984 59230 228993
rect 59174 228919 59230 228928
rect 59084 226296 59136 226302
rect 59084 226238 59136 226244
rect 59096 143585 59124 226238
rect 59082 143576 59138 143585
rect 59082 143511 59138 143520
rect 59096 109002 59124 143511
rect 59084 108996 59136 109002
rect 59084 108938 59136 108944
rect 59084 106956 59136 106962
rect 59084 106898 59136 106904
rect 59096 106350 59124 106898
rect 59084 106344 59136 106350
rect 59084 106286 59136 106292
rect 57888 100768 57940 100774
rect 57888 100710 57940 100716
rect 57796 100020 57848 100026
rect 57796 99962 57848 99968
rect 57704 97300 57756 97306
rect 57704 97242 57756 97248
rect 57244 96688 57296 96694
rect 57244 96630 57296 96636
rect 56506 89720 56562 89729
rect 56506 89655 56562 89664
rect 57256 86601 57284 96630
rect 57242 86592 57298 86601
rect 57242 86527 57298 86536
rect 57900 73137 57928 100710
rect 59096 74526 59124 106286
rect 59188 104854 59216 228919
rect 59176 104848 59228 104854
rect 59176 104790 59228 104796
rect 59280 101318 59308 249698
rect 60384 154630 60412 271895
rect 60476 229838 60504 287030
rect 60568 273329 60596 430578
rect 60648 427848 60700 427854
rect 60648 427790 60700 427796
rect 60554 273320 60610 273329
rect 60554 273255 60610 273264
rect 60660 270609 60688 427790
rect 60740 423496 60792 423502
rect 60740 423438 60792 423444
rect 60752 422958 60780 423438
rect 60740 422952 60792 422958
rect 60740 422894 60792 422900
rect 61384 325712 61436 325718
rect 61384 325654 61436 325660
rect 60646 270600 60702 270609
rect 60646 270535 60702 270544
rect 60660 258074 60688 270535
rect 60568 258046 60688 258074
rect 60464 229832 60516 229838
rect 60464 229774 60516 229780
rect 60568 160857 60596 258046
rect 61014 251288 61070 251297
rect 61014 251223 61070 251232
rect 61028 250782 61056 251223
rect 61396 250782 61424 325654
rect 61764 284345 61792 433298
rect 61856 423502 61884 537474
rect 61934 432848 61990 432857
rect 61934 432783 61990 432792
rect 61844 423496 61896 423502
rect 61844 423438 61896 423444
rect 61844 419552 61896 419558
rect 61844 419494 61896 419500
rect 61750 284336 61806 284345
rect 61750 284271 61806 284280
rect 61658 283248 61714 283257
rect 61658 283183 61714 283192
rect 61016 250776 61068 250782
rect 61016 250718 61068 250724
rect 61384 250776 61436 250782
rect 61384 250718 61436 250724
rect 61672 233918 61700 283183
rect 61750 273320 61806 273329
rect 61750 273255 61806 273264
rect 61660 233912 61712 233918
rect 61660 233854 61712 233860
rect 61764 190454 61792 273255
rect 61856 265198 61884 419494
rect 61948 276214 61976 432783
rect 62040 389298 62068 582422
rect 64788 579692 64840 579698
rect 64788 579634 64840 579640
rect 63406 578912 63462 578921
rect 63406 578847 63462 578856
rect 63316 554804 63368 554810
rect 63316 554746 63368 554752
rect 63328 490618 63356 554746
rect 63316 490612 63368 490618
rect 63316 490554 63368 490560
rect 63314 434752 63370 434761
rect 63314 434687 63370 434696
rect 63224 404388 63276 404394
rect 63224 404330 63276 404336
rect 62028 389292 62080 389298
rect 62028 389234 62080 389240
rect 63132 284436 63184 284442
rect 63132 284378 63184 284384
rect 61936 276208 61988 276214
rect 61936 276150 61988 276156
rect 61948 275330 61976 276150
rect 61936 275324 61988 275330
rect 61936 275266 61988 275272
rect 63038 268424 63094 268433
rect 63038 268359 63094 268368
rect 61844 265192 61896 265198
rect 61844 265134 61896 265140
rect 62026 263664 62082 263673
rect 62026 263599 62082 263608
rect 61844 251184 61896 251190
rect 61844 251126 61896 251132
rect 61856 248577 61884 251126
rect 61842 248568 61898 248577
rect 61842 248503 61898 248512
rect 61856 229022 61884 248503
rect 61936 248396 61988 248402
rect 61936 248338 61988 248344
rect 61948 248305 61976 248338
rect 61934 248296 61990 248305
rect 61934 248231 61990 248240
rect 61844 229016 61896 229022
rect 61844 228958 61896 228964
rect 61934 216744 61990 216753
rect 61934 216679 61990 216688
rect 61764 190426 61884 190454
rect 61856 169833 61884 190426
rect 61842 169824 61898 169833
rect 61842 169759 61898 169768
rect 60554 160848 60610 160857
rect 60554 160783 60610 160792
rect 60372 154624 60424 154630
rect 60372 154566 60424 154572
rect 60384 151814 60412 154566
rect 60384 151786 60504 151814
rect 60476 121446 60504 151786
rect 60464 121440 60516 121446
rect 60464 121382 60516 121388
rect 60568 121378 60596 160783
rect 60740 160744 60792 160750
rect 60740 160686 60792 160692
rect 60752 160138 60780 160686
rect 60740 160132 60792 160138
rect 60740 160074 60792 160080
rect 61752 160132 61804 160138
rect 61752 160074 61804 160080
rect 60646 155272 60702 155281
rect 60646 155207 60702 155216
rect 60556 121372 60608 121378
rect 60556 121314 60608 121320
rect 59268 101312 59320 101318
rect 59268 101254 59320 101260
rect 59084 74520 59136 74526
rect 59084 74462 59136 74468
rect 59096 73234 59124 74462
rect 58624 73228 58676 73234
rect 58624 73170 58676 73176
rect 59084 73228 59136 73234
rect 59084 73170 59136 73176
rect 57886 73128 57942 73137
rect 57886 73063 57942 73072
rect 57900 71913 57928 73063
rect 57242 71904 57298 71913
rect 57242 71839 57298 71848
rect 57886 71904 57942 71913
rect 57886 71839 57942 71848
rect 55128 50380 55180 50386
rect 55128 50322 55180 50328
rect 54484 33108 54536 33114
rect 54484 33050 54536 33056
rect 53748 29640 53800 29646
rect 53748 29582 53800 29588
rect 53576 16546 53696 16574
rect 52552 3596 52604 3602
rect 52552 3538 52604 3544
rect 48964 3528 49016 3534
rect 48964 3470 49016 3476
rect 49516 3528 49568 3534
rect 49516 3470 49568 3476
rect 50160 3528 50212 3534
rect 50160 3470 50212 3476
rect 50896 3528 50948 3534
rect 50896 3470 50948 3476
rect 48976 480 49004 3470
rect 50172 480 50200 3470
rect 51356 2100 51408 2106
rect 51356 2042 51408 2048
rect 51368 480 51396 2042
rect 52564 480 52592 3538
rect 53576 3482 53604 16546
rect 53760 6914 53788 29582
rect 55140 6914 55168 50322
rect 57256 45558 57284 71839
rect 57888 58676 57940 58682
rect 57888 58618 57940 58624
rect 57244 45552 57296 45558
rect 57244 45494 57296 45500
rect 53668 6886 53788 6914
rect 54956 6886 55168 6914
rect 53668 3602 53696 6886
rect 53656 3596 53708 3602
rect 53656 3538 53708 3544
rect 53576 3454 53788 3482
rect 53760 480 53788 3454
rect 54956 480 54984 6886
rect 56048 6180 56100 6186
rect 56048 6122 56100 6128
rect 56060 480 56088 6122
rect 57900 3534 57928 58618
rect 58636 6866 58664 73170
rect 59268 44872 59320 44878
rect 59268 44814 59320 44820
rect 58624 6860 58676 6866
rect 58624 6802 58676 6808
rect 59280 3534 59308 44814
rect 60660 3534 60688 155207
rect 61764 128314 61792 160074
rect 61752 128308 61804 128314
rect 61752 128250 61804 128256
rect 61856 124166 61884 169759
rect 61844 124160 61896 124166
rect 61844 124102 61896 124108
rect 60740 109744 60792 109750
rect 60740 109686 60792 109692
rect 60752 109070 60780 109686
rect 60740 109064 60792 109070
rect 60740 109006 60792 109012
rect 61384 109064 61436 109070
rect 61384 109006 61436 109012
rect 61396 85542 61424 109006
rect 61844 101312 61896 101318
rect 61844 101254 61896 101260
rect 61384 85536 61436 85542
rect 61384 85478 61436 85484
rect 61856 77178 61884 101254
rect 61948 99346 61976 216679
rect 62040 139505 62068 263599
rect 62120 242208 62172 242214
rect 62120 242150 62172 242156
rect 62132 241641 62160 242150
rect 62118 241632 62174 241641
rect 62118 241567 62174 241576
rect 63052 224262 63080 268359
rect 63144 238134 63172 284378
rect 63236 253910 63264 404330
rect 63328 282878 63356 434687
rect 63420 433362 63448 578847
rect 64696 571396 64748 571402
rect 64696 571338 64748 571344
rect 64604 457496 64656 457502
rect 64604 457438 64656 457444
rect 63408 433356 63460 433362
rect 63408 433298 63460 433304
rect 63406 420880 63462 420889
rect 63406 420815 63462 420824
rect 63316 282872 63368 282878
rect 63316 282814 63368 282820
rect 63420 267734 63448 420815
rect 64144 416900 64196 416906
rect 64144 416842 64196 416848
rect 64156 320210 64184 416842
rect 64616 411330 64644 457438
rect 64708 454714 64736 571338
rect 64800 458862 64828 579634
rect 65982 568848 66038 568857
rect 65982 568783 66038 568792
rect 65996 529242 66024 568783
rect 66088 546009 66116 702442
rect 67548 589960 67600 589966
rect 67548 589902 67600 589908
rect 66810 580000 66866 580009
rect 66810 579935 66866 579944
rect 66824 579698 66852 579935
rect 66812 579692 66864 579698
rect 66812 579634 66864 579640
rect 66810 578640 66866 578649
rect 66810 578575 66866 578584
rect 66534 575920 66590 575929
rect 66534 575855 66590 575864
rect 66548 575550 66576 575855
rect 66536 575544 66588 575550
rect 66536 575486 66588 575492
rect 66442 573200 66498 573209
rect 66442 573135 66498 573144
rect 66456 572014 66484 573135
rect 66444 572008 66496 572014
rect 66444 571950 66496 571956
rect 66718 571840 66774 571849
rect 66718 571775 66774 571784
rect 66732 571402 66760 571775
rect 66720 571396 66772 571402
rect 66720 571338 66772 571344
rect 66718 564768 66774 564777
rect 66718 564703 66774 564712
rect 66732 564466 66760 564703
rect 66720 564460 66772 564466
rect 66720 564402 66772 564408
rect 66444 564392 66496 564398
rect 66444 564334 66496 564340
rect 66456 564233 66484 564334
rect 66442 564224 66498 564233
rect 66442 564159 66498 564168
rect 66166 562048 66222 562057
rect 66166 561983 66222 561992
rect 66074 546000 66130 546009
rect 66074 545935 66130 545944
rect 65984 529236 66036 529242
rect 65984 529178 66036 529184
rect 66088 482322 66116 545935
rect 66076 482316 66128 482322
rect 66076 482258 66128 482264
rect 65984 466472 66036 466478
rect 65984 466414 66036 466420
rect 64788 458856 64840 458862
rect 64788 458798 64840 458804
rect 64696 454708 64748 454714
rect 64696 454650 64748 454656
rect 65890 449984 65946 449993
rect 65890 449919 65946 449928
rect 64788 418192 64840 418198
rect 64788 418134 64840 418140
rect 64604 411324 64656 411330
rect 64604 411266 64656 411272
rect 64604 320884 64656 320890
rect 64604 320826 64656 320832
rect 63500 320204 63552 320210
rect 63500 320146 63552 320152
rect 64144 320204 64196 320210
rect 64144 320146 64196 320152
rect 63512 319462 63540 320146
rect 63500 319456 63552 319462
rect 63500 319398 63552 319404
rect 64512 285728 64564 285734
rect 64512 285670 64564 285676
rect 63328 267706 63448 267734
rect 63328 266422 63356 267706
rect 63316 266416 63368 266422
rect 63316 266358 63368 266364
rect 63224 253904 63276 253910
rect 63224 253846 63276 253852
rect 63132 238128 63184 238134
rect 63132 238070 63184 238076
rect 63040 224256 63092 224262
rect 63040 224198 63092 224204
rect 63130 144936 63186 144945
rect 63130 144871 63186 144880
rect 62026 139496 62082 139505
rect 62026 139431 62082 139440
rect 62040 114510 62068 139431
rect 63144 117230 63172 144871
rect 63328 142225 63356 266358
rect 63406 241632 63462 241641
rect 63406 241567 63462 241576
rect 63314 142216 63370 142225
rect 63314 142154 63370 142160
rect 63236 142151 63370 142154
rect 63236 142126 63356 142151
rect 63236 117298 63264 142126
rect 63224 117292 63276 117298
rect 63224 117234 63276 117240
rect 63132 117224 63184 117230
rect 63132 117166 63184 117172
rect 62028 114504 62080 114510
rect 62028 114446 62080 114452
rect 62028 113824 62080 113830
rect 62028 113766 62080 113772
rect 61936 99340 61988 99346
rect 61936 99282 61988 99288
rect 62040 86902 62068 113766
rect 63316 107704 63368 107710
rect 63316 107646 63368 107652
rect 62028 86896 62080 86902
rect 62028 86838 62080 86844
rect 63328 81394 63356 107646
rect 63420 93838 63448 241567
rect 64524 240786 64552 285670
rect 64512 240780 64564 240786
rect 64512 240722 64564 240728
rect 64616 240009 64644 320826
rect 64694 284336 64750 284345
rect 64694 284271 64750 284280
rect 64708 276010 64736 284271
rect 64696 276004 64748 276010
rect 64696 275946 64748 275952
rect 64694 274816 64750 274825
rect 64694 274751 64750 274760
rect 64602 240000 64658 240009
rect 64602 239935 64658 239944
rect 64708 150550 64736 274751
rect 64800 263673 64828 418134
rect 65904 386374 65932 449919
rect 65996 425746 66024 466414
rect 66074 429312 66130 429321
rect 66074 429247 66130 429256
rect 65984 425740 66036 425746
rect 65984 425682 66036 425688
rect 65982 403744 66038 403753
rect 65982 403679 66038 403688
rect 65892 386368 65944 386374
rect 65892 386310 65944 386316
rect 65892 305652 65944 305658
rect 65892 305594 65944 305600
rect 65904 279478 65932 305594
rect 65892 279472 65944 279478
rect 65892 279414 65944 279420
rect 65708 265192 65760 265198
rect 65706 265160 65708 265169
rect 65760 265160 65762 265169
rect 65706 265095 65762 265104
rect 64786 263664 64842 263673
rect 64786 263599 64842 263608
rect 65892 262880 65944 262886
rect 65892 262822 65944 262828
rect 64788 251388 64840 251394
rect 64788 251330 64840 251336
rect 64696 150544 64748 150550
rect 64696 150486 64748 150492
rect 64512 140072 64564 140078
rect 64512 140014 64564 140020
rect 63408 93832 63460 93838
rect 63408 93774 63460 93780
rect 64524 91050 64552 140014
rect 64602 138816 64658 138825
rect 64602 138751 64658 138760
rect 64616 92449 64644 138751
rect 64708 124982 64736 150486
rect 64696 124976 64748 124982
rect 64696 124918 64748 124924
rect 64800 102406 64828 251330
rect 65904 233238 65932 262822
rect 65996 251394 66024 403679
rect 66088 271969 66116 429247
rect 66180 394641 66208 561983
rect 66534 549536 66590 549545
rect 66534 549471 66590 549480
rect 66548 549302 66576 549471
rect 66536 549296 66588 549302
rect 66536 549238 66588 549244
rect 66718 544640 66774 544649
rect 66718 544575 66774 544584
rect 66732 544406 66760 544575
rect 66720 544400 66772 544406
rect 66720 544342 66772 544348
rect 66258 433392 66314 433401
rect 66258 433327 66260 433336
rect 66312 433327 66314 433336
rect 66260 433298 66312 433304
rect 66442 432576 66498 432585
rect 66442 432511 66498 432520
rect 66456 432002 66484 432511
rect 66444 431996 66496 432002
rect 66444 431938 66496 431944
rect 66718 431488 66774 431497
rect 66718 431423 66774 431432
rect 66732 430642 66760 431423
rect 66720 430636 66772 430642
rect 66720 430578 66772 430584
rect 66718 430400 66774 430409
rect 66718 430335 66774 430344
rect 66732 429282 66760 430335
rect 66720 429276 66772 429282
rect 66720 429218 66772 429224
rect 66718 428224 66774 428233
rect 66718 428159 66774 428168
rect 66732 427854 66760 428159
rect 66720 427848 66772 427854
rect 66720 427790 66772 427796
rect 66718 427408 66774 427417
rect 66718 427343 66774 427352
rect 66732 426494 66760 427343
rect 66720 426488 66772 426494
rect 66720 426430 66772 426436
rect 66536 425740 66588 425746
rect 66536 425682 66588 425688
rect 66548 425241 66576 425682
rect 66534 425232 66590 425241
rect 66534 425167 66590 425176
rect 66718 424144 66774 424153
rect 66718 424079 66774 424088
rect 66732 423706 66760 424079
rect 66720 423700 66772 423706
rect 66720 423642 66772 423648
rect 66720 423496 66772 423502
rect 66720 423438 66772 423444
rect 66732 423337 66760 423438
rect 66718 423328 66774 423337
rect 66718 423263 66774 423272
rect 66626 418976 66682 418985
rect 66626 418911 66682 418920
rect 66640 418198 66668 418911
rect 66628 418192 66680 418198
rect 66628 418134 66680 418140
rect 66628 417444 66680 417450
rect 66628 417386 66680 417392
rect 66640 415993 66668 417386
rect 66626 415984 66682 415993
rect 66626 415919 66682 415928
rect 66718 414896 66774 414905
rect 66718 414831 66774 414840
rect 66732 414050 66760 414831
rect 66720 414044 66772 414050
rect 66720 413986 66772 413992
rect 66718 411904 66774 411913
rect 66718 411839 66774 411848
rect 66732 411330 66760 411839
rect 66720 411324 66772 411330
rect 66720 411266 66772 411272
rect 66260 409828 66312 409834
rect 66260 409770 66312 409776
rect 66272 408921 66300 409770
rect 66258 408912 66314 408921
rect 66258 408847 66314 408856
rect 66442 406736 66498 406745
rect 66442 406671 66498 406680
rect 66456 405754 66484 406671
rect 66444 405748 66496 405754
rect 66444 405690 66496 405696
rect 66824 402974 66852 578575
rect 67454 577280 67510 577289
rect 67454 577215 67510 577224
rect 66902 570208 66958 570217
rect 66902 570143 66958 570152
rect 66916 420186 66944 570143
rect 66994 567488 67050 567497
rect 66994 567423 67050 567432
rect 67008 567254 67036 567423
rect 66996 567248 67048 567254
rect 66996 567190 67048 567196
rect 66994 560688 67050 560697
rect 66994 560623 67050 560632
rect 67008 560318 67036 560623
rect 66996 560312 67048 560318
rect 66996 560254 67048 560260
rect 66994 559328 67050 559337
rect 66994 559263 67050 559272
rect 67008 558958 67036 559263
rect 66996 558952 67048 558958
rect 66996 558894 67048 558900
rect 66994 557968 67050 557977
rect 66994 557903 67050 557912
rect 67008 557598 67036 557903
rect 66996 557592 67048 557598
rect 66996 557534 67048 557540
rect 66994 555248 67050 555257
rect 66994 555183 67050 555192
rect 67008 554810 67036 555183
rect 66996 554804 67048 554810
rect 66996 554746 67048 554752
rect 66994 553616 67050 553625
rect 66994 553551 67050 553560
rect 67008 553450 67036 553551
rect 66996 553444 67048 553450
rect 66996 553386 67048 553392
rect 66994 546816 67050 546825
rect 66994 546751 67050 546760
rect 67008 546514 67036 546751
rect 66996 546508 67048 546514
rect 66996 546450 67048 546456
rect 67364 434036 67416 434042
rect 67364 433978 67416 433984
rect 66996 422272 67048 422278
rect 66996 422214 67048 422220
rect 67008 421161 67036 422214
rect 66994 421152 67050 421161
rect 66994 421087 67050 421096
rect 66916 420158 67036 420186
rect 66902 420064 66958 420073
rect 66902 419999 66958 420008
rect 66916 419558 66944 419999
rect 66904 419552 66956 419558
rect 66904 419494 66956 419500
rect 67008 419370 67036 420158
rect 66916 419342 67036 419370
rect 66916 418266 66944 419342
rect 66904 418260 66956 418266
rect 66904 418202 66956 418208
rect 66916 417081 66944 418202
rect 67376 418169 67404 433978
rect 66994 418160 67050 418169
rect 66994 418095 67050 418104
rect 67362 418160 67418 418169
rect 67362 418095 67418 418104
rect 66902 417072 66958 417081
rect 66902 417007 66958 417016
rect 67008 416906 67036 418095
rect 66996 416900 67048 416906
rect 66996 416842 67048 416848
rect 66904 414792 66956 414798
rect 66904 414734 66956 414740
rect 66916 414089 66944 414734
rect 66902 414080 66958 414089
rect 66902 414015 66958 414024
rect 66904 413296 66956 413302
rect 66904 413238 66956 413244
rect 66916 413001 66944 413238
rect 66902 412992 66958 413001
rect 66902 412927 66958 412936
rect 66904 411256 66956 411262
rect 66904 411198 66956 411204
rect 66916 410825 66944 411198
rect 66902 410816 66958 410825
rect 66902 410751 66958 410760
rect 66904 408468 66956 408474
rect 66904 408410 66956 408416
rect 66916 407833 66944 408410
rect 66902 407824 66958 407833
rect 66902 407759 66958 407768
rect 67468 405657 67496 577215
rect 67560 575385 67588 589902
rect 67546 575376 67602 575385
rect 67546 575311 67602 575320
rect 67652 566681 67680 702986
rect 70320 582457 70348 703258
rect 72988 702982 73016 703520
rect 71780 702976 71832 702982
rect 71780 702918 71832 702924
rect 72976 702976 73028 702982
rect 72976 702918 73028 702924
rect 84108 702976 84160 702982
rect 84108 702918 84160 702924
rect 71688 700324 71740 700330
rect 71688 700266 71740 700272
rect 71700 589966 71728 700266
rect 71688 589960 71740 589966
rect 71688 589902 71740 589908
rect 71792 584905 71820 702918
rect 77208 702704 77260 702710
rect 77208 702646 77260 702652
rect 77220 591161 77248 702646
rect 76470 591152 76526 591161
rect 76470 591087 76526 591096
rect 77206 591152 77262 591161
rect 77206 591087 77262 591096
rect 71778 584896 71834 584905
rect 71778 584831 71834 584840
rect 73528 583772 73580 583778
rect 73528 583714 73580 583720
rect 72422 582720 72478 582729
rect 72422 582655 72478 582664
rect 69478 582448 69534 582457
rect 70306 582448 70362 582457
rect 69478 582383 69534 582392
rect 69940 582412 69992 582418
rect 69492 580938 69520 582383
rect 70306 582383 70362 582392
rect 69940 582354 69992 582360
rect 69664 581120 69716 581126
rect 69664 581062 69716 581068
rect 69952 581074 69980 582354
rect 72436 581074 72464 582655
rect 73540 581074 73568 583714
rect 73804 582480 73856 582486
rect 73804 582422 73856 582428
rect 74906 582448 74962 582457
rect 69032 580910 69520 580938
rect 69032 580802 69060 580910
rect 68664 580774 69060 580802
rect 68664 578921 68692 580774
rect 69676 580718 69704 581062
rect 69952 581046 70288 581074
rect 72128 581046 72464 581074
rect 73232 581046 73568 581074
rect 73816 581074 73844 582422
rect 74906 582383 74962 582392
rect 76288 582412 76340 582418
rect 73816 581046 74152 581074
rect 74920 580938 74948 582383
rect 76288 582354 76340 582360
rect 76300 581074 76328 582354
rect 75992 581046 76328 581074
rect 76484 581074 76512 591087
rect 77220 590753 77248 591087
rect 77206 590744 77262 590753
rect 77206 590679 77262 590688
rect 84120 587926 84148 702918
rect 86224 702772 86276 702778
rect 86224 702714 86276 702720
rect 84108 587920 84160 587926
rect 84108 587862 84160 587868
rect 78588 585812 78640 585818
rect 78588 585754 78640 585760
rect 78600 585206 78628 585754
rect 82728 585268 82780 585274
rect 82728 585210 82780 585216
rect 77944 585200 77996 585206
rect 77944 585142 77996 585148
rect 78588 585200 78640 585206
rect 78588 585142 78640 585148
rect 76484 581046 76912 581074
rect 75366 580952 75422 580961
rect 74920 580910 75366 580938
rect 75366 580887 75422 580896
rect 70858 580816 70914 580825
rect 77956 580802 77984 585142
rect 81808 582616 81860 582622
rect 81808 582558 81860 582564
rect 80244 581120 80296 581126
rect 79046 581088 79102 581097
rect 78752 581046 79046 581074
rect 81820 581074 81848 582558
rect 82740 581074 82768 585210
rect 84120 582622 84148 587862
rect 86236 586514 86264 702714
rect 89180 699718 89208 703520
rect 90364 703248 90416 703254
rect 90364 703190 90416 703196
rect 87604 699712 87656 699718
rect 87604 699654 87656 699660
rect 89168 699712 89220 699718
rect 89168 699654 89220 699660
rect 86500 586560 86552 586566
rect 86236 586508 86500 586514
rect 86236 586502 86552 586508
rect 86236 586486 86540 586502
rect 84108 582616 84160 582622
rect 84108 582558 84160 582564
rect 83002 581224 83058 581233
rect 83002 581159 83058 581168
rect 80296 581068 80592 581074
rect 80244 581062 80592 581068
rect 80256 581046 80592 581062
rect 81512 581046 81848 581074
rect 82432 581046 82768 581074
rect 83016 581074 83044 581159
rect 86512 581074 86540 586486
rect 87616 585818 87644 699654
rect 90376 596174 90404 703190
rect 102048 703112 102100 703118
rect 102048 703054 102100 703060
rect 97264 702840 97316 702846
rect 97264 702782 97316 702788
rect 94688 702636 94740 702642
rect 94688 702578 94740 702584
rect 90376 596146 90496 596174
rect 87604 585812 87656 585818
rect 87604 585754 87656 585760
rect 87512 585200 87564 585206
rect 87512 585142 87564 585148
rect 87524 581074 87552 585142
rect 88246 582584 88302 582593
rect 88246 582519 88302 582528
rect 87880 582412 87932 582418
rect 87880 582354 87932 582360
rect 87892 581670 87920 582354
rect 87880 581664 87932 581670
rect 87880 581606 87932 581612
rect 88260 581074 88288 582519
rect 90272 582412 90324 582418
rect 90272 582354 90324 582360
rect 90284 581074 90312 582354
rect 83016 581046 83352 581074
rect 86296 581046 86540 581074
rect 87216 581046 87552 581074
rect 88136 581046 88288 581074
rect 89976 581046 90312 581074
rect 90468 581074 90496 596146
rect 92112 583840 92164 583846
rect 92112 583782 92164 583788
rect 92124 581074 92152 583782
rect 93768 582480 93820 582486
rect 93768 582422 93820 582428
rect 90468 581052 90896 581074
rect 90468 581046 90548 581052
rect 79046 581023 79102 581032
rect 90600 581046 90896 581052
rect 91816 581046 92152 581074
rect 90548 580994 90600 581000
rect 93780 580938 93808 582422
rect 93656 580910 93808 580938
rect 79782 580816 79838 580825
rect 70914 580774 71208 580802
rect 77832 580774 77984 580802
rect 79672 580774 79782 580802
rect 70858 580751 70914 580760
rect 79782 580751 79838 580760
rect 84198 580816 84254 580825
rect 88706 580816 88762 580825
rect 84254 580774 84456 580802
rect 85376 580774 85528 580802
rect 84198 580751 84254 580760
rect 85500 580718 85528 580774
rect 92386 580816 92442 580825
rect 88762 580774 89056 580802
rect 88706 580751 88762 580760
rect 92442 580774 92736 580802
rect 92386 580751 92442 580760
rect 69664 580712 69716 580718
rect 69664 580654 69716 580660
rect 85488 580712 85540 580718
rect 85488 580654 85540 580660
rect 94700 580514 94728 702578
rect 95332 588600 95384 588606
rect 95332 588542 95384 588548
rect 94688 580508 94740 580514
rect 94688 580450 94740 580456
rect 94576 580366 94820 580394
rect 94688 580304 94740 580310
rect 94688 580246 94740 580252
rect 68650 578912 68706 578921
rect 68650 578847 68706 578856
rect 67638 566672 67694 566681
rect 67638 566607 67694 566616
rect 67652 565894 67680 566607
rect 67640 565888 67692 565894
rect 67640 565830 67692 565836
rect 67822 556608 67878 556617
rect 67822 556543 67878 556552
rect 67730 552256 67786 552265
rect 67730 552191 67786 552200
rect 67638 550896 67694 550905
rect 67638 550831 67694 550840
rect 67652 440910 67680 550831
rect 67744 539850 67772 552191
rect 67732 539844 67784 539850
rect 67732 539786 67784 539792
rect 67836 539578 67864 556543
rect 94700 552537 94728 580246
rect 94792 574802 94820 580366
rect 95238 574832 95294 574841
rect 94780 574796 94832 574802
rect 95238 574767 95294 574776
rect 94780 574738 94832 574744
rect 94778 563680 94834 563689
rect 94778 563615 94834 563624
rect 94686 552528 94742 552537
rect 94686 552463 94742 552472
rect 94686 540288 94742 540297
rect 94686 540223 94742 540232
rect 94700 539850 94728 540223
rect 71780 539844 71832 539850
rect 71780 539786 71832 539792
rect 93216 539844 93268 539850
rect 93216 539786 93268 539792
rect 94688 539844 94740 539850
rect 94688 539786 94740 539792
rect 70306 539744 70362 539753
rect 70306 539679 70308 539688
rect 70360 539679 70362 539688
rect 70308 539650 70360 539656
rect 67824 539572 67876 539578
rect 67824 539514 67876 539520
rect 68928 539572 68980 539578
rect 68928 539514 68980 539520
rect 67744 539158 68816 539186
rect 67744 478174 67772 539158
rect 68940 538898 68968 539514
rect 69400 539158 69736 539186
rect 70656 539158 70716 539186
rect 68928 538892 68980 538898
rect 68928 538834 68980 538840
rect 69400 536722 69428 539158
rect 70688 538218 70716 539158
rect 70780 539158 71576 539186
rect 70676 538212 70728 538218
rect 70676 538154 70728 538160
rect 70688 536858 70716 538154
rect 70676 536852 70728 536858
rect 70676 536794 70728 536800
rect 69388 536716 69440 536722
rect 69388 536658 69440 536664
rect 70780 528554 70808 539158
rect 71136 536852 71188 536858
rect 71136 536794 71188 536800
rect 70504 528526 70808 528554
rect 67732 478168 67784 478174
rect 67732 478110 67784 478116
rect 70504 466478 70532 528526
rect 71044 520940 71096 520946
rect 71044 520882 71096 520888
rect 70492 466472 70544 466478
rect 70492 466414 70544 466420
rect 67732 460216 67784 460222
rect 67732 460158 67784 460164
rect 67640 440904 67692 440910
rect 67640 440846 67692 440852
rect 67454 405648 67510 405657
rect 67454 405583 67510 405592
rect 66902 404560 66958 404569
rect 66902 404495 66958 404504
rect 66916 404394 66944 404495
rect 66904 404388 66956 404394
rect 66904 404330 66956 404336
rect 67468 402974 67496 405583
rect 66732 402946 66852 402974
rect 67284 402946 67496 402974
rect 66732 402665 66760 402946
rect 66718 402656 66774 402665
rect 66718 402591 66774 402600
rect 66534 399664 66590 399673
rect 66534 399599 66590 399608
rect 66548 398886 66576 399599
rect 66536 398880 66588 398886
rect 66536 398822 66588 398828
rect 66626 398576 66682 398585
rect 66626 398511 66682 398520
rect 66640 396846 66668 398511
rect 66732 397458 66760 402591
rect 66902 401568 66958 401577
rect 66902 401503 66958 401512
rect 66810 400480 66866 400489
rect 66810 400415 66866 400424
rect 66824 400314 66852 400415
rect 66812 400308 66864 400314
rect 66812 400250 66864 400256
rect 66916 400246 66944 401503
rect 66904 400240 66956 400246
rect 66904 400182 66956 400188
rect 66720 397452 66772 397458
rect 66720 397394 66772 397400
rect 66628 396840 66680 396846
rect 66628 396782 66680 396788
rect 67088 396704 67140 396710
rect 67088 396646 67140 396652
rect 67100 396409 67128 396646
rect 67086 396400 67142 396409
rect 67086 396335 67142 396344
rect 66812 396024 66864 396030
rect 66812 395966 66864 395972
rect 66824 395321 66852 395966
rect 66810 395312 66866 395321
rect 66810 395247 66866 395256
rect 66166 394632 66222 394641
rect 66166 394567 66222 394576
rect 66350 394496 66406 394505
rect 66350 394431 66406 394440
rect 66364 392630 66392 394431
rect 66810 393408 66866 393417
rect 66810 393343 66812 393352
rect 66864 393343 66866 393352
rect 66812 393314 66864 393320
rect 66352 392624 66404 392630
rect 66352 392566 66404 392572
rect 66810 392320 66866 392329
rect 66810 392255 66866 392264
rect 66824 392018 66852 392255
rect 66812 392012 66864 392018
rect 66812 391954 66864 391960
rect 66810 391232 66866 391241
rect 66810 391167 66866 391176
rect 66824 385694 66852 391167
rect 66812 385688 66864 385694
rect 66812 385630 66864 385636
rect 67284 312594 67312 402946
rect 67744 397905 67772 460158
rect 68926 449984 68982 449993
rect 68926 449919 68928 449928
rect 68980 449919 68982 449928
rect 68928 449890 68980 449896
rect 71056 436257 71084 520882
rect 71148 485110 71176 536794
rect 71136 485104 71188 485110
rect 71136 485046 71188 485052
rect 71136 437436 71188 437442
rect 71136 437378 71188 437384
rect 68926 436248 68982 436257
rect 68926 436183 68982 436192
rect 71042 436248 71098 436257
rect 71042 436183 71098 436192
rect 68468 435396 68520 435402
rect 68468 435338 68520 435344
rect 68376 433764 68428 433770
rect 68376 433706 68428 433712
rect 68388 432018 68416 433706
rect 68480 432562 68508 435338
rect 68940 434194 68968 436183
rect 71148 436150 71176 437378
rect 71136 436144 71188 436150
rect 69938 436112 69994 436121
rect 71136 436086 71188 436092
rect 69938 436047 69994 436056
rect 69952 434330 69980 436047
rect 69952 434302 70288 434330
rect 71148 434194 71176 436086
rect 71792 435402 71820 539786
rect 72332 539708 72384 539714
rect 72332 539650 72384 539656
rect 72344 538214 72372 539650
rect 76746 539608 76802 539617
rect 76802 539566 77096 539594
rect 76746 539543 76802 539552
rect 72496 539158 72832 539186
rect 73416 539158 73476 539186
rect 74336 539158 74488 539186
rect 72344 538186 72648 538214
rect 72620 476785 72648 538186
rect 72804 535498 72832 539158
rect 73448 536790 73476 539158
rect 73436 536784 73488 536790
rect 73436 536726 73488 536732
rect 73448 535770 73476 536726
rect 73436 535764 73488 535770
rect 73436 535706 73488 535712
rect 72792 535492 72844 535498
rect 72792 535434 72844 535440
rect 73804 535492 73856 535498
rect 73804 535434 73856 535440
rect 72606 476776 72662 476785
rect 72606 476711 72662 476720
rect 73816 472666 73844 535434
rect 74460 534721 74488 539158
rect 74552 539158 75256 539186
rect 76176 539158 76512 539186
rect 74446 534712 74502 534721
rect 74446 534647 74502 534656
rect 73804 472660 73856 472666
rect 73804 472602 73856 472608
rect 73988 436212 74040 436218
rect 73988 436154 74040 436160
rect 71780 435396 71832 435402
rect 71780 435338 71832 435344
rect 72700 435396 72752 435402
rect 72700 435338 72752 435344
rect 72608 434852 72660 434858
rect 72608 434794 72660 434800
rect 72620 434330 72648 434794
rect 72312 434302 72648 434330
rect 72712 434330 72740 435338
rect 73434 434752 73490 434761
rect 73434 434687 73490 434696
rect 73448 434330 73476 434687
rect 74000 434330 74028 436154
rect 72712 434302 73048 434330
rect 73448 434302 73784 434330
rect 74000 434302 74336 434330
rect 68816 434166 68968 434194
rect 71024 434166 71176 434194
rect 68652 433696 68704 433702
rect 68940 433673 68968 434166
rect 74552 434042 74580 539158
rect 76484 536761 76512 539158
rect 76470 536752 76526 536761
rect 76470 536687 76526 536696
rect 76484 535673 76512 536687
rect 76564 535764 76616 535770
rect 76564 535706 76616 535712
rect 76470 535664 76526 535673
rect 76470 535599 76526 535608
rect 76102 535528 76158 535537
rect 76102 535463 76158 535472
rect 75184 526448 75236 526454
rect 75184 526390 75236 526396
rect 74724 438184 74776 438190
rect 74724 438126 74776 438132
rect 74736 434353 74764 438126
rect 75196 437442 75224 526390
rect 76116 441697 76144 535463
rect 76576 522345 76604 535706
rect 76760 535537 76788 539543
rect 77312 539158 78016 539186
rect 78692 539158 78936 539186
rect 80040 539158 80192 539186
rect 77206 535664 77262 535673
rect 77206 535599 77262 535608
rect 76746 535528 76802 535537
rect 76746 535463 76802 535472
rect 76562 522336 76618 522345
rect 76562 522271 76618 522280
rect 77220 473346 77248 535599
rect 77208 473340 77260 473346
rect 77208 473282 77260 473288
rect 77312 442270 77340 539158
rect 77944 473340 77996 473346
rect 77944 473282 77996 473288
rect 77300 442264 77352 442270
rect 77300 442206 77352 442212
rect 76102 441688 76158 441697
rect 76102 441623 76158 441632
rect 75184 437436 75236 437442
rect 75184 437378 75236 437384
rect 77390 437200 77446 437209
rect 77390 437135 77446 437144
rect 77404 436257 77432 437135
rect 77482 436384 77538 436393
rect 77482 436319 77538 436328
rect 77390 436248 77446 436257
rect 77390 436183 77446 436192
rect 76840 436144 76892 436150
rect 76840 436086 76892 436092
rect 74722 434344 74778 434353
rect 76194 434344 76250 434353
rect 74778 434302 75072 434330
rect 74722 434279 74778 434288
rect 76852 434330 76880 436086
rect 76250 434302 76880 434330
rect 76194 434279 76250 434288
rect 74736 434219 74764 434279
rect 77404 434194 77432 436183
rect 77496 434330 77524 436319
rect 77956 436218 77984 473282
rect 78692 449274 78720 539158
rect 80060 533384 80112 533390
rect 80060 533326 80112 533332
rect 79324 451920 79376 451926
rect 79324 451862 79376 451868
rect 78680 449268 78732 449274
rect 78680 449210 78732 449216
rect 78036 447908 78088 447914
rect 78036 447850 78088 447856
rect 78048 437209 78076 447850
rect 78404 440972 78456 440978
rect 78404 440914 78456 440920
rect 78416 437481 78444 440914
rect 78402 437472 78458 437481
rect 78402 437407 78458 437416
rect 78034 437200 78090 437209
rect 78034 437135 78090 437144
rect 77944 436212 77996 436218
rect 77944 436154 77996 436160
rect 79336 436150 79364 451862
rect 80072 450537 80100 533326
rect 80164 487830 80192 539158
rect 80624 539158 80960 539186
rect 81452 539158 81880 539186
rect 82800 539158 82860 539186
rect 83720 539158 84056 539186
rect 80624 533390 80652 539158
rect 80612 533384 80664 533390
rect 80612 533326 80664 533332
rect 80152 487824 80204 487830
rect 80152 487766 80204 487772
rect 81452 479505 81480 539158
rect 81438 479496 81494 479505
rect 81438 479431 81494 479440
rect 82832 467158 82860 539158
rect 82912 538892 82964 538898
rect 82912 538834 82964 538840
rect 82820 467152 82872 467158
rect 82820 467094 82872 467100
rect 80058 450528 80114 450537
rect 80058 450463 80114 450472
rect 80060 449948 80112 449954
rect 80060 449890 80112 449896
rect 79324 436144 79376 436150
rect 79324 436086 79376 436092
rect 80072 434602 80100 449890
rect 81440 443760 81492 443766
rect 81440 443702 81492 443708
rect 81452 441614 81480 443702
rect 82924 441614 82952 538834
rect 84028 533390 84056 539158
rect 84304 539158 84640 539186
rect 85560 539158 85620 539186
rect 86480 539158 86908 539186
rect 84304 533458 84332 539158
rect 84292 533452 84344 533458
rect 84292 533394 84344 533400
rect 84016 533384 84068 533390
rect 84016 533326 84068 533332
rect 85488 475176 85540 475182
rect 85488 475118 85540 475124
rect 85500 441614 85528 475118
rect 85592 463010 85620 539158
rect 86880 536790 86908 539158
rect 86972 539158 87400 539186
rect 88320 539158 88472 539186
rect 86868 536784 86920 536790
rect 86868 536726 86920 536732
rect 86316 464364 86368 464370
rect 86316 464306 86368 464312
rect 85580 463004 85632 463010
rect 85580 462946 85632 462952
rect 85672 449200 85724 449206
rect 85672 449142 85724 449148
rect 81452 441586 81664 441614
rect 82924 441586 83228 441614
rect 81346 438152 81402 438161
rect 81346 438087 81402 438096
rect 80242 435296 80298 435305
rect 80242 435231 80298 435240
rect 80026 434574 80100 434602
rect 77496 434302 77832 434330
rect 80026 434316 80054 434574
rect 80256 434330 80284 435231
rect 81360 434489 81388 438087
rect 81346 434480 81402 434489
rect 81402 434438 81480 434466
rect 81346 434415 81402 434424
rect 80256 434302 80592 434330
rect 81452 434194 81480 434438
rect 81636 434330 81664 441586
rect 82912 436212 82964 436218
rect 82912 436154 82964 436160
rect 81636 434302 82064 434330
rect 77280 434166 77432 434194
rect 81328 434166 81480 434194
rect 74540 434036 74592 434042
rect 74540 433978 74592 433984
rect 82924 433786 82952 436154
rect 83200 433809 83228 441586
rect 85224 441586 85528 441614
rect 85684 441614 85712 449142
rect 85684 441586 85896 441614
rect 83738 436112 83794 436121
rect 83738 436047 83794 436056
rect 83752 434330 83780 436047
rect 83752 434302 84088 434330
rect 83186 433800 83242 433809
rect 71240 433770 71576 433786
rect 71228 433764 71576 433770
rect 71280 433758 71576 433764
rect 82800 433758 83136 433786
rect 71228 433706 71280 433712
rect 69204 433696 69256 433702
rect 68652 433638 68704 433644
rect 68926 433664 68982 433673
rect 68664 432857 68692 433638
rect 83108 433673 83136 433758
rect 83242 433758 83536 433786
rect 83186 433735 83242 433744
rect 75458 433664 75514 433673
rect 69256 433644 69552 433650
rect 69204 433638 69552 433644
rect 69216 433622 69552 433638
rect 68926 433599 68982 433608
rect 78218 433664 78274 433673
rect 75514 433622 75808 433650
rect 75458 433599 75514 433608
rect 78954 433664 79010 433673
rect 78274 433622 78568 433650
rect 78218 433599 78274 433608
rect 83094 433664 83150 433673
rect 79010 433622 79304 433650
rect 78954 433599 79010 433608
rect 83094 433599 83150 433608
rect 84474 433664 84530 433673
rect 85224 433650 85252 441586
rect 85868 437474 85896 441586
rect 85868 437446 85988 437474
rect 85670 436112 85726 436121
rect 85670 436047 85726 436056
rect 85684 433673 85712 436047
rect 85960 433673 85988 437446
rect 86328 436121 86356 464306
rect 86880 457570 86908 536726
rect 86868 457564 86920 457570
rect 86868 457506 86920 457512
rect 86972 457502 87000 539158
rect 88248 538348 88300 538354
rect 88248 538290 88300 538296
rect 86960 457496 87012 457502
rect 86960 457438 87012 457444
rect 88260 436121 88288 538290
rect 88340 533452 88392 533458
rect 88340 533394 88392 533400
rect 88352 447846 88380 533394
rect 88444 468625 88472 539158
rect 88904 539158 89240 539186
rect 90160 539158 90404 539186
rect 88904 533458 88932 539158
rect 90376 538218 90404 539158
rect 91112 539158 91264 539186
rect 91572 539158 92184 539186
rect 92768 539158 93104 539186
rect 90364 538212 90416 538218
rect 90364 538154 90416 538160
rect 88892 533452 88944 533458
rect 88892 533394 88944 533400
rect 88430 468616 88486 468625
rect 88430 468551 88486 468560
rect 90376 451926 90404 538154
rect 91008 535492 91060 535498
rect 91008 535434 91060 535440
rect 90364 451920 90416 451926
rect 90364 451862 90416 451868
rect 88340 447840 88392 447846
rect 88340 447782 88392 447788
rect 91020 446486 91048 535434
rect 91112 447914 91140 539158
rect 91572 528554 91600 539158
rect 92768 535498 92796 539158
rect 92756 535492 92808 535498
rect 92756 535434 92808 535440
rect 91204 528526 91600 528554
rect 91204 520946 91232 528526
rect 91192 520940 91244 520946
rect 91192 520882 91244 520888
rect 93228 475182 93256 539786
rect 94024 539158 94544 539186
rect 93950 538928 94006 538937
rect 93950 538863 94006 538872
rect 93964 538286 93992 538863
rect 93952 538280 94004 538286
rect 93952 538222 94004 538228
rect 94516 534750 94544 539158
rect 94504 534744 94556 534750
rect 94504 534686 94556 534692
rect 93216 475176 93268 475182
rect 93216 475118 93268 475124
rect 92572 458856 92624 458862
rect 92572 458798 92624 458804
rect 91100 447908 91152 447914
rect 91100 447850 91152 447856
rect 91008 446480 91060 446486
rect 91008 446422 91060 446428
rect 88432 443692 88484 443698
rect 88432 443634 88484 443640
rect 88444 440337 88472 443634
rect 88430 440328 88486 440337
rect 88430 440263 88486 440272
rect 88444 437474 88472 440263
rect 88444 437446 88656 437474
rect 86314 436112 86370 436121
rect 86314 436047 86370 436056
rect 87142 436112 87198 436121
rect 87142 436047 87198 436056
rect 88246 436112 88302 436121
rect 88246 436047 88302 436056
rect 87156 433673 87184 436047
rect 88628 434330 88656 437446
rect 89902 436248 89958 436257
rect 89902 436183 89958 436192
rect 88628 434302 89056 434330
rect 89916 434058 89944 436183
rect 92584 434602 92612 458798
rect 93860 443012 93912 443018
rect 93860 442954 93912 442960
rect 93872 434602 93900 442954
rect 94516 437617 94544 534686
rect 94792 474065 94820 563615
rect 95148 546508 95200 546514
rect 95148 546450 95200 546456
rect 94778 474056 94834 474065
rect 94778 473991 94834 474000
rect 95160 443018 95188 546450
rect 95252 464370 95280 574767
rect 95344 558929 95372 588542
rect 96620 587172 96672 587178
rect 96620 587114 96672 587120
rect 96250 574832 96306 574841
rect 96250 574767 96306 574776
rect 96264 574122 96292 574767
rect 96252 574116 96304 574122
rect 96252 574058 96304 574064
rect 96632 569129 96660 587114
rect 96894 578912 96950 578921
rect 96894 578847 96950 578856
rect 96908 578270 96936 578847
rect 96896 578264 96948 578270
rect 96896 578206 96948 578212
rect 97078 577552 97134 577561
rect 97078 577487 97134 577496
rect 97092 576910 97120 577487
rect 97080 576904 97132 576910
rect 97080 576846 97132 576852
rect 97276 572257 97304 702782
rect 101404 587920 101456 587926
rect 101404 587862 101456 587868
rect 98644 585268 98696 585274
rect 98644 585210 98696 585216
rect 97908 576768 97960 576774
rect 97906 576736 97908 576745
rect 97960 576736 97962 576745
rect 97906 576671 97962 576680
rect 97906 573472 97962 573481
rect 97962 573430 98040 573458
rect 97906 573407 97962 573416
rect 97262 572248 97318 572257
rect 97262 572183 97318 572192
rect 96618 569120 96674 569129
rect 96618 569055 96674 569064
rect 95422 565856 95478 565865
rect 95422 565791 95478 565800
rect 95330 558920 95386 558929
rect 95330 558855 95386 558864
rect 95330 555520 95386 555529
rect 95330 555455 95386 555464
rect 95344 523705 95372 555455
rect 95436 538354 95464 565791
rect 96802 560960 96858 560969
rect 96802 560895 96858 560904
rect 95882 558920 95938 558929
rect 95882 558855 95938 558864
rect 95424 538348 95476 538354
rect 95424 538290 95476 538296
rect 95330 523696 95386 523705
rect 95330 523631 95386 523640
rect 95240 464364 95292 464370
rect 95240 464306 95292 464312
rect 95896 444446 95924 558855
rect 96710 556880 96766 556889
rect 96710 556815 96766 556824
rect 96618 552120 96674 552129
rect 96618 552055 96674 552064
rect 96632 547874 96660 552055
rect 96724 551834 96752 556815
rect 96816 551954 96844 560895
rect 97276 558210 97304 572183
rect 97906 570072 97962 570081
rect 97906 570007 97962 570016
rect 97920 569974 97948 570007
rect 97908 569968 97960 569974
rect 97908 569910 97960 569916
rect 97908 569220 97960 569226
rect 97908 569162 97960 569168
rect 97920 569129 97948 569162
rect 97906 569120 97962 569129
rect 97906 569055 97962 569064
rect 97354 562320 97410 562329
rect 97354 562255 97410 562264
rect 97264 558204 97316 558210
rect 97264 558146 97316 558152
rect 97368 555490 97396 562255
rect 97356 555484 97408 555490
rect 97356 555426 97408 555432
rect 96894 554160 96950 554169
rect 96894 554095 96950 554104
rect 96908 551970 96936 554095
rect 96986 552800 97042 552809
rect 96986 552735 97042 552744
rect 97000 552090 97028 552735
rect 96988 552084 97040 552090
rect 96988 552026 97040 552032
rect 96804 551948 96856 551954
rect 96908 551942 97028 551970
rect 96804 551890 96856 551896
rect 96724 551806 96936 551834
rect 96804 551744 96856 551750
rect 96804 551686 96856 551692
rect 96632 547846 96752 547874
rect 96724 546514 96752 547846
rect 96712 546508 96764 546514
rect 96712 546450 96764 546456
rect 96710 545728 96766 545737
rect 96710 545663 96766 545672
rect 96724 460222 96752 545663
rect 96816 526454 96844 551686
rect 96908 537538 96936 551806
rect 96896 537532 96948 537538
rect 96896 537474 96948 537480
rect 96804 526448 96856 526454
rect 96804 526390 96856 526396
rect 96712 460216 96764 460222
rect 96712 460158 96764 460164
rect 95976 446412 96028 446418
rect 95976 446354 96028 446360
rect 95884 444440 95936 444446
rect 95884 444382 95936 444388
rect 95148 443012 95200 443018
rect 95148 442954 95200 442960
rect 94502 437608 94558 437617
rect 94502 437543 94558 437552
rect 95988 437510 96016 446354
rect 96528 444440 96580 444446
rect 96528 444382 96580 444388
rect 96540 443766 96568 444382
rect 96528 443760 96580 443766
rect 96528 443702 96580 443708
rect 95976 437504 96028 437510
rect 95976 437446 96028 437452
rect 94410 436112 94466 436121
rect 94410 436047 94466 436056
rect 92538 434574 92612 434602
rect 93826 434574 93900 434602
rect 92538 434194 92566 434574
rect 93826 434316 93854 434574
rect 94424 434330 94452 436047
rect 95284 434616 95340 434625
rect 95988 434602 96016 437446
rect 95988 434574 96062 434602
rect 95284 434551 95340 434560
rect 94778 434344 94834 434353
rect 94424 434302 94778 434330
rect 95298 434316 95326 434551
rect 96034 434316 96062 434574
rect 96342 434344 96398 434353
rect 94778 434279 94834 434288
rect 97000 434330 97028 551942
rect 97906 550760 97962 550769
rect 97906 550695 97962 550704
rect 97920 550662 97948 550695
rect 97908 550656 97960 550662
rect 97908 550598 97960 550604
rect 97538 544368 97594 544377
rect 97538 544303 97594 544312
rect 97552 543794 97580 544303
rect 97540 543788 97592 543794
rect 97540 543730 97592 543736
rect 98012 518226 98040 573430
rect 98090 543008 98146 543017
rect 98090 542943 98146 542952
rect 98104 532030 98132 542943
rect 98092 532024 98144 532030
rect 98092 531966 98144 531972
rect 98000 518220 98052 518226
rect 98000 518162 98052 518168
rect 98656 439521 98684 585210
rect 100022 582584 100078 582593
rect 100022 582519 100078 582528
rect 98736 478168 98788 478174
rect 98736 478110 98788 478116
rect 98642 439512 98698 439521
rect 98642 439447 98698 439456
rect 97078 437472 97134 437481
rect 97078 437407 97134 437416
rect 96398 434302 97028 434330
rect 97092 434330 97120 437407
rect 98748 436150 98776 478110
rect 100036 443698 100064 582519
rect 101416 449206 101444 587862
rect 102060 576978 102088 703054
rect 105464 700330 105492 703520
rect 119344 703180 119396 703186
rect 119344 703122 119396 703128
rect 116584 702772 116636 702778
rect 116584 702714 116636 702720
rect 105636 702636 105688 702642
rect 105636 702578 105688 702584
rect 105452 700324 105504 700330
rect 105452 700266 105504 700272
rect 105544 582480 105596 582486
rect 105544 582422 105596 582428
rect 103520 582412 103572 582418
rect 103520 582354 103572 582360
rect 102782 581088 102838 581097
rect 102782 581023 102838 581032
rect 102048 576972 102100 576978
rect 102048 576914 102100 576920
rect 102060 576774 102088 576914
rect 102048 576768 102100 576774
rect 102048 576710 102100 576716
rect 101496 449268 101548 449274
rect 101496 449210 101548 449216
rect 101404 449200 101456 449206
rect 101404 449142 101456 449148
rect 100024 443692 100076 443698
rect 100024 443634 100076 443640
rect 100758 436384 100814 436393
rect 100758 436319 100814 436328
rect 98736 436144 98788 436150
rect 98736 436086 98788 436092
rect 99932 436144 99984 436150
rect 99932 436086 99984 436092
rect 97092 434302 97336 434330
rect 96342 434279 96398 434288
rect 92662 434208 92718 434217
rect 92538 434180 92662 434194
rect 92552 434166 92662 434180
rect 92662 434143 92718 434152
rect 96986 434208 97042 434217
rect 97092 434194 97120 434302
rect 97042 434166 97120 434194
rect 96986 434143 97042 434152
rect 89792 434030 89944 434058
rect 91466 433936 91522 433945
rect 99194 433936 99250 433945
rect 91522 433894 91816 433922
rect 91466 433871 91522 433880
rect 99250 433894 99544 433922
rect 99194 433871 99250 433880
rect 87326 433800 87382 433809
rect 92938 433800 92994 433809
rect 87382 433758 87584 433786
rect 87326 433735 87382 433744
rect 98366 433800 98422 433809
rect 92994 433758 93288 433786
rect 98072 433758 98366 433786
rect 92938 433735 92994 433744
rect 98366 433735 98422 433744
rect 99944 433673 99972 436086
rect 100772 434714 100800 436319
rect 101508 436150 101536 449210
rect 102796 439006 102824 581023
rect 103532 442950 103560 582354
rect 104348 457564 104400 457570
rect 104348 457506 104400 457512
rect 103520 442944 103572 442950
rect 103520 442886 103572 442892
rect 103532 441614 103560 442886
rect 103532 441586 103928 441614
rect 102600 439000 102652 439006
rect 102600 438942 102652 438948
rect 102784 439000 102836 439006
rect 102784 438942 102836 438948
rect 101496 436144 101548 436150
rect 101496 436086 101548 436092
rect 100680 434686 100800 434714
rect 100680 434058 100708 434686
rect 102612 434330 102640 438942
rect 103334 436384 103390 436393
rect 103334 436319 103390 436328
rect 103348 436121 103376 436319
rect 103704 436144 103756 436150
rect 103334 436112 103390 436121
rect 103704 436086 103756 436092
rect 103334 436047 103390 436056
rect 102304 434302 102640 434330
rect 103716 434058 103744 436086
rect 100680 434030 100832 434058
rect 103592 434030 103744 434058
rect 85670 433664 85726 433673
rect 84530 433622 85252 433650
rect 85560 433622 85670 433650
rect 84474 433599 84530 433608
rect 85670 433599 85726 433608
rect 85946 433664 86002 433673
rect 87142 433664 87198 433673
rect 86002 433622 86296 433650
rect 87032 433622 87142 433650
rect 85946 433599 86002 433608
rect 87142 433599 87198 433608
rect 87970 433664 88026 433673
rect 89994 433664 90050 433673
rect 88026 433622 88320 433650
rect 87970 433599 88026 433608
rect 91374 433664 91430 433673
rect 90050 433622 90344 433650
rect 91080 433622 91374 433650
rect 89994 433599 90050 433608
rect 91374 433599 91430 433608
rect 98458 433664 98514 433673
rect 99930 433664 99986 433673
rect 98514 433622 98808 433650
rect 98458 433599 98514 433608
rect 101218 433664 101274 433673
rect 99986 433622 100096 433650
rect 99930 433599 99986 433608
rect 102690 433664 102746 433673
rect 101274 433622 101568 433650
rect 101218 433599 101274 433608
rect 103900 433650 103928 441586
rect 104360 436121 104388 457506
rect 105556 441614 105584 582422
rect 105648 574122 105676 702578
rect 111064 583772 111116 583778
rect 111064 583714 111116 583720
rect 108304 581664 108356 581670
rect 108304 581606 108356 581612
rect 105636 574116 105688 574122
rect 105636 574058 105688 574064
rect 107568 570648 107620 570654
rect 107568 570590 107620 570596
rect 107580 569974 107608 570590
rect 107568 569968 107620 569974
rect 107568 569910 107620 569916
rect 106924 454708 106976 454714
rect 106924 454650 106976 454656
rect 106936 442338 106964 454650
rect 106280 442332 106332 442338
rect 106280 442274 106332 442280
rect 106924 442332 106976 442338
rect 106924 442274 106976 442280
rect 106292 441658 106320 442274
rect 106280 441652 106332 441658
rect 105556 441586 105952 441614
rect 106280 441594 106332 441600
rect 104898 436248 104954 436257
rect 104898 436183 104954 436192
rect 104346 436112 104402 436121
rect 104346 436047 104402 436056
rect 104912 434330 104940 436183
rect 104912 434302 105064 434330
rect 105924 434042 105952 441586
rect 106292 434602 106320 441594
rect 107580 437481 107608 569910
rect 108120 438932 108172 438938
rect 108120 438874 108172 438880
rect 107566 437472 107622 437481
rect 107566 437407 107622 437416
rect 106292 434574 106366 434602
rect 106338 434316 106366 434574
rect 108132 434330 108160 438874
rect 108316 437578 108344 581606
rect 109684 552084 109736 552090
rect 109684 552026 109736 552032
rect 108396 543788 108448 543794
rect 108396 543730 108448 543736
rect 108408 438938 108436 543730
rect 109696 521626 109724 552026
rect 109684 521620 109736 521626
rect 109684 521562 109736 521568
rect 109040 467152 109092 467158
rect 109040 467094 109092 467100
rect 109052 441614 109080 467094
rect 109052 441586 109448 441614
rect 108396 438932 108448 438938
rect 108396 438874 108448 438880
rect 108304 437572 108356 437578
rect 108304 437514 108356 437520
rect 107824 434302 108160 434330
rect 108316 434330 108344 437514
rect 109420 434353 109448 441586
rect 110418 436384 110474 436393
rect 110418 436319 110474 436328
rect 109406 434344 109462 434353
rect 108316 434302 108560 434330
rect 110432 434330 110460 436319
rect 111076 436150 111104 583714
rect 113456 579692 113508 579698
rect 113456 579634 113508 579640
rect 111800 521620 111852 521626
rect 111800 521562 111852 521568
rect 111064 436144 111116 436150
rect 111064 436086 111116 436092
rect 111076 434330 111104 436086
rect 111812 434790 111840 521562
rect 113272 447840 113324 447846
rect 113272 447782 113324 447788
rect 111800 434784 111852 434790
rect 111800 434726 111852 434732
rect 112444 434784 112496 434790
rect 112444 434726 112496 434732
rect 109462 434302 109848 434330
rect 110432 434302 110584 434330
rect 111076 434302 111320 434330
rect 109406 434279 109462 434288
rect 109420 434219 109448 434279
rect 108946 434072 109002 434081
rect 105912 434036 105964 434042
rect 112456 434058 112484 434726
rect 109002 434030 109296 434058
rect 112456 434030 112608 434058
rect 108946 434007 109002 434016
rect 105912 433978 105964 433984
rect 110880 433696 110932 433702
rect 104162 433664 104218 433673
rect 102746 433622 103040 433650
rect 103900 433622 104162 433650
rect 102690 433599 102746 433608
rect 105450 433664 105506 433673
rect 104218 433622 104328 433650
rect 104162 433599 104218 433608
rect 106738 433664 106794 433673
rect 105506 433622 105800 433650
rect 105450 433599 105506 433608
rect 110878 433664 110880 433673
rect 110932 433664 110934 433673
rect 106794 433622 107088 433650
rect 106738 433599 106794 433608
rect 110878 433599 110934 433608
rect 111890 433664 111946 433673
rect 111946 433622 112056 433650
rect 111890 433599 111946 433608
rect 112720 433288 112772 433294
rect 112720 433230 112772 433236
rect 68650 432848 68706 432857
rect 68650 432783 68706 432792
rect 68480 432534 68692 432562
rect 68388 431990 68600 432018
rect 67730 397896 67786 397905
rect 67730 397831 67786 397840
rect 67744 397594 67772 397831
rect 67364 397588 67416 397594
rect 67364 397530 67416 397536
rect 67732 397588 67784 397594
rect 67732 397530 67784 397536
rect 67272 312588 67324 312594
rect 67272 312530 67324 312536
rect 67284 312225 67312 312530
rect 67270 312216 67326 312225
rect 67270 312151 67326 312160
rect 66902 312080 66958 312089
rect 66902 312015 66958 312024
rect 66916 291145 66944 312015
rect 67376 309126 67404 397530
rect 67732 397452 67784 397458
rect 67732 397394 67784 397400
rect 67454 396400 67510 396409
rect 67454 396335 67510 396344
rect 67364 309120 67416 309126
rect 67364 309062 67416 309068
rect 66442 291136 66498 291145
rect 66442 291071 66498 291080
rect 66902 291136 66958 291145
rect 66902 291071 66958 291080
rect 66456 290465 66484 291071
rect 66442 290456 66498 290465
rect 66442 290391 66498 290400
rect 66812 283620 66864 283626
rect 66812 283562 66864 283568
rect 66168 283076 66220 283082
rect 66168 283018 66220 283024
rect 66074 271960 66130 271969
rect 66074 271895 66130 271904
rect 66074 252784 66130 252793
rect 66074 252719 66130 252728
rect 65984 251388 66036 251394
rect 65984 251330 66036 251336
rect 65892 233232 65944 233238
rect 65892 233174 65944 233180
rect 65982 147792 66038 147801
rect 65982 147727 66038 147736
rect 65890 144800 65946 144809
rect 65890 144735 65946 144744
rect 65904 143721 65932 144735
rect 65890 143712 65946 143721
rect 65890 143647 65946 143656
rect 65904 114617 65932 143647
rect 65996 118425 66024 147727
rect 66088 143614 66116 252719
rect 66180 241534 66208 283018
rect 66824 282985 66852 283562
rect 66810 282976 66866 282985
rect 66810 282911 66866 282920
rect 67272 280220 67324 280226
rect 67272 280162 67324 280168
rect 66536 279472 66588 279478
rect 66536 279414 66588 279420
rect 66548 278905 66576 279414
rect 66534 278896 66590 278905
rect 66534 278831 66590 278840
rect 66810 278080 66866 278089
rect 66810 278015 66812 278024
rect 66864 278015 66866 278024
rect 66812 277986 66864 277992
rect 66904 277364 66956 277370
rect 66904 277306 66956 277312
rect 66810 277264 66866 277273
rect 66810 277199 66866 277208
rect 66824 276214 66852 277199
rect 66916 276457 66944 277306
rect 66902 276448 66958 276457
rect 66902 276383 66958 276392
rect 66812 276208 66864 276214
rect 66812 276150 66864 276156
rect 66628 276004 66680 276010
rect 66628 275946 66680 275952
rect 66640 275641 66668 275946
rect 66626 275632 66682 275641
rect 66626 275567 66682 275576
rect 66810 273184 66866 273193
rect 66810 273119 66866 273128
rect 66824 272542 66852 273119
rect 66812 272536 66864 272542
rect 66812 272478 66864 272484
rect 66260 271176 66312 271182
rect 66260 271118 66312 271124
rect 66272 270745 66300 271118
rect 66258 270736 66314 270745
rect 66258 270671 66314 270680
rect 66272 269822 66300 270671
rect 66260 269816 66312 269822
rect 66260 269758 66312 269764
rect 66810 268288 66866 268297
rect 66810 268223 66866 268232
rect 66824 267782 66852 268223
rect 66812 267776 66864 267782
rect 66812 267718 66864 267724
rect 66810 266656 66866 266665
rect 66810 266591 66866 266600
rect 66824 266422 66852 266591
rect 66812 266416 66864 266422
rect 66812 266358 66864 266364
rect 66904 263560 66956 263566
rect 66904 263502 66956 263508
rect 66916 263401 66944 263502
rect 66902 263392 66958 263401
rect 66902 263327 66958 263336
rect 66536 262880 66588 262886
rect 66536 262822 66588 262828
rect 66548 262585 66576 262822
rect 66534 262576 66590 262585
rect 66534 262511 66590 262520
rect 66260 261520 66312 261526
rect 66260 261462 66312 261468
rect 66272 260953 66300 261462
rect 66258 260944 66314 260953
rect 66258 260879 66314 260888
rect 66272 260166 66300 260879
rect 66812 260228 66864 260234
rect 66812 260170 66864 260176
rect 66260 260160 66312 260166
rect 66824 260137 66852 260170
rect 66260 260102 66312 260108
rect 66810 260128 66866 260137
rect 66810 260063 66866 260072
rect 66444 259412 66496 259418
rect 66444 259354 66496 259360
rect 66260 258732 66312 258738
rect 66260 258674 66312 258680
rect 66272 256873 66300 258674
rect 66456 258097 66484 259354
rect 66442 258088 66498 258097
rect 66442 258023 66498 258032
rect 66810 257680 66866 257689
rect 66810 257615 66866 257624
rect 66824 257378 66852 257615
rect 66812 257372 66864 257378
rect 66812 257314 66864 257320
rect 66258 256864 66314 256873
rect 66258 256799 66314 256808
rect 66810 256048 66866 256057
rect 66810 255983 66866 255992
rect 66824 255338 66852 255983
rect 66812 255332 66864 255338
rect 66812 255274 66864 255280
rect 66812 254584 66864 254590
rect 66812 254526 66864 254532
rect 66824 254425 66852 254526
rect 66810 254416 66866 254425
rect 66810 254351 66866 254360
rect 66536 253904 66588 253910
rect 66536 253846 66588 253852
rect 66548 252793 66576 253846
rect 66534 252784 66590 252793
rect 66534 252719 66590 252728
rect 66258 251968 66314 251977
rect 66258 251903 66314 251912
rect 66272 251394 66300 251903
rect 66260 251388 66312 251394
rect 66260 251330 66312 251336
rect 66810 251152 66866 251161
rect 66810 251087 66866 251096
rect 66904 251116 66956 251122
rect 66824 250782 66852 251087
rect 66904 251058 66956 251064
rect 66812 250776 66864 250782
rect 66812 250718 66864 250724
rect 66916 250345 66944 251058
rect 66902 250336 66958 250345
rect 66902 250271 66958 250280
rect 66810 248704 66866 248713
rect 66810 248639 66866 248648
rect 66824 248470 66852 248639
rect 66812 248464 66864 248470
rect 66812 248406 66864 248412
rect 66904 248396 66956 248402
rect 66904 248338 66956 248344
rect 66916 247897 66944 248338
rect 66902 247888 66958 247897
rect 66902 247823 66958 247832
rect 67178 247072 67234 247081
rect 67178 247007 67234 247016
rect 66812 246356 66864 246362
rect 66812 246298 66864 246304
rect 66258 243808 66314 243817
rect 66258 243743 66314 243752
rect 66272 242962 66300 243743
rect 66824 243001 66852 246298
rect 66810 242992 66866 243001
rect 66260 242956 66312 242962
rect 66810 242927 66866 242936
rect 66260 242898 66312 242904
rect 66168 241528 66220 241534
rect 66168 241470 66220 241476
rect 66166 226400 66222 226409
rect 66166 226335 66222 226344
rect 66076 143608 66128 143614
rect 66076 143550 66128 143556
rect 65982 118416 66038 118425
rect 65982 118351 66038 118360
rect 65890 114608 65946 114617
rect 65890 114543 65946 114552
rect 65984 105596 66036 105602
rect 65984 105538 66036 105544
rect 64788 102400 64840 102406
rect 64788 102342 64840 102348
rect 64788 100020 64840 100026
rect 64788 99962 64840 99968
rect 64602 92440 64658 92449
rect 64602 92375 64658 92384
rect 64512 91044 64564 91050
rect 64512 90986 64564 90992
rect 63316 81388 63368 81394
rect 63316 81330 63368 81336
rect 64800 80034 64828 99962
rect 65996 82793 66024 105538
rect 66088 103193 66116 143550
rect 66180 111625 66208 226335
rect 66352 133204 66404 133210
rect 66352 133146 66404 133152
rect 66260 132456 66312 132462
rect 66260 132398 66312 132404
rect 66272 132025 66300 132398
rect 66258 132016 66314 132025
rect 66258 131951 66314 131960
rect 66364 131209 66392 133146
rect 66350 131200 66406 131209
rect 66350 131135 66406 131144
rect 66812 128308 66864 128314
rect 66812 128250 66864 128256
rect 66824 127673 66852 128250
rect 66810 127664 66866 127673
rect 66810 127599 66866 127608
rect 66812 126948 66864 126954
rect 66812 126890 66864 126896
rect 66824 126041 66852 126890
rect 66810 126032 66866 126041
rect 66810 125967 66866 125976
rect 66812 125588 66864 125594
rect 66812 125530 66864 125536
rect 66824 124409 66852 125530
rect 66904 124976 66956 124982
rect 66904 124918 66956 124924
rect 66810 124400 66866 124409
rect 66810 124335 66866 124344
rect 66628 124160 66680 124166
rect 66628 124102 66680 124108
rect 66640 123049 66668 124102
rect 66916 123865 66944 124918
rect 66902 123856 66958 123865
rect 66902 123791 66958 123800
rect 66626 123040 66682 123049
rect 66626 122975 66682 122984
rect 66812 122800 66864 122806
rect 66812 122742 66864 122748
rect 66824 122233 66852 122742
rect 66810 122224 66866 122233
rect 66810 122159 66866 122168
rect 66812 121440 66864 121446
rect 66810 121408 66812 121417
rect 66864 121408 66866 121417
rect 66628 121372 66680 121378
rect 66810 121343 66866 121352
rect 66628 121314 66680 121320
rect 66640 120601 66668 121314
rect 66902 120728 66958 120737
rect 66902 120663 66958 120672
rect 66626 120592 66682 120601
rect 66626 120527 66682 120536
rect 66812 120080 66864 120086
rect 66810 120048 66812 120057
rect 66864 120048 66866 120057
rect 66810 119983 66866 119992
rect 66916 119241 66944 120663
rect 66902 119232 66958 119241
rect 66902 119167 66958 119176
rect 66260 118584 66312 118590
rect 66260 118526 66312 118532
rect 66272 117609 66300 118526
rect 66258 117600 66314 117609
rect 66258 117535 66314 117544
rect 66260 117292 66312 117298
rect 66260 117234 66312 117240
rect 66272 116249 66300 117234
rect 66904 117224 66956 117230
rect 66904 117166 66956 117172
rect 66916 117065 66944 117166
rect 66902 117056 66958 117065
rect 66902 116991 66958 117000
rect 66258 116240 66314 116249
rect 66258 116175 66314 116184
rect 66812 115932 66864 115938
rect 66812 115874 66864 115880
rect 66824 115433 66852 115874
rect 66810 115424 66866 115433
rect 66810 115359 66866 115368
rect 66812 114504 66864 114510
rect 66812 114446 66864 114452
rect 66824 113801 66852 114446
rect 66904 113824 66956 113830
rect 66810 113792 66866 113801
rect 66904 113766 66956 113772
rect 66810 113727 66866 113736
rect 66916 113257 66944 113766
rect 66902 113248 66958 113257
rect 66902 113183 66958 113192
rect 66166 111616 66222 111625
rect 66166 111551 66222 111560
rect 66168 111104 66220 111110
rect 66168 111046 66220 111052
rect 66628 111104 66680 111110
rect 66628 111046 66680 111052
rect 66074 103184 66130 103193
rect 66074 103119 66130 103128
rect 66076 102400 66128 102406
rect 66076 102342 66128 102348
rect 65982 82784 66038 82793
rect 65982 82719 66038 82728
rect 64788 80028 64840 80034
rect 64788 79970 64840 79976
rect 62026 77888 62082 77897
rect 62026 77823 62082 77832
rect 61844 77172 61896 77178
rect 61844 77114 61896 77120
rect 61936 42084 61988 42090
rect 61936 42026 61988 42032
rect 61948 16574 61976 42026
rect 61856 16546 61976 16574
rect 60832 3596 60884 3602
rect 60832 3538 60884 3544
rect 57244 3528 57296 3534
rect 57244 3470 57296 3476
rect 57888 3528 57940 3534
rect 57888 3470 57940 3476
rect 58440 3528 58492 3534
rect 58440 3470 58492 3476
rect 59268 3528 59320 3534
rect 59268 3470 59320 3476
rect 59636 3528 59688 3534
rect 59636 3470 59688 3476
rect 60648 3528 60700 3534
rect 60648 3470 60700 3476
rect 57256 480 57284 3470
rect 58452 480 58480 3470
rect 59648 480 59676 3470
rect 60844 480 60872 3538
rect 61856 3482 61884 16546
rect 62040 6914 62068 77823
rect 66088 75886 66116 102342
rect 66076 75880 66128 75886
rect 66076 75822 66128 75828
rect 66180 74497 66208 111046
rect 66640 110809 66668 111046
rect 66626 110800 66682 110809
rect 66626 110735 66682 110744
rect 66810 110256 66866 110265
rect 66810 110191 66866 110200
rect 66824 109070 66852 110191
rect 66812 109064 66864 109070
rect 66812 109006 66864 109012
rect 66904 108996 66956 109002
rect 66904 108938 66956 108944
rect 66810 108624 66866 108633
rect 66810 108559 66866 108568
rect 66824 107710 66852 108559
rect 66916 107817 66944 108938
rect 66902 107808 66958 107817
rect 66902 107743 66958 107752
rect 66812 107704 66864 107710
rect 66812 107646 66864 107652
rect 66904 107636 66956 107642
rect 66904 107578 66956 107584
rect 66810 106992 66866 107001
rect 66810 106927 66866 106936
rect 66824 106350 66852 106927
rect 66916 106457 66944 107578
rect 66902 106448 66958 106457
rect 66902 106383 66958 106392
rect 66812 106344 66864 106350
rect 66812 106286 66864 106292
rect 66534 105632 66590 105641
rect 66534 105567 66536 105576
rect 66588 105567 66590 105576
rect 66536 105538 66588 105544
rect 66260 104848 66312 104854
rect 66258 104816 66260 104825
rect 66312 104816 66314 104825
rect 66258 104751 66314 104760
rect 66534 102640 66590 102649
rect 66534 102575 66590 102584
rect 66548 102406 66576 102575
rect 66536 102400 66588 102406
rect 66536 102342 66588 102348
rect 66810 101824 66866 101833
rect 66810 101759 66866 101768
rect 66444 101312 66496 101318
rect 66444 101254 66496 101260
rect 66456 101017 66484 101254
rect 66442 101008 66498 101017
rect 66442 100943 66498 100952
rect 66824 100774 66852 101759
rect 66812 100768 66864 100774
rect 66812 100710 66864 100716
rect 66812 100020 66864 100026
rect 66812 99962 66864 99968
rect 66824 99657 66852 99962
rect 66810 99648 66866 99657
rect 66810 99583 66866 99592
rect 66628 99340 66680 99346
rect 66628 99282 66680 99288
rect 66640 98841 66668 99282
rect 66626 98832 66682 98841
rect 66626 98767 66682 98776
rect 67192 98025 67220 247007
rect 67284 129849 67312 280162
rect 67376 247081 67404 309062
rect 67362 247072 67418 247081
rect 67362 247007 67418 247016
rect 67362 246256 67418 246265
rect 67468 246242 67496 396335
rect 67640 390176 67692 390182
rect 67640 390118 67692 390124
rect 67652 267734 67680 390118
rect 67744 325650 67772 397394
rect 67732 325644 67784 325650
rect 67732 325586 67784 325592
rect 67744 324970 67772 325586
rect 67732 324964 67784 324970
rect 67732 324906 67784 324912
rect 68468 318640 68520 318646
rect 68468 318582 68520 318588
rect 68006 280528 68062 280537
rect 68006 280463 68062 280472
rect 67652 267706 67864 267734
rect 67418 246214 67496 246242
rect 67362 246191 67418 246200
rect 67376 220794 67404 246191
rect 67548 244928 67600 244934
rect 67548 244870 67600 244876
rect 67560 244633 67588 244870
rect 67546 244624 67602 244633
rect 67546 244559 67602 244568
rect 67836 242962 67864 267706
rect 67914 257952 67970 257961
rect 67914 257887 67970 257896
rect 67824 242956 67876 242962
rect 67824 242898 67876 242904
rect 67638 233336 67694 233345
rect 67638 233271 67694 233280
rect 67652 233238 67680 233271
rect 67640 233232 67692 233238
rect 67640 233174 67692 233180
rect 67364 220788 67416 220794
rect 67364 220730 67416 220736
rect 67270 129840 67326 129849
rect 67270 129775 67326 129784
rect 67178 98016 67234 98025
rect 67178 97951 67234 97960
rect 66628 97300 66680 97306
rect 66628 97242 66680 97248
rect 66640 96393 66668 97242
rect 66626 96384 66682 96393
rect 66626 96319 66682 96328
rect 67192 89690 67220 97951
rect 67376 97209 67404 220730
rect 67546 147928 67602 147937
rect 67546 147863 67602 147872
rect 67560 147762 67588 147863
rect 67548 147756 67600 147762
rect 67548 147698 67600 147704
rect 67652 112441 67680 233174
rect 67836 203590 67864 242898
rect 67928 238649 67956 257887
rect 67914 238640 67970 238649
rect 67914 238575 67970 238584
rect 68020 229945 68048 280463
rect 68480 248414 68508 318582
rect 68572 284374 68600 431990
rect 68664 287054 68692 432534
rect 112732 432070 112760 433230
rect 112720 432064 112772 432070
rect 112720 432006 112772 432012
rect 113284 431225 113312 447782
rect 113364 442264 113416 442270
rect 113364 442206 113416 442212
rect 113270 431216 113326 431225
rect 113270 431151 113326 431160
rect 113270 427136 113326 427145
rect 113270 427071 113326 427080
rect 113178 420064 113234 420073
rect 113178 419999 113234 420008
rect 112720 407108 112772 407114
rect 112720 407050 112772 407056
rect 112732 405929 112760 407050
rect 112718 405920 112774 405929
rect 112718 405855 112774 405864
rect 87696 390992 87748 390998
rect 108672 390992 108724 390998
rect 87696 390934 87748 390940
rect 102414 390960 102470 390969
rect 84382 390688 84438 390697
rect 84382 390623 84438 390632
rect 80592 390510 80836 390538
rect 72330 390416 72386 390425
rect 68802 390182 68830 390388
rect 69032 390374 69368 390402
rect 69584 390374 70104 390402
rect 68790 390176 68842 390182
rect 68790 390118 68842 390124
rect 69032 292641 69060 390374
rect 69584 373994 69612 390374
rect 70826 390130 70854 390388
rect 69124 373966 69612 373994
rect 70780 390102 70854 390130
rect 71240 390374 71576 390402
rect 71884 390374 72330 390402
rect 69124 318646 69152 373966
rect 70306 364440 70362 364449
rect 70306 364375 70362 364384
rect 69112 318640 69164 318646
rect 69112 318582 69164 318588
rect 70214 317520 70270 317529
rect 70214 317455 70270 317464
rect 69754 317384 69810 317393
rect 69754 317319 69810 317328
rect 69768 316169 69796 317319
rect 69754 316160 69810 316169
rect 69754 316095 69810 316104
rect 69664 295384 69716 295390
rect 69664 295326 69716 295332
rect 69572 294024 69624 294030
rect 69572 293966 69624 293972
rect 69018 292632 69074 292641
rect 69018 292567 69074 292576
rect 68664 287026 68876 287054
rect 68560 284368 68612 284374
rect 68560 284310 68612 284316
rect 68572 279721 68600 284310
rect 68848 283626 68876 287026
rect 69110 285832 69166 285841
rect 69110 285767 69166 285776
rect 68836 283620 68888 283626
rect 68836 283562 68888 283568
rect 68848 281217 68876 283562
rect 69124 283370 69152 285767
rect 69202 285696 69258 285705
rect 69202 285631 69258 285640
rect 69216 283665 69244 285631
rect 69480 284980 69532 284986
rect 69480 284922 69532 284928
rect 69492 283778 69520 284922
rect 69584 284866 69612 293966
rect 69676 284986 69704 295326
rect 69768 285841 69796 316095
rect 70228 294030 70256 317455
rect 70320 317393 70348 364375
rect 70306 317384 70362 317393
rect 70306 317319 70362 317328
rect 70216 294024 70268 294030
rect 70216 293966 70268 293972
rect 69754 285832 69810 285841
rect 69754 285767 69810 285776
rect 69664 284980 69716 284986
rect 69664 284922 69716 284928
rect 69584 284838 69888 284866
rect 69492 283750 69704 283778
rect 69202 283656 69258 283665
rect 69202 283591 69258 283600
rect 69000 283342 69152 283370
rect 69216 283370 69244 283591
rect 69216 283342 69552 283370
rect 69676 283014 69704 283750
rect 69860 283506 69888 284838
rect 70780 283665 70808 390102
rect 71240 387841 71268 390374
rect 71778 389056 71834 389065
rect 71778 388991 71834 389000
rect 71688 387864 71740 387870
rect 71226 387832 71282 387841
rect 71688 387806 71740 387812
rect 71226 387767 71282 387776
rect 71042 298752 71098 298761
rect 71042 298687 71098 298696
rect 71056 288386 71084 298687
rect 71700 292670 71728 387806
rect 71792 381546 71820 388991
rect 71884 388929 71912 390374
rect 73986 390416 74042 390425
rect 72330 390351 72386 390360
rect 72528 390374 72864 390402
rect 73264 390374 73600 390402
rect 72528 389065 72556 390374
rect 72514 389056 72570 389065
rect 72514 388991 72570 389000
rect 71870 388920 71926 388929
rect 71870 388855 71926 388864
rect 73264 387870 73292 390374
rect 77206 390416 77262 390425
rect 74042 390374 74336 390402
rect 74552 390374 75072 390402
rect 75288 390374 75624 390402
rect 75932 390374 76360 390402
rect 76760 390374 77206 390402
rect 73986 390351 74042 390360
rect 73252 387864 73304 387870
rect 73252 387806 73304 387812
rect 73158 387696 73214 387705
rect 73158 387631 73214 387640
rect 72424 386368 72476 386374
rect 72424 386310 72476 386316
rect 71780 381540 71832 381546
rect 71780 381482 71832 381488
rect 72436 313313 72464 386310
rect 73066 380216 73122 380225
rect 73066 380151 73122 380160
rect 72422 313304 72478 313313
rect 72422 313239 72478 313248
rect 71870 299568 71926 299577
rect 71870 299503 71926 299512
rect 71688 292664 71740 292670
rect 71688 292606 71740 292612
rect 71044 288380 71096 288386
rect 71044 288322 71096 288328
rect 70766 283656 70822 283665
rect 70766 283591 70822 283600
rect 71056 283506 71084 288322
rect 71780 286340 71832 286346
rect 71780 286282 71832 286288
rect 71318 286104 71374 286113
rect 71318 286039 71374 286048
rect 69860 283478 70104 283506
rect 70656 283478 71084 283506
rect 71332 283370 71360 286039
rect 71792 283778 71820 286282
rect 71746 283750 71820 283778
rect 71746 283492 71774 283750
rect 71884 283506 71912 299503
rect 71964 292664 72016 292670
rect 71964 292606 72016 292612
rect 71976 284209 72004 292606
rect 72436 284442 72464 313239
rect 73080 299577 73108 380151
rect 73066 299568 73122 299577
rect 73066 299503 73122 299512
rect 72424 284436 72476 284442
rect 72424 284378 72476 284384
rect 71962 284200 72018 284209
rect 71962 284135 72018 284144
rect 72436 283506 72464 284378
rect 73172 283529 73200 387631
rect 74000 387122 74028 390351
rect 73988 387116 74040 387122
rect 73988 387058 74040 387064
rect 74552 366382 74580 390374
rect 75288 387569 75316 390374
rect 75274 387560 75330 387569
rect 75274 387495 75330 387504
rect 75184 386368 75236 386374
rect 75184 386310 75236 386316
rect 74540 366376 74592 366382
rect 74540 366318 74592 366324
rect 75196 320890 75224 386310
rect 75932 369170 75960 390374
rect 76760 389065 76788 390374
rect 79414 390416 79470 390425
rect 77206 390351 77262 390360
rect 77496 390374 77832 390402
rect 77956 390374 78384 390402
rect 78876 390374 79414 390402
rect 76010 389056 76066 389065
rect 76010 388991 76066 389000
rect 76746 389056 76802 389065
rect 76746 388991 76802 389000
rect 76024 374678 76052 388991
rect 77298 387968 77354 387977
rect 77298 387903 77354 387912
rect 77312 387682 77340 387903
rect 77128 387654 77340 387682
rect 76012 374672 76064 374678
rect 76012 374614 76064 374620
rect 75920 369164 75972 369170
rect 75920 369106 75972 369112
rect 75274 327040 75330 327049
rect 75274 326975 75330 326984
rect 75184 320884 75236 320890
rect 75184 320826 75236 320832
rect 74540 316940 74592 316946
rect 74540 316882 74592 316888
rect 73526 304192 73582 304201
rect 73526 304127 73582 304136
rect 73158 283520 73214 283529
rect 71884 283478 72312 283506
rect 72436 283478 72864 283506
rect 73540 283506 73568 304127
rect 74552 283778 74580 316882
rect 75288 285977 75316 326975
rect 77022 318744 77078 318753
rect 77022 318679 77078 318688
rect 76470 291272 76526 291281
rect 76470 291207 76526 291216
rect 75274 285968 75330 285977
rect 75274 285903 75330 285912
rect 74506 283750 74580 283778
rect 73214 283478 73416 283506
rect 73540 283478 73968 283506
rect 73158 283455 73214 283464
rect 73172 283395 73200 283455
rect 70964 283342 71360 283370
rect 69664 283008 69716 283014
rect 70964 282985 70992 283342
rect 74354 283248 74410 283257
rect 74506 283234 74534 283750
rect 75288 283506 75316 285903
rect 76484 283506 76512 291207
rect 77036 286346 77064 318679
rect 77128 314945 77156 387654
rect 77496 385801 77524 390374
rect 77482 385792 77538 385801
rect 77482 385727 77538 385736
rect 77956 373994 77984 390374
rect 78876 389065 78904 390374
rect 79856 390374 80008 390402
rect 79414 390351 79470 390360
rect 78862 389056 78918 389065
rect 78862 388991 78918 389000
rect 79980 387870 80008 390374
rect 80058 389056 80114 389065
rect 80058 388991 80114 389000
rect 79968 387864 80020 387870
rect 79968 387806 80020 387812
rect 79874 383752 79930 383761
rect 79874 383687 79930 383696
rect 79322 378720 79378 378729
rect 79322 378655 79378 378664
rect 77312 373966 77984 373994
rect 77206 365664 77262 365673
rect 77206 365599 77262 365608
rect 77114 314936 77170 314945
rect 77114 314871 77170 314880
rect 77128 291281 77156 314871
rect 77114 291272 77170 291281
rect 77114 291207 77170 291216
rect 77220 289921 77248 365599
rect 77312 360874 77340 373966
rect 77300 360868 77352 360874
rect 77300 360810 77352 360816
rect 78496 322788 78548 322794
rect 78496 322730 78548 322736
rect 78508 302258 78536 322730
rect 78586 318336 78642 318345
rect 78586 318271 78642 318280
rect 77300 302252 77352 302258
rect 77300 302194 77352 302200
rect 78496 302252 78548 302258
rect 78496 302194 78548 302200
rect 77206 289912 77262 289921
rect 77206 289847 77262 289856
rect 77220 288538 77248 289847
rect 77128 288510 77248 288538
rect 77024 286340 77076 286346
rect 77024 286282 77076 286288
rect 77128 283506 77156 288510
rect 77312 283778 77340 302194
rect 78600 288454 78628 318271
rect 79336 288522 79364 378655
rect 79414 323640 79470 323649
rect 79414 323575 79470 323584
rect 79324 288516 79376 288522
rect 79324 288458 79376 288464
rect 78588 288448 78640 288454
rect 78588 288390 78640 288396
rect 78126 286240 78182 286249
rect 78126 286175 78182 286184
rect 75072 283478 75316 283506
rect 76176 283478 76512 283506
rect 76728 283478 77156 283506
rect 77266 283750 77340 283778
rect 77266 283492 77294 283750
rect 78140 283506 78168 286175
rect 78600 283506 78628 288390
rect 79428 287094 79456 323575
rect 79888 318073 79916 383687
rect 79968 379568 80020 379574
rect 79968 379510 80020 379516
rect 79874 318064 79930 318073
rect 79874 317999 79930 318008
rect 79888 316034 79916 317999
rect 79520 316006 79916 316034
rect 79416 287088 79468 287094
rect 79416 287030 79468 287036
rect 79428 283778 79456 287030
rect 79520 286249 79548 316006
rect 79980 301510 80008 379510
rect 80072 378826 80100 388991
rect 80704 387864 80756 387870
rect 80704 387806 80756 387812
rect 80060 378820 80112 378826
rect 80060 378762 80112 378768
rect 80716 369170 80744 387806
rect 80808 386306 80836 390510
rect 81990 390416 82046 390425
rect 80992 390374 81328 390402
rect 81452 390374 81990 390402
rect 80992 389065 81020 390374
rect 80978 389056 81034 389065
rect 80978 388991 81034 389000
rect 81452 388793 81480 390374
rect 81990 390351 82046 390360
rect 82280 390374 82616 390402
rect 83016 390374 83352 390402
rect 81438 388784 81494 388793
rect 81438 388719 81494 388728
rect 80796 386300 80848 386306
rect 80796 386242 80848 386248
rect 81256 386300 81308 386306
rect 81256 386242 81308 386248
rect 81268 385665 81296 386242
rect 81254 385656 81310 385665
rect 81254 385591 81310 385600
rect 81452 379574 81480 388719
rect 82280 386374 82308 390374
rect 83016 389162 83044 390374
rect 84074 390130 84102 390388
rect 84074 390102 84148 390130
rect 83004 389156 83056 389162
rect 83004 389098 83056 389104
rect 84120 388482 84148 390102
rect 84108 388476 84160 388482
rect 84108 388418 84160 388424
rect 84200 387048 84252 387054
rect 84200 386990 84252 386996
rect 82268 386368 82320 386374
rect 82268 386310 82320 386316
rect 84212 381546 84240 386990
rect 84200 381540 84252 381546
rect 84200 381482 84252 381488
rect 81440 379568 81492 379574
rect 81440 379510 81492 379516
rect 84106 376000 84162 376009
rect 84106 375935 84162 375944
rect 80704 369164 80756 369170
rect 80704 369106 80756 369112
rect 83554 339552 83610 339561
rect 83554 339487 83556 339496
rect 83608 339487 83610 339496
rect 83556 339458 83608 339464
rect 84014 330440 84070 330449
rect 84014 330375 84070 330384
rect 81440 327752 81492 327758
rect 81440 327694 81492 327700
rect 80702 320784 80758 320793
rect 80702 320719 80758 320728
rect 80716 306374 80744 320719
rect 81346 319424 81402 319433
rect 81346 319359 81402 319368
rect 80716 306346 80836 306374
rect 79968 301504 80020 301510
rect 79968 301446 80020 301452
rect 79600 288516 79652 288522
rect 79600 288458 79652 288464
rect 79506 286240 79562 286249
rect 79506 286175 79562 286184
rect 79336 283750 79456 283778
rect 79336 283506 79364 283750
rect 79612 283506 79640 288458
rect 80334 288416 80390 288425
rect 80334 288351 80390 288360
rect 80348 287201 80376 288351
rect 80334 287192 80390 287201
rect 80334 287127 80390 287136
rect 80348 283506 80376 287127
rect 80808 285734 80836 306346
rect 81254 303648 81310 303657
rect 81254 303583 81310 303592
rect 80796 285728 80848 285734
rect 80796 285670 80848 285676
rect 77832 283478 78168 283506
rect 78384 283478 78628 283506
rect 78936 283478 79364 283506
rect 79488 283478 79640 283506
rect 80040 283478 80376 283506
rect 80808 283506 80836 285670
rect 80808 283478 81144 283506
rect 75734 283248 75790 283257
rect 74410 283220 74534 283234
rect 74410 283206 74520 283220
rect 75624 283206 75734 283234
rect 74354 283183 74410 283192
rect 75734 283183 75790 283192
rect 81268 282985 81296 303583
rect 81360 288425 81388 319359
rect 81346 288416 81402 288425
rect 81346 288351 81402 288360
rect 81452 283014 81480 327694
rect 81530 318200 81586 318209
rect 81530 318135 81586 318144
rect 81544 316946 81572 318135
rect 81532 316940 81584 316946
rect 81532 316882 81584 316888
rect 82912 316736 82964 316742
rect 82912 316678 82964 316684
rect 82820 296744 82872 296750
rect 82820 296686 82872 296692
rect 82728 289128 82780 289134
rect 82726 289096 82728 289105
rect 82780 289096 82782 289105
rect 82726 289031 82782 289040
rect 82450 285696 82506 285705
rect 82450 285631 82506 285640
rect 82464 283506 82492 285631
rect 82832 283778 82860 296686
rect 82924 284986 82952 316678
rect 84028 296750 84056 330375
rect 84016 296744 84068 296750
rect 84016 296686 84068 296692
rect 84120 289950 84148 375935
rect 84396 322794 84424 390623
rect 87708 390402 87736 390934
rect 93676 390924 93728 390930
rect 102414 390895 102470 390904
rect 106738 390960 106794 390969
rect 106794 390918 107516 390946
rect 108376 390940 108672 390946
rect 108376 390934 108724 390940
rect 108376 390918 108712 390934
rect 106738 390895 106794 390904
rect 93676 390866 93728 390872
rect 93688 390810 93716 390866
rect 93688 390796 93840 390810
rect 93688 390782 93854 390796
rect 84824 390374 84976 390402
rect 84948 387870 84976 390374
rect 85040 390374 85376 390402
rect 85592 390374 86112 390402
rect 84936 387864 84988 387870
rect 84936 387806 84988 387812
rect 85040 387054 85068 390374
rect 85028 387048 85080 387054
rect 85028 386990 85080 386996
rect 85592 367810 85620 390374
rect 86834 390130 86862 390388
rect 86972 390374 87584 390402
rect 87708 390374 88136 390402
rect 88444 390374 88872 390402
rect 89272 390374 89608 390402
rect 89732 390374 90344 390402
rect 91080 390374 91232 390402
rect 86834 390102 86908 390130
rect 86224 387864 86276 387870
rect 86224 387806 86276 387812
rect 85580 367804 85632 367810
rect 85580 367746 85632 367752
rect 86236 363662 86264 387806
rect 86880 387122 86908 390102
rect 86868 387116 86920 387122
rect 86868 387058 86920 387064
rect 86866 380216 86922 380225
rect 86866 380151 86922 380160
rect 86776 374672 86828 374678
rect 86776 374614 86828 374620
rect 86224 363656 86276 363662
rect 86224 363598 86276 363604
rect 85396 327072 85448 327078
rect 85396 327014 85448 327020
rect 84384 322788 84436 322794
rect 84384 322730 84436 322736
rect 84198 294672 84254 294681
rect 84198 294607 84254 294616
rect 83004 289944 83056 289950
rect 83004 289886 83056 289892
rect 84108 289944 84160 289950
rect 84108 289886 84160 289892
rect 82912 284980 82964 284986
rect 82912 284922 82964 284928
rect 82248 283478 82492 283506
rect 82786 283750 82860 283778
rect 82786 283492 82814 283750
rect 83016 283506 83044 289886
rect 83556 284980 83608 284986
rect 83556 284922 83608 284928
rect 83568 283506 83596 284922
rect 84212 283506 84240 294607
rect 84568 293276 84620 293282
rect 84568 293218 84620 293224
rect 84580 283506 84608 293218
rect 85408 283665 85436 327014
rect 85580 304292 85632 304298
rect 85580 304234 85632 304240
rect 85592 283778 85620 304234
rect 86788 288561 86816 374614
rect 86774 288552 86830 288561
rect 86774 288487 86830 288496
rect 86788 287054 86816 288487
rect 85546 283750 85620 283778
rect 86512 287026 86816 287054
rect 85394 283656 85450 283665
rect 85394 283591 85450 283600
rect 83016 283478 83352 283506
rect 83568 283478 83904 283506
rect 84212 283478 84456 283506
rect 84580 283478 85008 283506
rect 85546 283492 85574 283750
rect 86512 283506 86540 287026
rect 86880 284442 86908 380151
rect 86972 293185 87000 390374
rect 87708 377534 87736 390374
rect 88338 389056 88394 389065
rect 88338 388991 88394 389000
rect 88248 379500 88300 379506
rect 88248 379442 88300 379448
rect 87696 377528 87748 377534
rect 87696 377470 87748 377476
rect 88260 335850 88288 379442
rect 87604 335844 87656 335850
rect 87604 335786 87656 335792
rect 88248 335844 88300 335850
rect 88248 335786 88300 335792
rect 87050 316704 87106 316713
rect 87050 316639 87106 316648
rect 86958 293176 87014 293185
rect 86958 293111 87014 293120
rect 86868 284436 86920 284442
rect 86868 284378 86920 284384
rect 86880 283506 86908 284378
rect 86112 283478 86540 283506
rect 86664 283478 86908 283506
rect 87064 283506 87092 316639
rect 87616 293350 87644 335786
rect 88260 335374 88288 335786
rect 88248 335368 88300 335374
rect 88248 335310 88300 335316
rect 88352 327078 88380 388991
rect 88444 383654 88472 390374
rect 89272 389065 89300 390374
rect 89258 389056 89314 389065
rect 89258 388991 89314 389000
rect 89626 385656 89682 385665
rect 89626 385591 89682 385600
rect 88432 383648 88484 383654
rect 88432 383590 88484 383596
rect 88340 327072 88392 327078
rect 88340 327014 88392 327020
rect 89534 326360 89590 326369
rect 89534 326295 89590 326304
rect 89444 322924 89496 322930
rect 89444 322866 89496 322872
rect 88246 319560 88302 319569
rect 88246 319495 88302 319504
rect 87604 293344 87656 293350
rect 87604 293286 87656 293292
rect 88260 287054 88288 319495
rect 89456 312497 89484 322866
rect 89442 312488 89498 312497
rect 89442 312423 89498 312432
rect 89548 296714 89576 326295
rect 89272 296686 89576 296714
rect 89272 287337 89300 296686
rect 89534 288416 89590 288425
rect 89534 288351 89590 288360
rect 89258 287328 89314 287337
rect 89258 287263 89314 287272
rect 88168 287026 88288 287054
rect 87064 283478 87216 283506
rect 81440 283008 81492 283014
rect 69664 282950 69716 282956
rect 70950 282976 71006 282985
rect 80886 282976 80942 282985
rect 80592 282934 80886 282962
rect 70950 282911 71006 282920
rect 80886 282911 80942 282920
rect 81254 282976 81310 282985
rect 87878 282976 87934 282985
rect 81492 282956 81696 282962
rect 81440 282950 81696 282956
rect 81452 282934 81696 282950
rect 87768 282934 87878 282962
rect 81254 282911 81310 282920
rect 88168 282962 88196 287026
rect 89272 283506 89300 287263
rect 88872 283478 89300 283506
rect 88522 282976 88578 282985
rect 87934 282934 88196 282962
rect 88320 282934 88522 282962
rect 87878 282911 87934 282920
rect 89548 282962 89576 288351
rect 89640 285705 89668 385591
rect 89732 300801 89760 390374
rect 90364 387864 90416 387870
rect 90364 387806 90416 387812
rect 90376 322969 90404 387806
rect 91204 384402 91232 390374
rect 91388 390374 91632 390402
rect 91756 390374 92368 390402
rect 92492 390374 93104 390402
rect 91388 387870 91416 390374
rect 91376 387864 91428 387870
rect 91282 387832 91338 387841
rect 91376 387806 91428 387812
rect 91282 387767 91338 387776
rect 91192 384396 91244 384402
rect 91192 384338 91244 384344
rect 91006 373280 91062 373289
rect 91006 373215 91062 373224
rect 90362 322960 90418 322969
rect 90362 322895 90418 322904
rect 89812 320884 89864 320890
rect 89812 320826 89864 320832
rect 89824 306374 89852 320826
rect 89824 306346 90128 306374
rect 89718 300792 89774 300801
rect 89718 300727 89774 300736
rect 89626 285696 89682 285705
rect 89626 285631 89682 285640
rect 89950 283756 90002 283762
rect 89950 283698 90002 283704
rect 89810 283520 89866 283529
rect 89962 283506 89990 283698
rect 89866 283492 89990 283506
rect 90100 283506 90128 306346
rect 91020 283762 91048 373215
rect 91296 327758 91324 387767
rect 91756 383625 91784 390374
rect 92386 387016 92442 387025
rect 92386 386951 92442 386960
rect 91374 383616 91430 383625
rect 91374 383551 91430 383560
rect 91742 383616 91798 383625
rect 91742 383551 91798 383560
rect 91388 379506 91416 383551
rect 91376 379500 91428 379506
rect 91376 379442 91428 379448
rect 92296 378140 92348 378146
rect 92296 378082 92348 378088
rect 92308 377466 92336 378082
rect 92296 377460 92348 377466
rect 92296 377402 92348 377408
rect 91284 327752 91336 327758
rect 91284 327694 91336 327700
rect 92204 320952 92256 320958
rect 92204 320894 92256 320900
rect 92216 292574 92244 320894
rect 92308 308417 92336 377402
rect 92294 308408 92350 308417
rect 92294 308343 92350 308352
rect 92400 292574 92428 386951
rect 92492 385014 92520 390374
rect 93826 390130 93854 390782
rect 94378 390130 94406 390388
rect 94516 390374 95128 390402
rect 95252 390374 95864 390402
rect 93826 390102 93900 390130
rect 94378 390102 94452 390130
rect 93124 387864 93176 387870
rect 93124 387806 93176 387812
rect 92480 385008 92532 385014
rect 92480 384950 92532 384956
rect 92492 351937 92520 384950
rect 93136 378146 93164 387806
rect 93766 384296 93822 384305
rect 93766 384231 93822 384240
rect 93124 378140 93176 378146
rect 93124 378082 93176 378088
rect 93674 353968 93730 353977
rect 93674 353903 93730 353912
rect 92478 351928 92534 351937
rect 92478 351863 92534 351872
rect 93688 336802 93716 353903
rect 93124 336796 93176 336802
rect 93124 336738 93176 336744
rect 93676 336796 93728 336802
rect 93676 336738 93728 336744
rect 93030 293312 93086 293321
rect 93030 293247 93032 293256
rect 93084 293247 93086 293256
rect 93032 293218 93084 293224
rect 92032 292546 92244 292574
rect 92308 292546 92428 292574
rect 91468 291236 91520 291242
rect 91468 291178 91520 291184
rect 91374 285560 91430 285569
rect 91374 285495 91430 285504
rect 91388 284481 91416 285495
rect 91374 284472 91430 284481
rect 91374 284407 91430 284416
rect 91008 283756 91060 283762
rect 91008 283698 91060 283704
rect 91388 283506 91416 284407
rect 91480 284209 91508 291178
rect 91466 284200 91522 284209
rect 91466 284135 91522 284144
rect 92032 283506 92060 292546
rect 92308 285569 92336 292546
rect 93136 287026 93164 336738
rect 93676 331220 93728 331226
rect 93676 331162 93728 331168
rect 92388 287020 92440 287026
rect 92388 286962 92440 286968
rect 93124 287020 93176 287026
rect 93124 286962 93176 286968
rect 92294 285560 92350 285569
rect 92294 285495 92350 285504
rect 92400 283506 92428 286962
rect 93688 286113 93716 331162
rect 93780 287473 93808 384231
rect 93872 322930 93900 390102
rect 94424 387841 94452 390102
rect 94410 387832 94466 387841
rect 94410 387767 94466 387776
rect 94042 382256 94098 382265
rect 94042 382191 94098 382200
rect 94056 331226 94084 382191
rect 94516 380186 94544 390374
rect 94596 389496 94648 389502
rect 94596 389438 94648 389444
rect 94608 389366 94636 389438
rect 94596 389360 94648 389366
rect 94596 389302 94648 389308
rect 94504 380180 94556 380186
rect 94504 380122 94556 380128
rect 94044 331220 94096 331226
rect 94044 331162 94096 331168
rect 93860 322924 93912 322930
rect 93860 322866 93912 322872
rect 95252 321473 95280 390374
rect 96586 390130 96614 390388
rect 97000 390374 97336 390402
rect 97460 390374 97888 390402
rect 98288 390374 98624 390402
rect 99360 390374 99696 390402
rect 100096 390374 100432 390402
rect 96586 390102 96660 390130
rect 95330 389600 95386 389609
rect 95330 389535 95386 389544
rect 95344 374678 95372 389535
rect 96632 387802 96660 390102
rect 97000 387870 97028 390374
rect 97460 389722 97488 390374
rect 97184 389694 97488 389722
rect 96988 387864 97040 387870
rect 96988 387806 97040 387812
rect 96620 387796 96672 387802
rect 96620 387738 96672 387744
rect 96632 386442 96660 387738
rect 96620 386436 96672 386442
rect 96620 386378 96672 386384
rect 97184 376009 97212 389694
rect 98288 389366 98316 390374
rect 98276 389360 98328 389366
rect 98276 389302 98328 389308
rect 97264 389156 97316 389162
rect 97264 389098 97316 389104
rect 97170 376000 97226 376009
rect 97170 375935 97226 375944
rect 95332 374672 95384 374678
rect 95332 374614 95384 374620
rect 96526 374640 96582 374649
rect 96526 374575 96582 374584
rect 95238 321464 95294 321473
rect 95238 321399 95294 321408
rect 95884 317484 95936 317490
rect 95884 317426 95936 317432
rect 95896 304298 95924 317426
rect 95884 304292 95936 304298
rect 95884 304234 95936 304240
rect 96436 304292 96488 304298
rect 96436 304234 96488 304240
rect 94504 289876 94556 289882
rect 94504 289818 94556 289824
rect 94516 289134 94544 289818
rect 94504 289128 94556 289134
rect 94504 289070 94556 289076
rect 96448 288522 96476 304234
rect 95608 288516 95660 288522
rect 95608 288458 95660 288464
rect 96436 288516 96488 288522
rect 96436 288458 96488 288464
rect 93766 287464 93822 287473
rect 93766 287399 93822 287408
rect 93030 286104 93086 286113
rect 93030 286039 93086 286048
rect 93674 286104 93730 286113
rect 93674 286039 93730 286048
rect 89866 283478 89976 283492
rect 90100 283478 90528 283506
rect 91080 283478 91416 283506
rect 91632 283478 92060 283506
rect 92184 283478 92428 283506
rect 92570 283520 92626 283529
rect 89810 283455 89866 283464
rect 93044 283506 93072 286039
rect 93780 283778 93808 287399
rect 95148 287156 95200 287162
rect 95148 287098 95200 287104
rect 94688 287020 94740 287026
rect 94688 286962 94740 286968
rect 94134 286376 94190 286385
rect 94134 286311 94190 286320
rect 93688 283750 93808 283778
rect 93688 283506 93716 283750
rect 94148 283506 94176 286311
rect 94700 283506 94728 286962
rect 95160 283506 95188 287098
rect 95620 283506 95648 288458
rect 96540 287094 96568 374575
rect 96710 330304 96766 330313
rect 96710 330239 96766 330248
rect 96620 314696 96672 314702
rect 96620 314638 96672 314644
rect 96528 287088 96580 287094
rect 96528 287030 96580 287036
rect 96020 283792 96076 283801
rect 96632 283778 96660 314638
rect 96020 283727 96076 283736
rect 96586 283750 96660 283778
rect 92626 283478 93072 283506
rect 93288 283478 93716 283506
rect 93840 283478 94176 283506
rect 94392 283478 94728 283506
rect 94944 283478 95188 283506
rect 95496 283478 95648 283506
rect 96034 283492 96062 283727
rect 96586 283492 96614 283750
rect 96724 283506 96752 330239
rect 97276 291242 97304 389098
rect 99668 389065 99696 390374
rect 100298 390280 100354 390289
rect 100298 390215 100354 390224
rect 99654 389056 99710 389065
rect 99654 388991 99710 389000
rect 97356 386436 97408 386442
rect 97356 386378 97408 386384
rect 97368 345014 97396 386378
rect 100312 383654 100340 390215
rect 100404 386306 100432 390374
rect 100818 390130 100846 390388
rect 101384 390374 101720 390402
rect 102120 390374 102272 390402
rect 100772 390102 100846 390130
rect 100772 389434 100800 390102
rect 100760 389428 100812 389434
rect 100760 389370 100812 389376
rect 100772 389065 100800 389370
rect 101692 389230 101720 390374
rect 102048 389836 102100 389842
rect 102048 389778 102100 389784
rect 101680 389224 101732 389230
rect 101680 389166 101732 389172
rect 100482 389056 100538 389065
rect 100482 388991 100538 389000
rect 100758 389056 100814 389065
rect 100758 388991 100814 389000
rect 100392 386300 100444 386306
rect 100392 386242 100444 386248
rect 100312 383626 100432 383654
rect 97816 378276 97868 378282
rect 97816 378218 97868 378224
rect 97368 344986 97764 345014
rect 97736 342310 97764 344986
rect 97724 342304 97776 342310
rect 97724 342246 97776 342252
rect 97736 309806 97764 342246
rect 97828 330313 97856 378218
rect 97906 376000 97962 376009
rect 97906 375935 97962 375944
rect 97814 330304 97870 330313
rect 97814 330239 97870 330248
rect 97828 329905 97856 330239
rect 97814 329896 97870 329905
rect 97814 329831 97870 329840
rect 97920 315314 97948 375935
rect 100024 334008 100076 334014
rect 100024 333950 100076 333956
rect 99288 332648 99340 332654
rect 99286 332616 99288 332625
rect 99340 332616 99342 332625
rect 99286 332551 99342 332560
rect 98090 327720 98146 327729
rect 98090 327655 98146 327664
rect 97908 315308 97960 315314
rect 97908 315250 97960 315256
rect 97920 314702 97948 315250
rect 97908 314696 97960 314702
rect 97908 314638 97960 314644
rect 97724 309800 97776 309806
rect 97724 309742 97776 309748
rect 97264 291236 97316 291242
rect 97264 291178 97316 291184
rect 97998 287464 98054 287473
rect 97998 287399 98054 287408
rect 96724 283478 97152 283506
rect 92570 283455 92626 283464
rect 89628 283008 89680 283014
rect 89424 282956 89628 282962
rect 97906 282976 97962 282985
rect 89424 282950 89680 282956
rect 89424 282934 89668 282950
rect 97704 282934 97906 282962
rect 88522 282911 88578 282920
rect 97906 282911 97962 282920
rect 69020 282736 69072 282742
rect 69018 282704 69020 282713
rect 69072 282704 69074 282713
rect 69018 282639 69074 282648
rect 98012 282266 98040 287399
rect 98104 282826 98132 327655
rect 98368 319524 98420 319530
rect 98368 319466 98420 319472
rect 98104 282812 98256 282826
rect 98104 282798 98270 282812
rect 98242 282554 98270 282798
rect 98242 282526 98316 282554
rect 98000 282260 98052 282266
rect 98000 282202 98052 282208
rect 68834 281208 68890 281217
rect 68834 281143 68890 281152
rect 68848 280226 68876 281143
rect 68836 280220 68888 280226
rect 68836 280162 68888 280168
rect 68558 279712 68614 279721
rect 68558 279647 68614 279656
rect 98182 270736 98238 270745
rect 98182 270671 98238 270680
rect 68480 248386 68968 248414
rect 68468 242956 68520 242962
rect 68468 242898 68520 242904
rect 68480 242298 68508 242898
rect 68480 242270 68816 242298
rect 68940 241482 68968 248386
rect 98090 247072 98146 247081
rect 98090 247007 98146 247016
rect 69018 244352 69074 244361
rect 69018 244287 69074 244296
rect 69032 243574 69060 244287
rect 69020 243568 69072 243574
rect 69020 243510 69072 243516
rect 96896 241800 96948 241806
rect 69478 241768 69534 241777
rect 69184 241726 69478 241754
rect 70950 241768 71006 241777
rect 69478 241703 69534 241712
rect 70412 241726 70950 241754
rect 70030 241632 70086 241641
rect 69308 241590 69736 241618
rect 69860 241590 70030 241618
rect 69308 241482 69336 241590
rect 69860 241482 69888 241590
rect 70086 241590 70288 241618
rect 70030 241567 70086 241576
rect 68940 241454 69336 241482
rect 69492 241454 69888 241482
rect 69940 241528 69992 241534
rect 69940 241470 69992 241476
rect 68006 229936 68062 229945
rect 68006 229871 68062 229880
rect 67824 203584 67876 203590
rect 67824 203526 67876 203532
rect 67732 149728 67784 149734
rect 67732 149670 67784 149676
rect 67744 133657 67772 149670
rect 69032 142154 69060 241454
rect 69492 229770 69520 241454
rect 69952 238754 69980 241470
rect 69664 238740 69716 238746
rect 69664 238682 69716 238688
rect 69860 238726 69980 238754
rect 69480 229764 69532 229770
rect 69480 229706 69532 229712
rect 69676 208457 69704 238682
rect 69860 238066 69888 238726
rect 69848 238060 69900 238066
rect 69848 238002 69900 238008
rect 69662 208448 69718 208457
rect 69662 208383 69718 208392
rect 69664 142860 69716 142866
rect 69664 142802 69716 142808
rect 68664 142126 69060 142154
rect 67824 139460 67876 139466
rect 67824 139402 67876 139408
rect 67730 133648 67786 133657
rect 67730 133583 67786 133592
rect 67730 129024 67786 129033
rect 67730 128959 67786 128968
rect 67638 112432 67694 112441
rect 67638 112367 67694 112376
rect 67362 97200 67418 97209
rect 67362 97135 67418 97144
rect 67376 92478 67404 97135
rect 67454 95840 67510 95849
rect 67454 95775 67510 95784
rect 67364 92472 67416 92478
rect 67364 92414 67416 92420
rect 67180 89684 67232 89690
rect 67180 89626 67232 89632
rect 67468 85474 67496 95775
rect 67546 94208 67602 94217
rect 67546 94143 67602 94152
rect 67560 92410 67588 94143
rect 67548 92404 67600 92410
rect 67548 92346 67600 92352
rect 67548 90364 67600 90370
rect 67548 90306 67600 90312
rect 67456 85468 67508 85474
rect 67456 85410 67508 85416
rect 66166 74488 66222 74497
rect 66166 74423 66222 74432
rect 67560 66910 67588 90306
rect 67548 66904 67600 66910
rect 67548 66846 67600 66852
rect 66168 36576 66220 36582
rect 66168 36518 66220 36524
rect 64786 10296 64842 10305
rect 64786 10231 64842 10240
rect 61948 6886 62068 6914
rect 61948 3602 61976 6886
rect 63222 4040 63278 4049
rect 63222 3975 63278 3984
rect 61936 3596 61988 3602
rect 61936 3538 61988 3544
rect 61856 3454 62068 3482
rect 62040 480 62068 3454
rect 63236 480 63264 3975
rect 64800 3534 64828 10231
rect 66180 3534 66208 36518
rect 67744 33794 67772 128959
rect 67836 128217 67864 139402
rect 67822 128208 67878 128217
rect 67822 128143 67878 128152
rect 68664 113174 68692 142126
rect 69294 138000 69350 138009
rect 69294 137935 69350 137944
rect 69308 134722 69336 137935
rect 69388 137828 69440 137834
rect 69388 137770 69440 137776
rect 69000 134694 69336 134722
rect 68836 134632 68888 134638
rect 68836 134574 68888 134580
rect 69400 134586 69428 137770
rect 69572 135924 69624 135930
rect 69572 135866 69624 135872
rect 69584 135017 69612 135866
rect 69570 135008 69626 135017
rect 69570 134943 69626 134952
rect 69676 134722 69704 142802
rect 70308 141432 70360 141438
rect 70306 141400 70308 141409
rect 70360 141400 70362 141409
rect 70306 141335 70362 141344
rect 70412 140078 70440 241726
rect 70950 241703 71006 241712
rect 72330 241768 72386 241777
rect 73894 241768 73950 241777
rect 72386 241726 72832 241754
rect 72330 241703 72386 241712
rect 70964 241670 70992 241703
rect 70952 241664 71004 241670
rect 70952 241606 71004 241612
rect 71056 241590 71544 241618
rect 71056 241369 71084 241590
rect 71042 241360 71098 241369
rect 71042 241295 71098 241304
rect 71516 240825 71544 241590
rect 71792 241590 71944 241618
rect 71502 240816 71558 240825
rect 71502 240751 71558 240760
rect 71792 240038 71820 241590
rect 71780 240032 71832 240038
rect 71780 239974 71832 239980
rect 72516 240032 72568 240038
rect 72516 239974 72568 239980
rect 72424 238128 72476 238134
rect 72424 238070 72476 238076
rect 72436 161673 72464 238070
rect 72528 229770 72556 239974
rect 72804 238754 72832 241726
rect 83370 241768 83426 241777
rect 73950 241740 74152 241754
rect 73950 241726 74166 241740
rect 73894 241703 73950 241712
rect 74138 241618 74166 241726
rect 84934 241768 84990 241777
rect 83426 241726 83536 241754
rect 83370 241703 83426 241712
rect 85946 241768 86002 241777
rect 84990 241726 85192 241754
rect 85592 241726 85946 241754
rect 84934 241703 84990 241712
rect 75550 241632 75606 241641
rect 72896 241590 73048 241618
rect 73172 241590 73600 241618
rect 74138 241604 74304 241618
rect 74152 241590 74304 241604
rect 74704 241590 74764 241618
rect 72896 240009 72924 241590
rect 72882 240000 72938 240009
rect 72882 239935 72938 239944
rect 72804 238726 73108 238754
rect 72516 229764 72568 229770
rect 72516 229706 72568 229712
rect 73080 211138 73108 238726
rect 73172 234598 73200 241590
rect 74276 239426 74304 241590
rect 74264 239420 74316 239426
rect 74264 239362 74316 239368
rect 74736 238105 74764 241590
rect 74920 241590 75256 241618
rect 75380 241590 75550 241618
rect 74920 238882 74948 241590
rect 74908 238876 74960 238882
rect 74908 238818 74960 238824
rect 75380 238754 75408 241590
rect 75606 241590 75808 241618
rect 76024 241590 76360 241618
rect 75550 241567 75606 241576
rect 75920 239964 75972 239970
rect 75920 239906 75972 239912
rect 75288 238726 75408 238754
rect 74722 238096 74778 238105
rect 74722 238031 74778 238040
rect 73160 234592 73212 234598
rect 73160 234534 73212 234540
rect 75184 233912 75236 233918
rect 75184 233854 75236 233860
rect 74538 230616 74594 230625
rect 74538 230551 74594 230560
rect 73068 211132 73120 211138
rect 73068 211074 73120 211080
rect 73068 162920 73120 162926
rect 73068 162862 73120 162868
rect 72422 161664 72478 161673
rect 72422 161599 72478 161608
rect 71320 140752 71372 140758
rect 71320 140694 71372 140700
rect 70400 140072 70452 140078
rect 70400 140014 70452 140020
rect 70858 137184 70914 137193
rect 70858 137119 70914 137128
rect 70872 134722 70900 137119
rect 71332 134722 71360 140694
rect 72330 137864 72386 137873
rect 72330 137799 72386 137808
rect 71686 137320 71742 137329
rect 71686 137255 71742 137264
rect 71700 134722 71728 137255
rect 72344 134722 72372 137799
rect 72436 137193 72464 161599
rect 73080 142154 73108 162862
rect 73342 159352 73398 159361
rect 73342 159287 73398 159296
rect 72988 142126 73108 142154
rect 72516 138712 72568 138718
rect 72516 138654 72568 138660
rect 72422 137184 72478 137193
rect 72422 137119 72478 137128
rect 69676 134694 70104 134722
rect 70656 134694 70900 134722
rect 71024 134694 71360 134722
rect 71576 134694 71728 134722
rect 72128 134694 72372 134722
rect 72528 134722 72556 138654
rect 72988 137986 73016 142126
rect 73066 140856 73122 140865
rect 73066 140791 73122 140800
rect 73080 140758 73108 140791
rect 73068 140752 73120 140758
rect 73068 140694 73120 140700
rect 72988 137970 73200 137986
rect 72976 137964 73200 137970
rect 73028 137958 73200 137964
rect 72976 137906 73028 137912
rect 72988 137875 73016 137906
rect 73172 134994 73200 137958
rect 73172 134966 73246 134994
rect 72528 134694 72680 134722
rect 73218 134708 73246 134966
rect 73356 134722 73384 159287
rect 74262 141536 74318 141545
rect 74262 141471 74318 141480
rect 74276 134722 74304 141471
rect 73356 134694 73600 134722
rect 74152 134694 74304 134722
rect 74552 134638 74580 230551
rect 75196 157486 75224 233854
rect 75288 200802 75316 238726
rect 75932 237386 75960 239906
rect 75920 237380 75972 237386
rect 75920 237322 75972 237328
rect 76024 231810 76052 241590
rect 76898 241466 76926 241604
rect 77404 241590 77464 241618
rect 77588 241590 78016 241618
rect 78140 241590 78568 241618
rect 78692 241590 79120 241618
rect 79672 241590 79732 241618
rect 76564 241460 76616 241466
rect 76564 241402 76616 241408
rect 76886 241460 76938 241466
rect 76886 241402 76938 241408
rect 76012 231804 76064 231810
rect 76012 231746 76064 231752
rect 76576 214033 76604 241402
rect 77404 240038 77432 241590
rect 77588 240258 77616 241590
rect 78140 240938 78168 241590
rect 77496 240230 77616 240258
rect 77680 240910 78168 240938
rect 77392 240032 77444 240038
rect 77392 239974 77444 239980
rect 77496 239970 77524 240230
rect 77484 239964 77536 239970
rect 77484 239906 77536 239912
rect 77680 238754 77708 240910
rect 77944 240780 77996 240786
rect 77944 240722 77996 240728
rect 77588 238726 77708 238754
rect 77208 237380 77260 237386
rect 77208 237322 77260 237328
rect 76840 236700 76892 236706
rect 76840 236642 76892 236648
rect 76852 236065 76880 236642
rect 76838 236056 76894 236065
rect 76838 235991 76894 236000
rect 77220 231130 77248 237322
rect 77588 235278 77616 238726
rect 77576 235272 77628 235278
rect 77576 235214 77628 235220
rect 77208 231124 77260 231130
rect 77208 231066 77260 231072
rect 76748 229832 76800 229838
rect 76748 229774 76800 229780
rect 76562 214024 76618 214033
rect 76562 213959 76618 213968
rect 75276 200796 75328 200802
rect 75276 200738 75328 200744
rect 75920 173460 75972 173466
rect 75920 173402 75972 173408
rect 75276 165640 75328 165646
rect 75276 165582 75328 165588
rect 75184 157480 75236 157486
rect 75184 157422 75236 157428
rect 75196 137873 75224 157422
rect 75182 137864 75238 137873
rect 75288 137834 75316 165582
rect 75826 138680 75882 138689
rect 75826 138615 75882 138624
rect 75840 138038 75868 138615
rect 75828 138032 75880 138038
rect 75550 138000 75606 138009
rect 75828 137974 75880 137980
rect 75550 137935 75606 137944
rect 75182 137799 75238 137808
rect 75276 137828 75328 137834
rect 75276 137770 75328 137776
rect 74998 135960 75054 135969
rect 74998 135895 75054 135904
rect 75012 134722 75040 135895
rect 75564 134722 75592 137935
rect 75644 135244 75696 135250
rect 75644 135186 75696 135192
rect 74704 134694 75040 134722
rect 75256 134694 75592 134722
rect 75656 134638 75684 135186
rect 75840 134994 75868 137974
rect 75794 134966 75868 134994
rect 75794 134708 75822 134966
rect 75932 134722 75960 173402
rect 76576 138825 76604 213959
rect 76656 199436 76708 199442
rect 76656 199378 76708 199384
rect 76668 140185 76696 199378
rect 76760 173466 76788 229774
rect 76748 173460 76800 173466
rect 76748 173402 76800 173408
rect 76760 173194 76788 173402
rect 76748 173188 76800 173194
rect 76748 173130 76800 173136
rect 77956 170406 77984 240722
rect 78692 236065 78720 241590
rect 79704 240145 79732 241590
rect 80072 241590 80224 241618
rect 80348 241590 80776 241618
rect 79690 240136 79746 240145
rect 79690 240071 79746 240080
rect 79324 238060 79376 238066
rect 79324 238002 79376 238008
rect 78678 236056 78734 236065
rect 78678 235991 78734 236000
rect 78864 175296 78916 175302
rect 78864 175238 78916 175244
rect 77944 170400 77996 170406
rect 77944 170342 77996 170348
rect 77956 169794 77984 170342
rect 77392 169788 77444 169794
rect 77392 169730 77444 169736
rect 77944 169788 77996 169794
rect 77944 169730 77996 169736
rect 77298 153776 77354 153785
rect 77298 153711 77354 153720
rect 76654 140176 76710 140185
rect 76654 140111 76710 140120
rect 76562 138816 76618 138825
rect 76562 138751 76618 138760
rect 76668 134994 76696 140111
rect 77312 134994 77340 153711
rect 77404 151814 77432 169730
rect 77404 151786 77984 151814
rect 77852 137896 77904 137902
rect 77852 137838 77904 137844
rect 77864 134994 77892 137838
rect 76668 134966 76742 134994
rect 75932 134694 76176 134722
rect 76714 134708 76742 134966
rect 77266 134966 77340 134994
rect 77818 134966 77892 134994
rect 77266 134708 77294 134966
rect 77818 134708 77846 134966
rect 77956 134722 77984 151786
rect 78876 138106 78904 175238
rect 78956 142180 79008 142186
rect 78956 142122 79008 142128
rect 78864 138100 78916 138106
rect 78864 138042 78916 138048
rect 78864 137964 78916 137970
rect 78864 137906 78916 137912
rect 78876 134722 78904 137906
rect 77956 134694 78200 134722
rect 78752 134694 78904 134722
rect 78968 134722 78996 142122
rect 79336 137970 79364 238002
rect 80072 237318 80100 241590
rect 80348 238746 80376 241590
rect 81314 241466 81342 241604
rect 81452 241590 81880 241618
rect 82004 241590 82432 241618
rect 82832 241590 82984 241618
rect 83660 241590 84088 241618
rect 84212 241590 84640 241618
rect 81302 241460 81354 241466
rect 81302 241402 81354 241408
rect 81346 241360 81402 241369
rect 81346 241295 81402 241304
rect 80336 238740 80388 238746
rect 80336 238682 80388 238688
rect 80060 237312 80112 237318
rect 80060 237254 80112 237260
rect 79966 236872 80022 236881
rect 79966 236807 80022 236816
rect 79980 236065 80008 236807
rect 79966 236056 80022 236065
rect 80072 236026 80100 237254
rect 79966 235991 80022 236000
rect 80060 236020 80112 236026
rect 79980 195294 80008 235991
rect 80060 235962 80112 235968
rect 80704 236020 80756 236026
rect 80704 235962 80756 235968
rect 80716 206417 80744 235962
rect 80702 206408 80758 206417
rect 80702 206343 80758 206352
rect 79968 195288 80020 195294
rect 79968 195230 80020 195236
rect 80520 150476 80572 150482
rect 80520 150418 80572 150424
rect 80428 141500 80480 141506
rect 80428 141442 80480 141448
rect 79508 138100 79560 138106
rect 79508 138042 79560 138048
rect 79324 137964 79376 137970
rect 79324 137906 79376 137912
rect 79336 137766 79364 137906
rect 79324 137760 79376 137766
rect 79324 137702 79376 137708
rect 79520 134722 79548 138042
rect 80440 134994 80468 141442
rect 80394 134966 80468 134994
rect 78968 134694 79304 134722
rect 79520 134694 79856 134722
rect 80394 134708 80422 134966
rect 80532 134722 80560 150418
rect 81360 141409 81388 241295
rect 81452 235958 81480 241590
rect 82004 238754 82032 241590
rect 82082 240136 82138 240145
rect 82082 240071 82138 240080
rect 81544 238726 82032 238754
rect 81544 238678 81572 238726
rect 81532 238672 81584 238678
rect 81532 238614 81584 238620
rect 81440 235952 81492 235958
rect 81440 235894 81492 235900
rect 82096 180130 82124 240071
rect 82832 236042 82860 241590
rect 83660 240122 83688 241590
rect 82740 236014 82860 236042
rect 82924 240094 83688 240122
rect 82740 220114 82768 236014
rect 82924 233238 82952 240094
rect 83004 240032 83056 240038
rect 83004 239974 83056 239980
rect 83016 235890 83044 239974
rect 84212 235929 84240 241590
rect 84290 240136 84346 240145
rect 85592 240122 85620 241726
rect 85946 241703 86002 241712
rect 86682 241768 86738 241777
rect 88062 241768 88118 241777
rect 86738 241740 86848 241754
rect 86738 241726 86862 241740
rect 87952 241726 88062 241754
rect 86682 241703 86738 241712
rect 86834 241618 86862 241726
rect 96434 241768 96490 241777
rect 88118 241726 88288 241754
rect 96232 241740 96434 241754
rect 88062 241703 88118 241712
rect 84290 240071 84346 240080
rect 85500 240094 85620 240122
rect 85868 241590 86296 241618
rect 86834 241604 86908 241618
rect 86848 241590 86908 241604
rect 84198 235920 84254 235929
rect 83004 235884 83056 235890
rect 83004 235826 83056 235832
rect 83924 235884 83976 235890
rect 84198 235855 84254 235864
rect 83924 235826 83976 235832
rect 83936 234462 83964 235826
rect 84304 234546 84332 240071
rect 84028 234518 84332 234546
rect 83924 234456 83976 234462
rect 83924 234398 83976 234404
rect 82912 233232 82964 233238
rect 82912 233174 82964 233180
rect 82728 220108 82780 220114
rect 82728 220050 82780 220056
rect 84028 218754 84056 234518
rect 84108 234456 84160 234462
rect 84108 234398 84160 234404
rect 84016 218748 84068 218754
rect 84016 218690 84068 218696
rect 84120 192574 84148 234398
rect 84108 192568 84160 192574
rect 84108 192510 84160 192516
rect 82084 180124 82136 180130
rect 82084 180066 82136 180072
rect 82820 177336 82872 177342
rect 82820 177278 82872 177284
rect 81440 171148 81492 171154
rect 81440 171090 81492 171096
rect 81346 141400 81402 141409
rect 81346 141335 81402 141344
rect 81360 137902 81388 141335
rect 81348 137896 81400 137902
rect 81348 137838 81400 137844
rect 81348 136672 81400 136678
rect 81348 136614 81400 136620
rect 81360 134858 81388 136614
rect 81314 134830 81388 134858
rect 80532 134694 80776 134722
rect 81314 134708 81342 134830
rect 81452 134722 81480 171090
rect 82082 168464 82138 168473
rect 82082 168399 82138 168408
rect 81990 146976 82046 146985
rect 81990 146911 82046 146920
rect 82004 134722 82032 146911
rect 82096 138009 82124 168399
rect 82082 138000 82138 138009
rect 82082 137935 82138 137944
rect 82832 134994 82860 177278
rect 82912 173936 82964 173942
rect 82912 173878 82964 173884
rect 82924 142154 82952 173878
rect 83464 158772 83516 158778
rect 83464 158714 83516 158720
rect 83476 142866 83504 158714
rect 83556 147008 83608 147014
rect 83556 146950 83608 146956
rect 83464 142860 83516 142866
rect 83464 142802 83516 142808
rect 82924 142126 83504 142154
rect 83372 136740 83424 136746
rect 83372 136682 83424 136688
rect 82786 134966 82860 134994
rect 81452 134694 81880 134722
rect 82004 134694 82432 134722
rect 82786 134708 82814 134966
rect 83384 134858 83412 136682
rect 83338 134830 83412 134858
rect 83338 134708 83366 134830
rect 83476 134722 83504 142126
rect 83568 136678 83596 146950
rect 85500 145625 85528 240094
rect 85868 238754 85896 241590
rect 86224 240100 86276 240106
rect 86224 240042 86276 240048
rect 85592 238726 85896 238754
rect 85592 236609 85620 238726
rect 85578 236600 85634 236609
rect 85578 236535 85634 236544
rect 86236 233170 86264 240042
rect 86880 240009 86908 241590
rect 87064 241590 87400 241618
rect 87064 240106 87092 241590
rect 87052 240100 87104 240106
rect 87052 240042 87104 240048
rect 86866 240000 86922 240009
rect 86866 239935 86922 239944
rect 86224 233164 86276 233170
rect 86224 233106 86276 233112
rect 86236 199442 86264 233106
rect 86868 229764 86920 229770
rect 86868 229706 86920 229712
rect 86224 199436 86276 199442
rect 86224 199378 86276 199384
rect 86224 170468 86276 170474
rect 86224 170410 86276 170416
rect 85486 145616 85542 145625
rect 85486 145551 85542 145560
rect 84566 143712 84622 143721
rect 84566 143647 84622 143656
rect 84474 139632 84530 139641
rect 84474 139567 84530 139576
rect 83556 136672 83608 136678
rect 83556 136614 83608 136620
rect 84488 134994 84516 139567
rect 84442 134966 84516 134994
rect 83476 134694 83904 134722
rect 84442 134708 84470 134966
rect 84580 134722 84608 143647
rect 86040 142860 86092 142866
rect 86040 142802 86092 142808
rect 85486 136776 85542 136785
rect 85486 136711 85542 136720
rect 85500 134722 85528 136711
rect 85948 136672 86000 136678
rect 85948 136614 86000 136620
rect 85960 134858 85988 136614
rect 84580 134694 85008 134722
rect 85376 134694 85528 134722
rect 85914 134830 85988 134858
rect 85914 134708 85942 134830
rect 86052 134722 86080 142802
rect 86236 136746 86264 170410
rect 86316 165708 86368 165714
rect 86316 165650 86368 165656
rect 86328 137329 86356 165650
rect 86774 156632 86830 156641
rect 86774 156567 86830 156576
rect 86788 142866 86816 156567
rect 86880 152590 86908 229706
rect 88260 205018 88288 241726
rect 96218 241726 96434 241740
rect 92110 241632 92166 241641
rect 88504 241590 88564 241618
rect 88536 239494 88564 241590
rect 88628 241590 89056 241618
rect 89608 241590 89668 241618
rect 90160 241590 90312 241618
rect 88524 239488 88576 239494
rect 88524 239430 88576 239436
rect 88628 238754 88656 241590
rect 89640 239873 89668 241590
rect 89626 239864 89682 239873
rect 89626 239799 89682 239808
rect 90284 239737 90312 241590
rect 90376 241590 90712 241618
rect 91112 241590 91264 241618
rect 91664 241590 91816 241618
rect 90270 239728 90326 239737
rect 90270 239663 90326 239672
rect 88352 238726 88656 238754
rect 88352 234433 88380 238726
rect 90376 234614 90404 241590
rect 91006 235784 91062 235793
rect 91006 235719 91062 235728
rect 89732 234586 90404 234614
rect 88338 234424 88394 234433
rect 88338 234359 88394 234368
rect 89732 215286 89760 234586
rect 89720 215280 89772 215286
rect 89720 215222 89772 215228
rect 88248 205012 88300 205018
rect 88248 204954 88300 204960
rect 91020 178090 91048 235719
rect 91112 232558 91140 241590
rect 91664 240145 91692 241590
rect 92166 241590 92428 241618
rect 92110 241567 92166 241576
rect 91650 240136 91706 240145
rect 91650 240071 91706 240080
rect 91100 232552 91152 232558
rect 91100 232494 91152 232500
rect 92400 211041 92428 241590
rect 92906 241505 92934 241604
rect 93136 241590 93472 241618
rect 94024 241590 94360 241618
rect 94576 241590 95004 241618
rect 92892 241496 92948 241505
rect 92892 241431 92948 241440
rect 93136 241233 93164 241590
rect 93122 241224 93178 241233
rect 93122 241159 93178 241168
rect 92386 211032 92442 211041
rect 92386 210967 92442 210976
rect 93136 206310 93164 241159
rect 94332 240145 94360 241590
rect 94318 240136 94374 240145
rect 94318 240071 94374 240080
rect 94870 240136 94926 240145
rect 94870 240071 94926 240080
rect 93766 237008 93822 237017
rect 93766 236943 93822 236952
rect 93124 206304 93176 206310
rect 93124 206246 93176 206252
rect 93780 180878 93808 236943
rect 94884 234614 94912 240071
rect 94976 238082 95004 241590
rect 95068 241590 95128 241618
rect 95680 241590 95924 241618
rect 95068 238513 95096 241590
rect 95332 241528 95384 241534
rect 95332 241470 95384 241476
rect 95054 238504 95110 238513
rect 95054 238439 95110 238448
rect 95068 238241 95096 238439
rect 95054 238232 95110 238241
rect 95054 238167 95110 238176
rect 94976 238054 95188 238082
rect 94884 234586 95096 234614
rect 95068 209774 95096 234586
rect 95160 227050 95188 238054
rect 95238 237280 95294 237289
rect 95238 237215 95294 237224
rect 95252 236706 95280 237215
rect 95240 236700 95292 236706
rect 95240 236642 95292 236648
rect 95344 234614 95372 241470
rect 95896 241398 95924 241590
rect 96218 241534 96246 241726
rect 96434 241703 96490 241712
rect 96770 241760 96896 241788
rect 96206 241528 96258 241534
rect 96206 241470 96258 241476
rect 96770 241482 96798 241760
rect 96896 241742 96948 241748
rect 96908 241590 97336 241618
rect 97736 241590 97888 241618
rect 96770 241454 96844 241482
rect 95884 241392 95936 241398
rect 95884 241334 95936 241340
rect 95252 234586 95372 234614
rect 95148 227044 95200 227050
rect 95148 226986 95200 226992
rect 95148 225616 95200 225622
rect 95148 225558 95200 225564
rect 94700 209746 95096 209774
rect 94700 207058 94728 209746
rect 94688 207052 94740 207058
rect 94688 206994 94740 207000
rect 93124 180872 93176 180878
rect 93124 180814 93176 180820
rect 93768 180872 93820 180878
rect 93768 180814 93820 180820
rect 90364 178084 90416 178090
rect 90364 178026 90416 178032
rect 91008 178084 91060 178090
rect 91008 178026 91060 178032
rect 87602 176760 87658 176769
rect 87602 176695 87658 176704
rect 86958 167104 87014 167113
rect 86958 167039 87014 167048
rect 86868 152584 86920 152590
rect 86868 152526 86920 152532
rect 86776 142860 86828 142866
rect 86776 142802 86828 142808
rect 86314 137320 86370 137329
rect 86314 137255 86370 137264
rect 86224 136740 86276 136746
rect 86224 136682 86276 136688
rect 86972 134994 87000 167039
rect 87144 159384 87196 159390
rect 87144 159326 87196 159332
rect 87052 138644 87104 138650
rect 87052 138586 87104 138592
rect 87064 136678 87092 138586
rect 87052 136672 87104 136678
rect 87052 136614 87104 136620
rect 86972 134966 87046 134994
rect 86052 134694 86480 134722
rect 87018 134708 87046 134966
rect 87156 134722 87184 159326
rect 87512 145580 87564 145586
rect 87512 145522 87564 145528
rect 87524 144906 87552 145522
rect 87512 144900 87564 144906
rect 87512 144842 87564 144848
rect 87524 138014 87552 144842
rect 87616 139641 87644 176695
rect 88982 174040 89038 174049
rect 88982 173975 89038 173984
rect 88340 152516 88392 152522
rect 88340 152458 88392 152464
rect 87602 139632 87658 139641
rect 87602 139567 87658 139576
rect 87524 137986 87736 138014
rect 87708 134722 87736 137986
rect 88352 134722 88380 152458
rect 88996 136785 89024 173975
rect 89166 143712 89222 143721
rect 89166 143647 89222 143656
rect 89180 142769 89208 143647
rect 89166 142760 89222 142769
rect 89166 142695 89222 142704
rect 89626 140856 89682 140865
rect 89626 140791 89682 140800
rect 89352 137012 89404 137018
rect 89352 136954 89404 136960
rect 88982 136776 89038 136785
rect 88982 136711 89038 136720
rect 89364 134722 89392 136954
rect 89640 134994 89668 140791
rect 90376 137018 90404 178026
rect 91744 172576 91796 172582
rect 91744 172518 91796 172524
rect 91008 164960 91060 164966
rect 91008 164902 91060 164908
rect 90456 157412 90508 157418
rect 90456 157354 90508 157360
rect 90468 147014 90496 157354
rect 90456 147008 90508 147014
rect 90456 146950 90508 146956
rect 90916 146940 90968 146946
rect 90916 146882 90968 146888
rect 90824 138712 90876 138718
rect 90824 138654 90876 138660
rect 90364 137012 90416 137018
rect 90364 136954 90416 136960
rect 90272 136672 90324 136678
rect 90272 136614 90324 136620
rect 87156 134694 87584 134722
rect 87708 134694 87952 134722
rect 88352 134694 88504 134722
rect 89056 134694 89392 134722
rect 89594 134966 89668 134994
rect 89594 134708 89622 134966
rect 90284 134722 90312 136614
rect 90836 134722 90864 138654
rect 90928 136082 90956 146882
rect 91020 138014 91048 164902
rect 91652 143608 91704 143614
rect 91652 143550 91704 143556
rect 91020 137986 91140 138014
rect 91112 136105 91140 137986
rect 91664 136610 91692 143550
rect 91756 136678 91784 172518
rect 92478 171184 92534 171193
rect 92478 171119 92534 171128
rect 91744 136672 91796 136678
rect 91744 136614 91796 136620
rect 92388 136672 92440 136678
rect 92388 136614 92440 136620
rect 91652 136604 91704 136610
rect 91652 136546 91704 136552
rect 91098 136096 91154 136105
rect 90928 136054 91048 136082
rect 91020 135998 91048 136054
rect 91098 136031 91154 136040
rect 91282 136096 91338 136105
rect 91282 136031 91338 136040
rect 91008 135992 91060 135998
rect 91060 135940 91140 135946
rect 91008 135934 91140 135940
rect 91020 135918 91140 135934
rect 91112 134994 91140 135918
rect 89976 134694 90312 134722
rect 90528 134694 90864 134722
rect 91066 134966 91140 134994
rect 91066 134708 91094 134966
rect 91296 134722 91324 136031
rect 92400 134722 92428 136614
rect 92492 134994 92520 171119
rect 92662 161528 92718 161537
rect 92662 161463 92718 161472
rect 92492 134966 92566 134994
rect 91296 134694 91632 134722
rect 92184 134694 92428 134722
rect 92538 134708 92566 134966
rect 92676 134722 92704 161463
rect 93030 144120 93086 144129
rect 93030 144055 93086 144064
rect 93044 134858 93072 144055
rect 93136 136678 93164 180814
rect 93860 169040 93912 169046
rect 93860 168982 93912 168988
rect 93124 136672 93176 136678
rect 93124 136614 93176 136620
rect 93044 134830 93256 134858
rect 93228 134722 93256 134830
rect 93872 134722 93900 168982
rect 94700 138014 94728 206994
rect 94962 143984 95018 143993
rect 94962 143919 95018 143928
rect 94700 137986 94820 138014
rect 94136 135244 94188 135250
rect 94136 135186 94188 135192
rect 94148 135153 94176 135186
rect 94134 135144 94190 135153
rect 94134 135079 94190 135088
rect 92676 134694 93104 134722
rect 93228 134694 93656 134722
rect 93872 134694 94208 134722
rect 74540 134632 74592 134638
rect 68848 133385 68876 134574
rect 69400 134558 69552 134586
rect 74540 134574 74592 134580
rect 75644 134632 75696 134638
rect 75644 134574 75696 134580
rect 94576 134014 94728 134042
rect 94700 133958 94728 134014
rect 94688 133952 94740 133958
rect 94688 133894 94740 133900
rect 68834 133376 68890 133385
rect 68834 133311 68890 133320
rect 94594 124944 94650 124953
rect 94594 124879 94650 124888
rect 94608 124166 94636 124879
rect 94596 124160 94648 124166
rect 94596 124102 94648 124108
rect 68664 113146 68968 113174
rect 67824 93832 67876 93838
rect 67824 93774 67876 93780
rect 67836 93401 67864 93774
rect 67822 93392 67878 93401
rect 67822 93327 67878 93336
rect 67836 60625 67864 93327
rect 68480 92806 68816 92834
rect 68006 91760 68062 91769
rect 68006 91695 68062 91704
rect 68020 91089 68048 91695
rect 68006 91080 68062 91089
rect 68006 91015 68062 91024
rect 68480 90370 68508 92806
rect 68940 92750 68968 113146
rect 94608 93854 94636 124102
rect 94792 122834 94820 137986
rect 94976 126954 95004 143919
rect 95160 138281 95188 225558
rect 95146 138272 95202 138281
rect 95146 138207 95202 138216
rect 94964 126948 95016 126954
rect 94964 126890 95016 126896
rect 94700 122806 94820 122834
rect 94700 113174 94728 122806
rect 94700 113146 94820 113174
rect 94608 93826 94728 93854
rect 68928 92744 68980 92750
rect 68928 92686 68980 92692
rect 69170 92562 69198 92820
rect 69722 92750 69750 92820
rect 69710 92744 69762 92750
rect 69710 92686 69762 92692
rect 70274 92698 70302 92820
rect 69722 92562 69750 92686
rect 70274 92670 70348 92698
rect 69170 92534 69244 92562
rect 69722 92534 69796 92562
rect 70320 92546 70348 92670
rect 70826 92562 70854 92820
rect 71194 92562 71222 92820
rect 68468 90364 68520 90370
rect 68468 90306 68520 90312
rect 69216 88330 69244 92534
rect 69204 88324 69256 88330
rect 69204 88266 69256 88272
rect 69662 87544 69718 87553
rect 69662 87479 69718 87488
rect 67822 60616 67878 60625
rect 67822 60551 67878 60560
rect 68928 47592 68980 47598
rect 68928 47534 68980 47540
rect 67732 33788 67784 33794
rect 67732 33730 67784 33736
rect 68940 3534 68968 47534
rect 69676 20670 69704 87479
rect 69768 70281 69796 92534
rect 70308 92540 70360 92546
rect 70308 92482 70360 92488
rect 70780 92534 70854 92562
rect 71148 92534 71222 92562
rect 71746 92562 71774 92820
rect 72298 92562 72326 92820
rect 72850 92750 72878 92820
rect 72838 92744 72890 92750
rect 72976 92744 73028 92750
rect 72838 92686 72890 92692
rect 72974 92712 72976 92721
rect 73028 92712 73030 92721
rect 72974 92647 73030 92656
rect 73402 92562 73430 92820
rect 71746 92534 71820 92562
rect 70320 91225 70348 92482
rect 70306 91216 70362 91225
rect 70306 91151 70362 91160
rect 70780 91050 70808 92534
rect 71042 91216 71098 91225
rect 71042 91151 71098 91160
rect 70768 91044 70820 91050
rect 70768 90986 70820 90992
rect 71056 71777 71084 91151
rect 71148 91089 71176 92534
rect 71134 91080 71190 91089
rect 71134 91015 71190 91024
rect 71792 84182 71820 92534
rect 71884 92534 72326 92562
rect 73172 92534 73430 92562
rect 73770 92562 73798 92820
rect 74322 92562 74350 92820
rect 74874 92698 74902 92820
rect 74828 92670 74902 92698
rect 73770 92534 73844 92562
rect 71780 84176 71832 84182
rect 71780 84118 71832 84124
rect 71686 76528 71742 76537
rect 71686 76463 71742 76472
rect 71042 71768 71098 71777
rect 71042 71703 71098 71712
rect 69754 70272 69810 70281
rect 69754 70207 69810 70216
rect 70308 28280 70360 28286
rect 70308 28222 70360 28228
rect 69664 20664 69716 20670
rect 69664 20606 69716 20612
rect 70122 14512 70178 14521
rect 70122 14447 70178 14456
rect 69112 3596 69164 3602
rect 69112 3538 69164 3544
rect 64328 3528 64380 3534
rect 64328 3470 64380 3476
rect 64788 3528 64840 3534
rect 64788 3470 64840 3476
rect 65524 3528 65576 3534
rect 65524 3470 65576 3476
rect 66168 3528 66220 3534
rect 66168 3470 66220 3476
rect 67916 3528 67968 3534
rect 67916 3470 67968 3476
rect 68928 3528 68980 3534
rect 68928 3470 68980 3476
rect 64340 480 64368 3470
rect 65536 480 65564 3470
rect 66720 3460 66772 3466
rect 66720 3402 66772 3408
rect 66732 480 66760 3402
rect 67928 480 67956 3470
rect 69124 480 69152 3538
rect 70136 3482 70164 14447
rect 70320 6914 70348 28222
rect 71700 6914 71728 76463
rect 71884 63510 71912 92534
rect 73172 84114 73200 92534
rect 73816 86970 73844 92534
rect 74276 92534 74350 92562
rect 74540 92608 74592 92614
rect 74540 92550 74592 92556
rect 74276 90953 74304 92534
rect 74262 90944 74318 90953
rect 74262 90879 74318 90888
rect 73804 86964 73856 86970
rect 73804 86906 73856 86912
rect 74276 84194 74304 90879
rect 73816 84166 74304 84194
rect 73160 84108 73212 84114
rect 73160 84050 73212 84056
rect 71872 63504 71924 63510
rect 71872 63446 71924 63452
rect 73816 56574 73844 84166
rect 74552 64802 74580 92550
rect 74828 91089 74856 92670
rect 75426 92562 75454 92820
rect 75794 92614 75822 92820
rect 75782 92608 75834 92614
rect 75426 92534 75500 92562
rect 76346 92562 76374 92820
rect 76898 92562 76926 92820
rect 77450 92562 77478 92820
rect 75782 92550 75834 92556
rect 74814 91080 74870 91089
rect 74814 91015 74870 91024
rect 75472 89622 75500 92534
rect 76300 92534 76374 92562
rect 76576 92534 76926 92562
rect 77312 92534 77478 92562
rect 78002 92562 78030 92820
rect 78370 92562 78398 92820
rect 78922 92562 78950 92820
rect 79474 92562 79502 92820
rect 80026 92562 80054 92820
rect 80578 92562 80606 92820
rect 80946 92562 80974 92820
rect 81498 92562 81526 92820
rect 78002 92534 78076 92562
rect 78370 92534 78444 92562
rect 78922 92534 78996 92562
rect 79474 92534 79548 92562
rect 80026 92534 80100 92562
rect 76300 92449 76328 92534
rect 76286 92440 76342 92449
rect 76286 92375 76342 92384
rect 75460 89616 75512 89622
rect 75460 89558 75512 89564
rect 76576 84194 76604 92534
rect 75932 84166 76604 84194
rect 75932 82822 75960 84166
rect 75920 82816 75972 82822
rect 75920 82758 75972 82764
rect 77312 81326 77340 92534
rect 78048 89865 78076 92534
rect 78034 89856 78090 89865
rect 78034 89791 78090 89800
rect 78416 85513 78444 92534
rect 78968 90953 78996 92534
rect 79520 92177 79548 92534
rect 79506 92168 79562 92177
rect 79506 92103 79562 92112
rect 78954 90944 79010 90953
rect 78954 90879 79010 90888
rect 80072 88262 80100 92534
rect 80164 92534 80606 92562
rect 80716 92534 80974 92562
rect 81452 92534 81526 92562
rect 82050 92562 82078 92820
rect 82602 92562 82630 92820
rect 82970 92698 82998 92820
rect 82970 92670 83044 92698
rect 82050 92534 82124 92562
rect 80060 88256 80112 88262
rect 80060 88198 80112 88204
rect 78402 85504 78458 85513
rect 78402 85439 78458 85448
rect 77300 81320 77352 81326
rect 77300 81262 77352 81268
rect 75828 75200 75880 75206
rect 75828 75142 75880 75148
rect 74540 64796 74592 64802
rect 74540 64738 74592 64744
rect 73804 56568 73856 56574
rect 73804 56510 73856 56516
rect 73068 49020 73120 49026
rect 73068 48962 73120 48968
rect 70228 6886 70348 6914
rect 71516 6886 71728 6914
rect 70228 3602 70256 6886
rect 70216 3596 70268 3602
rect 70216 3538 70268 3544
rect 70136 3454 70348 3482
rect 70320 480 70348 3454
rect 71516 480 71544 6886
rect 73080 3534 73108 48962
rect 75840 3534 75868 75142
rect 80164 68950 80192 92534
rect 80716 84194 80744 92534
rect 80256 84166 80744 84194
rect 80256 78606 80284 84166
rect 80244 78600 80296 78606
rect 80244 78542 80296 78548
rect 80152 68944 80204 68950
rect 80152 68886 80204 68892
rect 81452 66230 81480 92534
rect 82096 89457 82124 92534
rect 82280 92534 82630 92562
rect 82082 89448 82138 89457
rect 82082 89383 82138 89392
rect 82280 88233 82308 92534
rect 83016 89321 83044 92670
rect 83522 92562 83550 92820
rect 83200 92534 83550 92562
rect 84074 92562 84102 92820
rect 84626 92698 84654 92820
rect 84626 92670 84700 92698
rect 84074 92534 84148 92562
rect 83002 89312 83058 89321
rect 83002 89247 83058 89256
rect 82266 88224 82322 88233
rect 82266 88159 82322 88168
rect 82280 84194 82308 88159
rect 83200 84194 83228 92534
rect 84120 88097 84148 92534
rect 84672 91050 84700 92670
rect 85178 92562 85206 92820
rect 84856 92534 85206 92562
rect 85546 92562 85574 92820
rect 86098 92698 86126 92820
rect 86098 92670 86172 92698
rect 85546 92534 85620 92562
rect 84660 91044 84712 91050
rect 84660 90986 84712 90992
rect 84106 88088 84162 88097
rect 84106 88023 84162 88032
rect 84856 84194 84884 92534
rect 82096 84166 82308 84194
rect 82832 84166 83228 84194
rect 84212 84166 84884 84194
rect 81440 66224 81492 66230
rect 81440 66166 81492 66172
rect 82096 57934 82124 84166
rect 82832 81433 82860 84166
rect 82818 81424 82874 81433
rect 82818 81359 82874 81368
rect 83462 62792 83518 62801
rect 83462 62727 83518 62736
rect 82084 57928 82136 57934
rect 82084 57870 82136 57876
rect 77208 54528 77260 54534
rect 77208 54470 77260 54476
rect 77220 3534 77248 54470
rect 79968 31068 80020 31074
rect 79968 31010 80020 31016
rect 78588 18624 78640 18630
rect 78588 18566 78640 18572
rect 72608 3528 72660 3534
rect 72608 3470 72660 3476
rect 73068 3528 73120 3534
rect 75000 3528 75052 3534
rect 73068 3470 73120 3476
rect 73802 3496 73858 3505
rect 72620 480 72648 3470
rect 75000 3470 75052 3476
rect 75828 3528 75880 3534
rect 75828 3470 75880 3476
rect 76196 3528 76248 3534
rect 76196 3470 76248 3476
rect 77208 3528 77260 3534
rect 77208 3470 77260 3476
rect 73802 3431 73858 3440
rect 73816 480 73844 3431
rect 75012 480 75040 3470
rect 76208 480 76236 3470
rect 77392 3052 77444 3058
rect 77392 2994 77444 3000
rect 77404 480 77432 2994
rect 78600 480 78628 18566
rect 79322 15872 79378 15881
rect 79322 15807 79378 15816
rect 79336 3058 79364 15807
rect 79980 6914 80008 31010
rect 82082 8936 82138 8945
rect 82082 8871 82138 8880
rect 79704 6886 80008 6914
rect 79324 3052 79376 3058
rect 79324 2994 79376 3000
rect 79704 480 79732 6886
rect 80888 3596 80940 3602
rect 80888 3538 80940 3544
rect 80900 480 80928 3538
rect 82096 480 82124 8871
rect 83476 3602 83504 62727
rect 84212 57866 84240 84166
rect 85592 62082 85620 92534
rect 86144 86873 86172 92670
rect 86650 92562 86678 92820
rect 87202 92698 87230 92820
rect 87202 92670 87276 92698
rect 86328 92534 86678 92562
rect 86130 86864 86186 86873
rect 86130 86799 86186 86808
rect 86328 84194 86356 92534
rect 87248 85377 87276 92670
rect 87570 92562 87598 92820
rect 88122 92562 88150 92820
rect 88674 92562 88702 92820
rect 87340 92534 87598 92562
rect 87800 92534 88150 92562
rect 88352 92534 88702 92562
rect 89226 92562 89254 92820
rect 89778 92562 89806 92820
rect 90146 92682 90174 92820
rect 90134 92676 90186 92682
rect 90134 92618 90186 92624
rect 90698 92562 90726 92820
rect 91008 92676 91060 92682
rect 91008 92618 91060 92624
rect 89226 92534 89300 92562
rect 89778 92534 89852 92562
rect 87234 85368 87290 85377
rect 87234 85303 87290 85312
rect 87340 85218 87368 92534
rect 85684 84166 86356 84194
rect 86972 85190 87368 85218
rect 85684 79966 85712 84166
rect 85672 79960 85724 79966
rect 85672 79902 85724 79908
rect 86868 72480 86920 72486
rect 86868 72422 86920 72428
rect 85580 62076 85632 62082
rect 85580 62018 85632 62024
rect 84200 57860 84252 57866
rect 84200 57802 84252 57808
rect 86776 26920 86828 26926
rect 86776 26862 86828 26868
rect 84108 25560 84160 25566
rect 84108 25502 84160 25508
rect 83464 3596 83516 3602
rect 83464 3538 83516 3544
rect 84120 3534 84148 25502
rect 85486 17232 85542 17241
rect 85486 17167 85542 17176
rect 85500 3534 85528 17167
rect 86788 3534 86816 26862
rect 83280 3528 83332 3534
rect 83280 3470 83332 3476
rect 84108 3528 84160 3534
rect 84108 3470 84160 3476
rect 84476 3528 84528 3534
rect 84476 3470 84528 3476
rect 85488 3528 85540 3534
rect 85488 3470 85540 3476
rect 85672 3528 85724 3534
rect 85672 3470 85724 3476
rect 86776 3528 86828 3534
rect 86776 3470 86828 3476
rect 83292 480 83320 3470
rect 84488 480 84516 3470
rect 85684 480 85712 3470
rect 86880 480 86908 72422
rect 86972 66162 87000 85190
rect 87800 84194 87828 92534
rect 87064 84166 87828 84194
rect 87064 78674 87092 84166
rect 88246 82104 88302 82113
rect 88246 82039 88302 82048
rect 87052 78668 87104 78674
rect 87052 78610 87104 78616
rect 86960 66156 87012 66162
rect 86960 66098 87012 66104
rect 88260 6914 88288 82039
rect 88352 60722 88380 92534
rect 89272 88233 89300 92534
rect 89258 88224 89314 88233
rect 89258 88159 89314 88168
rect 89824 86737 89852 92534
rect 89916 92534 90726 92562
rect 89810 86728 89866 86737
rect 89810 86663 89866 86672
rect 89628 73840 89680 73846
rect 89628 73782 89680 73788
rect 88340 60716 88392 60722
rect 88340 60658 88392 60664
rect 87984 6886 88288 6914
rect 87984 480 88012 6886
rect 89640 3534 89668 73782
rect 89916 69018 89944 92534
rect 91020 92449 91048 92618
rect 91250 92562 91278 92820
rect 91802 92562 91830 92820
rect 92354 92562 92382 92820
rect 92722 92562 92750 92820
rect 93274 92721 93302 92820
rect 93260 92712 93316 92721
rect 93826 92698 93854 92820
rect 94378 92750 94406 92820
rect 94366 92744 94418 92750
rect 93826 92670 93900 92698
rect 94366 92686 94418 92692
rect 93260 92647 93316 92656
rect 91250 92534 91324 92562
rect 91802 92534 91876 92562
rect 92354 92534 92428 92562
rect 91006 92440 91062 92449
rect 91006 92375 91062 92384
rect 89904 69012 89956 69018
rect 89904 68954 89956 68960
rect 91020 67590 91048 92375
rect 91296 89593 91324 92534
rect 91848 92313 91876 92534
rect 92400 92449 92428 92534
rect 92492 92534 92750 92562
rect 93274 92562 93302 92647
rect 93274 92534 93348 92562
rect 92386 92440 92442 92449
rect 92386 92375 92442 92384
rect 91834 92304 91890 92313
rect 91834 92239 91890 92248
rect 91282 89584 91338 89593
rect 91282 89519 91338 89528
rect 92492 82754 92520 92534
rect 93320 84194 93348 92534
rect 93872 90302 93900 92670
rect 93860 90296 93912 90302
rect 93860 90238 93912 90244
rect 94700 86601 94728 93826
rect 94792 92449 94820 113146
rect 95148 93152 95200 93158
rect 95148 93094 95200 93100
rect 94778 92440 94834 92449
rect 94778 92375 94834 92384
rect 95056 90296 95108 90302
rect 95056 90238 95108 90244
rect 94686 86592 94742 86601
rect 94686 86527 94742 86536
rect 95068 84194 95096 90238
rect 95160 88262 95188 93094
rect 95252 92750 95280 234586
rect 95516 147076 95568 147082
rect 95516 147018 95568 147024
rect 95422 138272 95478 138281
rect 95422 138207 95478 138216
rect 95436 124137 95464 138207
rect 95528 127673 95556 147018
rect 95514 127664 95570 127673
rect 95514 127599 95570 127608
rect 95422 124128 95478 124137
rect 95422 124063 95478 124072
rect 95330 120320 95386 120329
rect 95330 120255 95386 120264
rect 95240 92744 95292 92750
rect 95240 92686 95292 92692
rect 95148 88256 95200 88262
rect 95148 88198 95200 88204
rect 93320 84166 93716 84194
rect 95068 84166 95188 84194
rect 92480 82748 92532 82754
rect 92480 82690 92532 82696
rect 91008 67584 91060 67590
rect 91008 67526 91060 67532
rect 93688 64870 93716 84166
rect 95160 77246 95188 84166
rect 95148 77240 95200 77246
rect 95148 77182 95200 77188
rect 95344 71738 95372 120255
rect 95896 90302 95924 241334
rect 96816 240145 96844 241454
rect 96802 240136 96858 240145
rect 96802 240071 96858 240080
rect 96908 234614 96936 241590
rect 97736 241369 97764 241590
rect 97722 241360 97778 241369
rect 97722 241295 97778 241304
rect 96632 234586 96936 234614
rect 96632 204950 96660 234586
rect 97736 233481 97764 241295
rect 98000 239488 98052 239494
rect 98000 239430 98052 239436
rect 98012 236774 98040 239430
rect 98000 236768 98052 236774
rect 98000 236710 98052 236716
rect 97816 236020 97868 236026
rect 97816 235962 97868 235968
rect 97262 233472 97318 233481
rect 97262 233407 97318 233416
rect 97722 233472 97778 233481
rect 97722 233407 97778 233416
rect 97276 211818 97304 233407
rect 97264 211812 97316 211818
rect 97264 211754 97316 211760
rect 96620 204944 96672 204950
rect 96620 204886 96672 204892
rect 97828 166297 97856 235962
rect 97908 233912 97960 233918
rect 97908 233854 97960 233860
rect 97262 166288 97318 166297
rect 97262 166223 97318 166232
rect 97814 166288 97870 166297
rect 97814 166223 97870 166232
rect 96526 147112 96582 147121
rect 96526 147047 96528 147056
rect 96580 147047 96582 147056
rect 96528 147018 96580 147024
rect 96712 135244 96764 135250
rect 96712 135186 96764 135192
rect 96724 133929 96752 135186
rect 96710 133920 96766 133929
rect 96710 133855 96766 133864
rect 96712 133340 96764 133346
rect 96712 133282 96764 133288
rect 96724 133113 96752 133282
rect 96710 133104 96766 133113
rect 96710 133039 96766 133048
rect 96620 132456 96672 132462
rect 96620 132398 96672 132404
rect 96632 131481 96660 132398
rect 96618 131472 96674 131481
rect 96618 131407 96674 131416
rect 96620 131028 96672 131034
rect 96620 130970 96672 130976
rect 96632 130121 96660 130970
rect 96618 130112 96674 130121
rect 96618 130047 96674 130056
rect 96712 129668 96764 129674
rect 96712 129610 96764 129616
rect 96724 128489 96752 129610
rect 96710 128480 96766 128489
rect 96710 128415 96766 128424
rect 97172 126880 97224 126886
rect 97172 126822 97224 126828
rect 97184 126313 97212 126822
rect 97170 126304 97226 126313
rect 97170 126239 97226 126248
rect 97276 122505 97304 166223
rect 97920 162858 97948 233854
rect 98104 202230 98132 247007
rect 98196 233918 98224 270671
rect 98288 264246 98316 282526
rect 98276 264240 98328 264246
rect 98276 264182 98328 264188
rect 98380 248414 98408 319466
rect 99288 316804 99340 316810
rect 99288 316746 99340 316752
rect 99300 292574 99328 316746
rect 99024 292546 99328 292574
rect 98460 284436 98512 284442
rect 98460 284378 98512 284384
rect 98472 278050 98500 284378
rect 99024 283506 99052 292546
rect 98624 283478 99052 283506
rect 98736 282260 98788 282266
rect 98736 282202 98788 282208
rect 98460 278044 98512 278050
rect 98460 277986 98512 277992
rect 98748 268433 98776 282202
rect 99380 278724 99432 278730
rect 99380 278666 99432 278672
rect 99392 277817 99420 278666
rect 99378 277808 99434 277817
rect 99378 277743 99434 277752
rect 99288 271584 99340 271590
rect 99288 271526 99340 271532
rect 99300 271289 99328 271526
rect 99286 271280 99342 271289
rect 99286 271215 99342 271224
rect 98734 268424 98790 268433
rect 98734 268359 98790 268368
rect 99288 263628 99340 263634
rect 99288 263570 99340 263576
rect 98380 248386 98500 248414
rect 98472 242570 98500 248386
rect 99196 248396 99248 248402
rect 99196 248338 99248 248344
rect 99208 247625 99236 248338
rect 99194 247616 99250 247625
rect 99194 247551 99250 247560
rect 98426 242542 98500 242570
rect 98426 241890 98454 242542
rect 98288 241876 98454 241890
rect 98288 241862 98440 241876
rect 98288 240106 98316 241862
rect 98276 240100 98328 240106
rect 98276 240042 98328 240048
rect 98184 233912 98236 233918
rect 98184 233854 98236 233860
rect 98644 213920 98696 213926
rect 98644 213862 98696 213868
rect 98092 202224 98144 202230
rect 98092 202166 98144 202172
rect 98104 200114 98132 202166
rect 98012 200086 98132 200114
rect 97448 162852 97500 162858
rect 97448 162794 97500 162800
rect 97908 162852 97960 162858
rect 97908 162794 97960 162800
rect 97460 162178 97488 162794
rect 97448 162172 97500 162178
rect 97448 162114 97500 162120
rect 97460 128354 97488 162114
rect 97540 144356 97592 144362
rect 97540 144298 97592 144304
rect 97552 129305 97580 144298
rect 97906 130928 97962 130937
rect 97906 130863 97962 130872
rect 97920 129742 97948 130863
rect 97908 129736 97960 129742
rect 97908 129678 97960 129684
rect 97538 129296 97594 129305
rect 97538 129231 97594 129240
rect 97368 128326 97488 128354
rect 97920 128330 97948 129678
rect 97368 123321 97396 128326
rect 97644 128302 97948 128330
rect 97448 125588 97500 125594
rect 97448 125530 97500 125536
rect 97460 124681 97488 125530
rect 97446 124672 97502 124681
rect 97446 124607 97502 124616
rect 97354 123312 97410 123321
rect 97354 123247 97410 123256
rect 97644 122834 97672 128302
rect 97908 128240 97960 128246
rect 97908 128182 97960 128188
rect 97920 127129 97948 128182
rect 97906 127120 97962 127129
rect 97906 127055 97962 127064
rect 97368 122806 97672 122834
rect 97262 122496 97318 122505
rect 97262 122431 97318 122440
rect 97172 121440 97224 121446
rect 97172 121382 97224 121388
rect 97184 120873 97212 121382
rect 97170 120864 97226 120873
rect 97170 120799 97226 120808
rect 96068 120352 96120 120358
rect 96066 120320 96068 120329
rect 96120 120320 96122 120329
rect 96066 120255 96122 120264
rect 97264 118720 97316 118726
rect 97264 118662 97316 118668
rect 97276 114073 97304 118662
rect 97262 114064 97318 114073
rect 97262 113999 97318 114008
rect 96804 111104 96856 111110
rect 96802 111072 96804 111081
rect 96856 111072 96858 111081
rect 96802 111007 96858 111016
rect 97170 109712 97226 109721
rect 97170 109647 97226 109656
rect 97184 109070 97212 109647
rect 97172 109064 97224 109070
rect 97172 109006 97224 109012
rect 95976 108316 96028 108322
rect 95976 108258 96028 108264
rect 95884 90296 95936 90302
rect 95884 90238 95936 90244
rect 95988 89622 96016 108258
rect 96620 97708 96672 97714
rect 96620 97650 96672 97656
rect 96632 96665 96660 97650
rect 96618 96656 96674 96665
rect 96618 96591 96674 96600
rect 95976 89616 96028 89622
rect 95976 89558 96028 89564
rect 97276 73001 97304 113999
rect 97368 87553 97396 122806
rect 97908 122800 97960 122806
rect 97908 122742 97960 122748
rect 97920 121689 97948 122742
rect 97906 121680 97962 121689
rect 97906 121615 97962 121624
rect 97814 118688 97870 118697
rect 97814 118623 97870 118632
rect 97908 118652 97960 118658
rect 97828 118250 97856 118623
rect 97908 118594 97960 118600
rect 97816 118244 97868 118250
rect 97816 118186 97868 118192
rect 97920 117881 97948 118594
rect 97906 117872 97962 117881
rect 97906 117807 97962 117816
rect 97908 117292 97960 117298
rect 97908 117234 97960 117240
rect 97816 117224 97868 117230
rect 97816 117166 97868 117172
rect 97828 116521 97856 117166
rect 97920 117065 97948 117234
rect 97906 117056 97962 117065
rect 97906 116991 97962 117000
rect 97814 116512 97870 116521
rect 97814 116447 97870 116456
rect 97908 115932 97960 115938
rect 97908 115874 97960 115880
rect 97816 115864 97868 115870
rect 97816 115806 97868 115812
rect 97828 114889 97856 115806
rect 97920 115705 97948 115874
rect 97906 115696 97962 115705
rect 97906 115631 97962 115640
rect 97814 114880 97870 114889
rect 97814 114815 97870 114824
rect 97538 113520 97594 113529
rect 97538 113455 97594 113464
rect 97552 113218 97580 113455
rect 97540 113212 97592 113218
rect 97540 113154 97592 113160
rect 97814 112704 97870 112713
rect 97814 112639 97870 112648
rect 97828 111858 97856 112639
rect 97908 111920 97960 111926
rect 97906 111888 97908 111897
rect 97960 111888 97962 111897
rect 97816 111852 97868 111858
rect 97906 111823 97962 111832
rect 97816 111794 97868 111800
rect 97448 110288 97500 110294
rect 97446 110256 97448 110265
rect 97500 110256 97502 110265
rect 97446 110191 97502 110200
rect 97908 108384 97960 108390
rect 97908 108326 97960 108332
rect 97920 108089 97948 108326
rect 97906 108080 97962 108089
rect 97906 108015 97962 108024
rect 97538 107264 97594 107273
rect 97538 107199 97594 107208
rect 97552 106418 97580 107199
rect 97906 106720 97962 106729
rect 97906 106655 97962 106664
rect 97540 106412 97592 106418
rect 97540 106354 97592 106360
rect 97920 106350 97948 106655
rect 97908 106344 97960 106350
rect 97908 106286 97960 106292
rect 97540 106276 97592 106282
rect 97540 106218 97592 106224
rect 97552 105097 97580 106218
rect 97906 105904 97962 105913
rect 97906 105839 97962 105848
rect 97920 105602 97948 105839
rect 97908 105596 97960 105602
rect 97908 105538 97960 105544
rect 97538 105088 97594 105097
rect 97538 105023 97594 105032
rect 97906 104272 97962 104281
rect 97906 104207 97962 104216
rect 97920 104174 97948 104207
rect 97908 104168 97960 104174
rect 97908 104110 97960 104116
rect 97908 103488 97960 103494
rect 97722 103456 97778 103465
rect 97908 103430 97960 103436
rect 97722 103391 97724 103400
rect 97776 103391 97778 103400
rect 97724 103362 97776 103368
rect 97920 102921 97948 103430
rect 97906 102912 97962 102921
rect 97906 102847 97962 102856
rect 97630 102096 97686 102105
rect 97630 102031 97686 102040
rect 97644 100774 97672 102031
rect 97906 101280 97962 101289
rect 98012 101266 98040 200086
rect 97962 101238 98040 101266
rect 97906 101215 97962 101224
rect 97632 100768 97684 100774
rect 97632 100710 97684 100716
rect 97814 100464 97870 100473
rect 97814 100399 97870 100408
rect 97828 99482 97856 100399
rect 97906 99648 97962 99657
rect 97906 99583 97962 99592
rect 97816 99476 97868 99482
rect 97816 99418 97868 99424
rect 97920 99414 97948 99583
rect 97908 99408 97960 99414
rect 97908 99350 97960 99356
rect 97816 99340 97868 99346
rect 97816 99282 97868 99288
rect 97540 99136 97592 99142
rect 97538 99104 97540 99113
rect 97592 99104 97594 99113
rect 97538 99039 97594 99048
rect 97828 98297 97856 99282
rect 97814 98288 97870 98297
rect 97814 98223 97870 98232
rect 98656 97714 98684 213862
rect 99300 155990 99328 263570
rect 98736 155984 98788 155990
rect 98736 155926 98788 155932
rect 99288 155984 99340 155990
rect 99288 155926 99340 155932
rect 98748 120358 98776 155926
rect 99392 144362 99420 277743
rect 99470 270464 99526 270473
rect 99470 270399 99526 270408
rect 99484 236026 99512 270399
rect 99562 242584 99618 242593
rect 99562 242519 99618 242528
rect 99576 241806 99604 242519
rect 99564 241800 99616 241806
rect 99564 241742 99616 241748
rect 100036 241398 100064 333950
rect 100114 284472 100170 284481
rect 100114 284407 100170 284416
rect 100128 275330 100156 284407
rect 100116 275324 100168 275330
rect 100116 275266 100168 275272
rect 100300 270496 100352 270502
rect 100298 270464 100300 270473
rect 100352 270464 100354 270473
rect 100298 270399 100354 270408
rect 100404 256737 100432 383626
rect 100496 378826 100524 388991
rect 100576 387864 100628 387870
rect 100576 387806 100628 387812
rect 100484 378820 100536 378826
rect 100484 378762 100536 378768
rect 100588 334014 100616 387806
rect 101864 387184 101916 387190
rect 101864 387126 101916 387132
rect 101772 382968 101824 382974
rect 101772 382910 101824 382916
rect 100576 334008 100628 334014
rect 100576 333950 100628 333956
rect 101784 296714 101812 382910
rect 101416 296686 101812 296714
rect 101416 292534 101444 296686
rect 101404 292528 101456 292534
rect 101404 292470 101456 292476
rect 100758 282704 100814 282713
rect 100758 282639 100814 282648
rect 100772 281586 100800 282639
rect 100760 281580 100812 281586
rect 100760 281522 100812 281528
rect 100760 281444 100812 281450
rect 100760 281386 100812 281392
rect 100772 281081 100800 281386
rect 100758 281072 100814 281081
rect 100758 281007 100814 281016
rect 100760 280084 100812 280090
rect 100760 280026 100812 280032
rect 100772 279449 100800 280026
rect 100758 279440 100814 279449
rect 100758 279375 100814 279384
rect 100758 276992 100814 277001
rect 100758 276927 100814 276936
rect 100772 276690 100800 276927
rect 100760 276684 100812 276690
rect 100760 276626 100812 276632
rect 100852 275392 100904 275398
rect 100852 275334 100904 275340
rect 100760 274644 100812 274650
rect 100760 274586 100812 274592
rect 100772 273737 100800 274586
rect 100864 274553 100892 275334
rect 100850 274544 100906 274553
rect 100850 274479 100906 274488
rect 100758 273728 100814 273737
rect 100758 273663 100814 273672
rect 100760 273216 100812 273222
rect 100760 273158 100812 273164
rect 100772 272921 100800 273158
rect 100758 272912 100814 272921
rect 100758 272847 100814 272856
rect 101126 272096 101182 272105
rect 101126 272031 101128 272040
rect 101180 272031 101182 272040
rect 101128 272002 101180 272008
rect 100758 268832 100814 268841
rect 100758 268767 100814 268776
rect 100772 268394 100800 268767
rect 101220 268456 101272 268462
rect 101220 268398 101272 268404
rect 100760 268388 100812 268394
rect 100760 268330 100812 268336
rect 101232 268025 101260 268398
rect 101218 268016 101274 268025
rect 101218 267951 101274 267960
rect 100760 267708 100812 267714
rect 100760 267650 100812 267656
rect 100772 267209 100800 267650
rect 100758 267200 100814 267209
rect 100758 267135 100814 267144
rect 100852 266348 100904 266354
rect 100852 266290 100904 266296
rect 100864 265577 100892 266290
rect 100850 265568 100906 265577
rect 100850 265503 100906 265512
rect 100760 264920 100812 264926
rect 100760 264862 100812 264868
rect 100772 263945 100800 264862
rect 100758 263936 100814 263945
rect 100758 263871 100814 263880
rect 101232 263634 101260 267951
rect 101220 263628 101272 263634
rect 101220 263570 101272 263576
rect 100758 262304 100814 262313
rect 100758 262239 100760 262248
rect 100812 262239 100814 262248
rect 100760 262210 100812 262216
rect 101416 261497 101444 292470
rect 101876 291961 101904 387126
rect 101956 373312 102008 373318
rect 101956 373254 102008 373260
rect 101862 291952 101918 291961
rect 101862 291887 101918 291896
rect 101496 291848 101548 291854
rect 101496 291790 101548 291796
rect 101508 280265 101536 291790
rect 101494 280256 101550 280265
rect 101494 280191 101550 280200
rect 101968 277394 101996 373254
rect 102060 278730 102088 389778
rect 102244 388550 102272 390374
rect 102428 389174 102456 390895
rect 103886 390688 103942 390697
rect 103942 390646 104144 390674
rect 103886 390623 103942 390632
rect 102336 389146 102456 389174
rect 102520 390374 102856 390402
rect 102232 388544 102284 388550
rect 102232 388486 102284 388492
rect 102336 378282 102364 389146
rect 102520 387870 102548 390374
rect 103578 390130 103606 390388
rect 104880 390374 105216 390402
rect 103532 390102 103606 390130
rect 102508 387864 102560 387870
rect 102508 387806 102560 387812
rect 102782 387832 102838 387841
rect 102782 387767 102838 387776
rect 102324 378276 102376 378282
rect 102324 378218 102376 378224
rect 102140 369164 102192 369170
rect 102140 369106 102192 369112
rect 102048 278724 102100 278730
rect 102048 278666 102100 278672
rect 101876 277366 101996 277394
rect 101876 272066 101904 277366
rect 101864 272060 101916 272066
rect 101864 272002 101916 272008
rect 101680 263560 101732 263566
rect 101680 263502 101732 263508
rect 101692 263129 101720 263502
rect 101678 263120 101734 263129
rect 101678 263055 101734 263064
rect 100942 261488 100998 261497
rect 100942 261423 100998 261432
rect 101402 261488 101458 261497
rect 101402 261423 101458 261432
rect 100760 260840 100812 260846
rect 100760 260782 100812 260788
rect 100772 260681 100800 260782
rect 100758 260672 100814 260681
rect 100758 260607 100814 260616
rect 100760 259412 100812 259418
rect 100760 259354 100812 259360
rect 100772 259049 100800 259354
rect 100758 259040 100814 259049
rect 100758 258975 100814 258984
rect 100760 258256 100812 258262
rect 100758 258224 100760 258233
rect 100812 258224 100814 258233
rect 100758 258159 100814 258168
rect 100772 258074 100800 258159
rect 100680 258046 100800 258074
rect 100390 256728 100446 256737
rect 100390 256663 100446 256672
rect 100114 242584 100170 242593
rect 100114 242519 100170 242528
rect 100128 241777 100156 242519
rect 100114 241768 100170 241777
rect 100114 241703 100170 241712
rect 100024 241392 100076 241398
rect 100024 241334 100076 241340
rect 99472 236020 99524 236026
rect 99472 235962 99524 235968
rect 100022 234560 100078 234569
rect 100022 234495 100078 234504
rect 99380 144356 99432 144362
rect 99380 144298 99432 144304
rect 98736 120352 98788 120358
rect 98736 120294 98788 120300
rect 98736 118992 98788 118998
rect 98736 118934 98788 118940
rect 98644 97708 98696 97714
rect 98644 97650 98696 97656
rect 97906 97472 97962 97481
rect 97906 97407 97962 97416
rect 97920 96694 97948 97407
rect 97908 96688 97960 96694
rect 97908 96630 97960 96636
rect 97448 95940 97500 95946
rect 97448 95882 97500 95888
rect 97354 87544 97410 87553
rect 97354 87479 97410 87488
rect 97460 85474 97488 95882
rect 97906 95296 97962 95305
rect 97906 95231 97908 95240
rect 97960 95231 97962 95240
rect 97908 95202 97960 95208
rect 97816 95192 97868 95198
rect 97816 95134 97868 95140
rect 97828 94489 97856 95134
rect 97814 94480 97870 94489
rect 97814 94415 97870 94424
rect 98748 92313 98776 118934
rect 98828 101448 98880 101454
rect 98828 101390 98880 101396
rect 98734 92304 98790 92313
rect 98734 92239 98790 92248
rect 97448 85468 97500 85474
rect 97448 85410 97500 85416
rect 98840 80073 98868 101390
rect 100036 99142 100064 234495
rect 100680 147694 100708 258046
rect 100760 257440 100812 257446
rect 100758 257408 100760 257417
rect 100812 257408 100814 257417
rect 100758 257343 100814 257352
rect 100850 254960 100906 254969
rect 100850 254895 100906 254904
rect 100760 254584 100812 254590
rect 100760 254526 100812 254532
rect 100772 254153 100800 254526
rect 100758 254144 100814 254153
rect 100758 254079 100814 254088
rect 100864 253978 100892 254895
rect 100852 253972 100904 253978
rect 100852 253914 100904 253920
rect 100760 253904 100812 253910
rect 100760 253846 100812 253852
rect 100772 253337 100800 253846
rect 100758 253328 100814 253337
rect 100758 253263 100814 253272
rect 100852 253224 100904 253230
rect 100852 253166 100904 253172
rect 100864 252521 100892 253166
rect 100850 252512 100906 252521
rect 100850 252447 100906 252456
rect 100758 250880 100814 250889
rect 100758 250815 100814 250824
rect 100772 249830 100800 250815
rect 100760 249824 100812 249830
rect 100760 249766 100812 249772
rect 100760 249688 100812 249694
rect 100760 249630 100812 249636
rect 100116 147688 100168 147694
rect 100116 147630 100168 147636
rect 100668 147688 100720 147694
rect 100668 147630 100720 147636
rect 100128 111110 100156 147630
rect 100208 139460 100260 139466
rect 100208 139402 100260 139408
rect 100220 128314 100248 139402
rect 100208 128308 100260 128314
rect 100208 128250 100260 128256
rect 100116 111104 100168 111110
rect 100116 111046 100168 111052
rect 100772 110294 100800 249630
rect 100760 110288 100812 110294
rect 100760 110230 100812 110236
rect 100864 105602 100892 252447
rect 100956 118726 100984 261423
rect 101220 259888 101272 259894
rect 101218 259856 101220 259865
rect 101272 259856 101274 259865
rect 101218 259791 101274 259800
rect 101128 257440 101180 257446
rect 101128 257382 101180 257388
rect 101036 256692 101088 256698
rect 101036 256634 101088 256640
rect 101048 255785 101076 256634
rect 101034 255776 101090 255785
rect 101034 255711 101090 255720
rect 101140 249694 101168 257382
rect 101956 250504 102008 250510
rect 101956 250446 102008 250452
rect 101968 250073 101996 250446
rect 101954 250064 102010 250073
rect 101954 249999 102010 250008
rect 101128 249688 101180 249694
rect 101128 249630 101180 249636
rect 101680 249076 101732 249082
rect 101680 249018 101732 249024
rect 101692 248441 101720 249018
rect 101678 248432 101734 248441
rect 101968 248414 101996 249999
rect 101968 248386 102088 248414
rect 101678 248367 101734 248376
rect 101128 247036 101180 247042
rect 101128 246978 101180 246984
rect 101034 246800 101090 246809
rect 101034 246735 101090 246744
rect 101048 246362 101076 246735
rect 101036 246356 101088 246362
rect 101036 246298 101088 246304
rect 101140 245993 101168 246978
rect 101126 245984 101182 245993
rect 101126 245919 101182 245928
rect 101034 242720 101090 242729
rect 101034 242655 101090 242664
rect 101048 241738 101076 242655
rect 101036 241732 101088 241738
rect 101036 241674 101088 241680
rect 102060 137902 102088 248386
rect 102152 235890 102180 369106
rect 102796 284209 102824 387767
rect 103532 327078 103560 390102
rect 104164 388476 104216 388482
rect 104164 388418 104216 388424
rect 103520 327072 103572 327078
rect 103520 327014 103572 327020
rect 103426 318336 103482 318345
rect 103426 318271 103482 318280
rect 102782 284200 102838 284209
rect 102782 284135 102838 284144
rect 102232 279472 102284 279478
rect 102232 279414 102284 279420
rect 102244 276185 102272 279414
rect 102230 276176 102286 276185
rect 102230 276111 102286 276120
rect 102782 268560 102838 268569
rect 102782 268495 102838 268504
rect 102796 259894 102824 268495
rect 103440 263566 103468 318271
rect 104176 310486 104204 388418
rect 105188 384334 105216 390374
rect 105280 390374 105616 390402
rect 105280 389065 105308 390374
rect 106338 390130 106366 390388
rect 106292 390102 106366 390130
rect 105266 389056 105322 389065
rect 105266 388991 105322 389000
rect 105544 388476 105596 388482
rect 105544 388418 105596 388424
rect 105176 384328 105228 384334
rect 105176 384270 105228 384276
rect 104808 328772 104860 328778
rect 104808 328714 104860 328720
rect 104164 310480 104216 310486
rect 104164 310422 104216 310428
rect 103612 301504 103664 301510
rect 103612 301446 103664 301452
rect 103520 289944 103572 289950
rect 103520 289886 103572 289892
rect 103428 263560 103480 263566
rect 103428 263502 103480 263508
rect 103428 261588 103480 261594
rect 103428 261530 103480 261536
rect 102784 259888 102836 259894
rect 102784 259830 102836 259836
rect 102414 245712 102470 245721
rect 102414 245647 102470 245656
rect 102322 245168 102378 245177
rect 102322 245103 102378 245112
rect 102232 244928 102284 244934
rect 102232 244870 102284 244876
rect 102244 243545 102272 244870
rect 102230 243536 102286 243545
rect 102230 243471 102286 243480
rect 102336 238754 102364 245103
rect 102428 244361 102456 245647
rect 102414 244352 102470 244361
rect 102414 244287 102470 244296
rect 102244 238726 102364 238754
rect 102140 235884 102192 235890
rect 102140 235826 102192 235832
rect 102244 234569 102272 238726
rect 102230 234560 102286 234569
rect 102230 234495 102286 234504
rect 102796 229090 102824 259830
rect 103336 251932 103388 251938
rect 103336 251874 103388 251880
rect 103348 249082 103376 251874
rect 103336 249076 103388 249082
rect 103336 249018 103388 249024
rect 103440 245721 103468 261530
rect 103426 245712 103482 245721
rect 103426 245647 103482 245656
rect 103426 241632 103482 241641
rect 103426 241567 103482 241576
rect 103440 241369 103468 241567
rect 103426 241360 103482 241369
rect 103426 241295 103482 241304
rect 103428 236292 103480 236298
rect 103428 236234 103480 236240
rect 102784 229084 102836 229090
rect 102784 229026 102836 229032
rect 102782 162888 102838 162897
rect 102782 162823 102838 162832
rect 102140 152584 102192 152590
rect 102140 152526 102192 152532
rect 101404 137896 101456 137902
rect 101404 137838 101456 137844
rect 102048 137896 102100 137902
rect 102048 137838 102100 137844
rect 100944 118720 100996 118726
rect 100944 118662 100996 118668
rect 100852 105596 100904 105602
rect 100852 105538 100904 105544
rect 101416 103426 101444 137838
rect 101496 106412 101548 106418
rect 101496 106354 101548 106360
rect 101404 103420 101456 103426
rect 101404 103362 101456 103368
rect 100114 102232 100170 102241
rect 100114 102167 100170 102176
rect 99288 99136 99340 99142
rect 99288 99078 99340 99084
rect 100024 99136 100076 99142
rect 100024 99078 100076 99084
rect 99010 96112 99066 96121
rect 99010 96047 99066 96056
rect 99024 92449 99052 96047
rect 99010 92440 99066 92449
rect 99010 92375 99066 92384
rect 99300 80073 99328 99078
rect 100024 97300 100076 97306
rect 100024 97242 100076 97248
rect 100036 86902 100064 97242
rect 100024 86896 100076 86902
rect 100024 86838 100076 86844
rect 98826 80064 98882 80073
rect 98826 79999 98882 80008
rect 99286 80064 99342 80073
rect 99286 79999 99342 80008
rect 100128 77178 100156 102167
rect 101404 98048 101456 98054
rect 101404 97990 101456 97996
rect 100758 91080 100814 91089
rect 100758 91015 100760 91024
rect 100812 91015 100814 91024
rect 100760 90986 100812 90992
rect 101416 89690 101444 97990
rect 101404 89684 101456 89690
rect 101404 89626 101456 89632
rect 100116 77172 100168 77178
rect 100116 77114 100168 77120
rect 101508 75857 101536 106354
rect 102152 84182 102180 152526
rect 102796 133346 102824 162823
rect 103440 159361 103468 236234
rect 103426 159352 103482 159361
rect 103426 159287 103482 159296
rect 103426 156632 103482 156641
rect 103426 156567 103482 156576
rect 102874 139496 102930 139505
rect 102874 139431 102930 139440
rect 102784 133340 102836 133346
rect 102784 133282 102836 133288
rect 102888 120766 102916 139431
rect 102876 120760 102928 120766
rect 102876 120702 102928 120708
rect 102140 84176 102192 84182
rect 102140 84118 102192 84124
rect 101494 75848 101550 75857
rect 101494 75783 101550 75792
rect 97262 72992 97318 73001
rect 97262 72927 97318 72936
rect 95332 71732 95384 71738
rect 95332 71674 95384 71680
rect 93768 71052 93820 71058
rect 93768 70994 93820 71000
rect 93676 64864 93728 64870
rect 93676 64806 93728 64812
rect 90362 61432 90418 61441
rect 90362 61367 90418 61376
rect 90376 6914 90404 61367
rect 91008 21412 91060 21418
rect 91008 21354 91060 21360
rect 90284 6886 90404 6914
rect 89168 3528 89220 3534
rect 89168 3470 89220 3476
rect 89628 3528 89680 3534
rect 89628 3470 89680 3476
rect 89180 480 89208 3470
rect 90284 3466 90312 6886
rect 91020 3534 91048 21354
rect 93780 3534 93808 70994
rect 96528 69692 96580 69698
rect 96528 69634 96580 69640
rect 95146 55856 95202 55865
rect 95146 55791 95202 55800
rect 95056 11756 95108 11762
rect 95056 11698 95108 11704
rect 95068 3534 95096 11698
rect 90364 3528 90416 3534
rect 90364 3470 90416 3476
rect 91008 3528 91060 3534
rect 91008 3470 91060 3476
rect 92756 3528 92808 3534
rect 92756 3470 92808 3476
rect 93768 3528 93820 3534
rect 93768 3470 93820 3476
rect 93952 3528 94004 3534
rect 93952 3470 94004 3476
rect 95056 3528 95108 3534
rect 95056 3470 95108 3476
rect 90272 3460 90324 3466
rect 90272 3402 90324 3408
rect 90376 480 90404 3470
rect 91560 3460 91612 3466
rect 91560 3402 91612 3408
rect 91572 480 91600 3402
rect 92768 480 92796 3470
rect 93964 480 93992 3470
rect 95160 480 95188 55791
rect 96540 6914 96568 69634
rect 97276 7614 97304 72927
rect 99932 66904 99984 66910
rect 99286 66872 99342 66881
rect 99932 66846 99984 66852
rect 99286 66807 99342 66816
rect 97264 7608 97316 7614
rect 97264 7550 97316 7556
rect 97448 7608 97500 7614
rect 97448 7550 97500 7556
rect 96264 6886 96568 6914
rect 96264 480 96292 6886
rect 97460 480 97488 7550
rect 99300 3534 99328 66807
rect 99944 59362 99972 66846
rect 99932 59356 99984 59362
rect 99932 59298 99984 59304
rect 101404 53100 101456 53106
rect 101404 53042 101456 53048
rect 100668 19984 100720 19990
rect 100668 19926 100720 19932
rect 100680 3534 100708 19926
rect 98644 3528 98696 3534
rect 98644 3470 98696 3476
rect 99288 3528 99340 3534
rect 99288 3470 99340 3476
rect 99840 3528 99892 3534
rect 99840 3470 99892 3476
rect 100668 3528 100720 3534
rect 100668 3470 100720 3476
rect 98656 480 98684 3470
rect 99852 480 99880 3470
rect 101034 3360 101090 3369
rect 101034 3295 101090 3304
rect 101048 480 101076 3295
rect 101416 2106 101444 53042
rect 103440 6914 103468 156567
rect 103532 141506 103560 289886
rect 103624 237153 103652 301446
rect 103702 291272 103758 291281
rect 103702 291207 103758 291216
rect 103610 237144 103666 237153
rect 103610 237079 103666 237088
rect 103716 236298 103744 291207
rect 104820 246362 104848 328714
rect 104900 272060 104952 272066
rect 104900 272002 104952 272008
rect 104808 246356 104860 246362
rect 104808 246298 104860 246304
rect 104164 241732 104216 241738
rect 104164 241674 104216 241680
rect 103704 236292 103756 236298
rect 103704 236234 103756 236240
rect 104176 213926 104204 241674
rect 104912 225622 104940 272002
rect 105556 271590 105584 388418
rect 106188 371204 106240 371210
rect 106188 371146 106240 371152
rect 105728 327752 105780 327758
rect 105728 327694 105780 327700
rect 105636 313336 105688 313342
rect 105636 313278 105688 313284
rect 105544 271584 105596 271590
rect 105544 271526 105596 271532
rect 105544 265668 105596 265674
rect 105544 265610 105596 265616
rect 105556 257446 105584 265610
rect 105648 258262 105676 313278
rect 105740 273222 105768 327694
rect 106200 313342 106228 371146
rect 106292 319530 106320 390102
rect 106372 388544 106424 388550
rect 106372 388486 106424 388492
rect 106280 319524 106332 319530
rect 106280 319466 106332 319472
rect 106188 313336 106240 313342
rect 106188 313278 106240 313284
rect 105818 284200 105874 284209
rect 105818 284135 105874 284144
rect 105728 273216 105780 273222
rect 105728 273158 105780 273164
rect 105636 258256 105688 258262
rect 105636 258198 105688 258204
rect 105544 257440 105596 257446
rect 105544 257382 105596 257388
rect 105544 247716 105596 247722
rect 105544 247658 105596 247664
rect 105556 235958 105584 247658
rect 105544 235952 105596 235958
rect 105544 235894 105596 235900
rect 105832 234666 105860 284135
rect 106188 272604 106240 272610
rect 106188 272546 106240 272552
rect 106200 272066 106228 272546
rect 106188 272060 106240 272066
rect 106188 272002 106240 272008
rect 106186 271144 106242 271153
rect 106186 271079 106242 271088
rect 106200 270502 106228 271079
rect 106188 270496 106240 270502
rect 106188 270438 106240 270444
rect 106188 251864 106240 251870
rect 106188 251806 106240 251812
rect 106200 251705 106228 251806
rect 106186 251696 106242 251705
rect 106186 251631 106242 251640
rect 106280 251184 106332 251190
rect 106280 251126 106332 251132
rect 106292 249830 106320 251126
rect 106280 249824 106332 249830
rect 106280 249766 106332 249772
rect 106188 236768 106240 236774
rect 106188 236710 106240 236716
rect 105636 234660 105688 234666
rect 105636 234602 105688 234608
rect 105820 234660 105872 234666
rect 105820 234602 105872 234608
rect 105648 234433 105676 234602
rect 105634 234424 105690 234433
rect 105634 234359 105690 234368
rect 104900 225616 104952 225622
rect 104900 225558 104952 225564
rect 104164 213920 104216 213926
rect 104164 213862 104216 213868
rect 105634 206408 105690 206417
rect 105634 206343 105690 206352
rect 103704 206304 103756 206310
rect 103704 206246 103756 206252
rect 103612 199436 103664 199442
rect 103612 199378 103664 199384
rect 103520 141500 103572 141506
rect 103520 141442 103572 141448
rect 103624 86873 103652 199378
rect 103716 118998 103744 206246
rect 105648 205737 105676 206343
rect 104990 205728 105046 205737
rect 104990 205663 105046 205672
rect 105634 205728 105690 205737
rect 105634 205663 105690 205672
rect 104900 205012 104952 205018
rect 104900 204954 104952 204960
rect 104806 203552 104862 203561
rect 104806 203487 104862 203496
rect 104716 141500 104768 141506
rect 104716 141442 104768 141448
rect 104728 140826 104756 141442
rect 104716 140820 104768 140826
rect 104716 140762 104768 140768
rect 104162 138136 104218 138145
rect 104162 138071 104218 138080
rect 104176 131102 104204 138071
rect 104164 131096 104216 131102
rect 104164 131038 104216 131044
rect 103704 118992 103756 118998
rect 103704 118934 103756 118940
rect 103610 86864 103666 86873
rect 103610 86799 103666 86808
rect 104714 86864 104770 86873
rect 104714 86799 104770 86808
rect 104728 86601 104756 86799
rect 104714 86592 104770 86601
rect 104714 86527 104770 86536
rect 104820 6914 104848 203487
rect 104912 79966 104940 204954
rect 105004 124273 105032 205663
rect 106096 205012 106148 205018
rect 106096 204954 106148 204960
rect 106108 204338 106136 204954
rect 106096 204332 106148 204338
rect 106096 204274 106148 204280
rect 106200 199442 106228 236710
rect 106188 199436 106240 199442
rect 106188 199378 106240 199384
rect 105544 160200 105596 160206
rect 105544 160142 105596 160148
rect 105082 142216 105138 142225
rect 105082 142151 105138 142160
rect 105096 141438 105124 142151
rect 105084 141432 105136 141438
rect 105084 141374 105136 141380
rect 105556 126886 105584 160142
rect 105544 126880 105596 126886
rect 105544 126822 105596 126828
rect 105636 126268 105688 126274
rect 105636 126210 105688 126216
rect 104990 124264 105046 124273
rect 104990 124199 105046 124208
rect 105648 118250 105676 126210
rect 105636 118244 105688 118250
rect 105636 118186 105688 118192
rect 106292 104174 106320 249766
rect 106384 238513 106412 388486
rect 107488 383654 107516 390918
rect 107750 390552 107806 390561
rect 107640 390510 107750 390538
rect 107750 390487 107806 390496
rect 107658 390280 107714 390289
rect 107658 390215 107714 390224
rect 107672 387190 107700 390215
rect 107764 389201 107792 390487
rect 111706 390416 111762 390425
rect 109098 390130 109126 390388
rect 109848 390374 110184 390402
rect 109052 390102 109126 390130
rect 107750 389192 107806 389201
rect 107750 389127 107806 389136
rect 107660 387184 107712 387190
rect 107660 387126 107712 387132
rect 107488 383626 107608 383654
rect 106924 367804 106976 367810
rect 106924 367746 106976 367752
rect 106648 254584 106700 254590
rect 106646 254552 106648 254561
rect 106700 254552 106702 254561
rect 106646 254487 106702 254496
rect 106936 248470 106964 367746
rect 107014 292632 107070 292641
rect 107014 292567 107070 292576
rect 107028 281518 107056 292567
rect 107016 281512 107068 281518
rect 107016 281454 107068 281460
rect 107580 258074 107608 383626
rect 107764 373994 107792 389127
rect 107488 258046 107608 258074
rect 107672 373966 107792 373994
rect 107488 251297 107516 258046
rect 107474 251288 107530 251297
rect 107474 251223 107530 251232
rect 106924 248464 106976 248470
rect 106924 248406 106976 248412
rect 106936 238678 106964 248406
rect 107488 241913 107516 251223
rect 107474 241904 107530 241913
rect 107474 241839 107530 241848
rect 107672 241738 107700 373966
rect 108304 366376 108356 366382
rect 108304 366318 108356 366324
rect 108212 261520 108264 261526
rect 108212 261462 108264 261468
rect 108224 260846 108252 261462
rect 108212 260840 108264 260846
rect 108212 260782 108264 260788
rect 108316 242962 108344 366318
rect 108488 325032 108540 325038
rect 108488 324974 108540 324980
rect 108396 310480 108448 310486
rect 108396 310422 108448 310428
rect 108408 244322 108436 310422
rect 108500 304298 108528 324974
rect 108488 304292 108540 304298
rect 108488 304234 108540 304240
rect 109052 261594 109080 390102
rect 110156 389094 110184 390374
rect 110386 390130 110414 390388
rect 110524 390374 111136 390402
rect 110386 390102 110460 390130
rect 110144 389088 110196 389094
rect 110144 389030 110196 389036
rect 109132 384396 109184 384402
rect 109132 384338 109184 384344
rect 109040 261588 109092 261594
rect 109040 261530 109092 261536
rect 108948 255332 109000 255338
rect 108948 255274 109000 255280
rect 108960 248402 108988 255274
rect 109040 255196 109092 255202
rect 109040 255138 109092 255144
rect 109052 253978 109080 255138
rect 109040 253972 109092 253978
rect 109040 253914 109092 253920
rect 108948 248396 109000 248402
rect 108948 248338 109000 248344
rect 108960 247790 108988 248338
rect 108948 247784 109000 247790
rect 108948 247726 109000 247732
rect 108396 244316 108448 244322
rect 108396 244258 108448 244264
rect 108304 242956 108356 242962
rect 108304 242898 108356 242904
rect 107660 241732 107712 241738
rect 107660 241674 107712 241680
rect 106924 238672 106976 238678
rect 106924 238614 106976 238620
rect 106370 238504 106426 238513
rect 106370 238439 106426 238448
rect 107568 238060 107620 238066
rect 107568 238002 107620 238008
rect 106922 213208 106978 213217
rect 106922 213143 106978 213152
rect 106280 104168 106332 104174
rect 106280 104110 106332 104116
rect 106292 103514 106320 104110
rect 106200 103486 106320 103514
rect 106200 94518 106228 103486
rect 106188 94512 106240 94518
rect 106188 94454 106240 94460
rect 104900 79960 104952 79966
rect 104900 79902 104952 79908
rect 106188 13116 106240 13122
rect 106188 13058 106240 13064
rect 103348 6886 103468 6914
rect 104544 6886 104848 6914
rect 102232 3528 102284 3534
rect 102232 3470 102284 3476
rect 101404 2100 101456 2106
rect 101404 2042 101456 2048
rect 102244 480 102272 3470
rect 103348 480 103376 6886
rect 104544 480 104572 6886
rect 106200 3602 106228 13058
rect 106936 6914 106964 213143
rect 107016 192568 107068 192574
rect 107016 192510 107068 192516
rect 107028 92546 107056 192510
rect 107016 92540 107068 92546
rect 107016 92482 107068 92488
rect 106844 6886 106964 6914
rect 105728 3596 105780 3602
rect 105728 3538 105780 3544
rect 106188 3596 106240 3602
rect 106188 3538 106240 3544
rect 105740 480 105768 3538
rect 106844 3534 106872 6886
rect 107580 3534 107608 238002
rect 108316 234598 108344 242898
rect 108408 238746 108436 244258
rect 108396 238740 108448 238746
rect 108396 238682 108448 238688
rect 108946 236600 109002 236609
rect 108946 236535 109002 236544
rect 108960 236026 108988 236535
rect 108948 236020 109000 236026
rect 108948 235962 109000 235968
rect 108304 234592 108356 234598
rect 108304 234534 108356 234540
rect 108396 231124 108448 231130
rect 108396 231066 108448 231072
rect 108302 229800 108358 229809
rect 108302 229735 108358 229744
rect 107660 200796 107712 200802
rect 107660 200738 107712 200744
rect 107672 108322 107700 200738
rect 107660 108316 107712 108322
rect 107660 108258 107712 108264
rect 107660 92540 107712 92546
rect 107660 92482 107712 92488
rect 107672 82822 107700 92482
rect 107660 82816 107712 82822
rect 107660 82758 107712 82764
rect 108316 3534 108344 229735
rect 108408 90409 108436 231066
rect 108960 202230 108988 235962
rect 108948 202224 109000 202230
rect 108948 202166 109000 202172
rect 108486 154592 108542 154601
rect 108486 154527 108542 154536
rect 108500 118658 108528 154527
rect 108488 118652 108540 118658
rect 108488 118594 108540 118600
rect 109052 108390 109080 253914
rect 109144 236026 109172 384338
rect 109684 311160 109736 311166
rect 109684 311102 109736 311108
rect 109696 251190 109724 311102
rect 110432 253978 110460 390102
rect 110524 328778 110552 390374
rect 111762 390388 111872 390402
rect 111762 390374 111886 390388
rect 111706 390351 111762 390360
rect 111858 390130 111886 390374
rect 112272 390374 112608 390402
rect 111858 390102 111932 390130
rect 111800 387048 111852 387054
rect 111800 386990 111852 386996
rect 110604 360868 110656 360874
rect 110604 360810 110656 360816
rect 110512 328772 110564 328778
rect 110512 328714 110564 328720
rect 110510 288552 110566 288561
rect 110510 288487 110566 288496
rect 110420 253972 110472 253978
rect 110420 253914 110472 253920
rect 109684 251184 109736 251190
rect 109684 251126 109736 251132
rect 109132 236020 109184 236026
rect 109132 235962 109184 235968
rect 110420 195288 110472 195294
rect 110420 195230 110472 195236
rect 109132 180124 109184 180130
rect 109132 180066 109184 180072
rect 109040 108384 109092 108390
rect 109040 108326 109092 108332
rect 109144 90953 109172 180066
rect 109684 108384 109736 108390
rect 109684 108326 109736 108332
rect 109130 90944 109186 90953
rect 109130 90879 109186 90888
rect 108394 90400 108450 90409
rect 108394 90335 108450 90344
rect 108408 81326 108436 90335
rect 108396 81320 108448 81326
rect 108396 81262 108448 81268
rect 109696 77178 109724 108326
rect 110432 85513 110460 195230
rect 110524 177342 110552 288487
rect 110616 238754 110644 360810
rect 110696 327072 110748 327078
rect 110696 327014 110748 327020
rect 110708 325718 110736 327014
rect 110696 325712 110748 325718
rect 110696 325654 110748 325660
rect 110708 242593 110736 325654
rect 111064 253972 111116 253978
rect 111064 253914 111116 253920
rect 111076 247042 111104 253914
rect 111812 251938 111840 386990
rect 111904 255338 111932 390102
rect 112272 387054 112300 390374
rect 112260 387048 112312 387054
rect 112260 386990 112312 386996
rect 112732 382974 112760 405855
rect 112720 382968 112772 382974
rect 112720 382910 112772 382916
rect 113192 373318 113220 419999
rect 113284 389842 113312 427071
rect 113376 424969 113404 442206
rect 113362 424960 113418 424969
rect 113362 424895 113418 424904
rect 113468 416809 113496 579634
rect 115204 558204 115256 558210
rect 115204 558146 115256 558152
rect 115216 442950 115244 558146
rect 115940 550656 115992 550662
rect 115940 550598 115992 550604
rect 115296 443692 115348 443698
rect 115296 443634 115348 443640
rect 115204 442944 115256 442950
rect 115204 442886 115256 442892
rect 114560 440904 114612 440910
rect 114560 440846 114612 440852
rect 113822 430128 113878 430137
rect 113822 430063 113878 430072
rect 113454 416800 113510 416809
rect 113454 416735 113510 416744
rect 113272 389836 113324 389842
rect 113272 389778 113324 389784
rect 113180 373312 113232 373318
rect 113180 373254 113232 373260
rect 112444 363656 112496 363662
rect 112444 363598 112496 363604
rect 111892 255332 111944 255338
rect 111892 255274 111944 255280
rect 111800 251932 111852 251938
rect 111800 251874 111852 251880
rect 111064 247036 111116 247042
rect 111064 246978 111116 246984
rect 110694 242584 110750 242593
rect 110694 242519 110750 242528
rect 112456 241466 112484 363598
rect 113836 325694 113864 430063
rect 114572 421977 114600 440846
rect 114650 437472 114706 437481
rect 114650 437407 114706 437416
rect 114664 424153 114692 437407
rect 114650 424144 114706 424153
rect 114650 424079 114706 424088
rect 114558 421968 114614 421977
rect 114558 421903 114614 421912
rect 114572 421598 114600 421903
rect 114560 421592 114612 421598
rect 114560 421534 114612 421540
rect 114650 418976 114706 418985
rect 114650 418911 114706 418920
rect 114664 402974 114692 418911
rect 115308 414050 115336 443634
rect 115570 432304 115626 432313
rect 115570 432239 115626 432248
rect 115584 432002 115612 432239
rect 115572 431996 115624 432002
rect 115572 431938 115624 431944
rect 115846 431216 115902 431225
rect 115846 431151 115902 431160
rect 115860 430642 115888 431151
rect 115848 430636 115900 430642
rect 115848 430578 115900 430584
rect 115756 430568 115808 430574
rect 115756 430510 115808 430516
rect 115768 429321 115796 430510
rect 115754 429312 115810 429321
rect 115754 429247 115810 429256
rect 115848 429140 115900 429146
rect 115848 429082 115900 429088
rect 115860 428233 115888 429082
rect 115846 428224 115902 428233
rect 115846 428159 115902 428168
rect 115846 426048 115902 426057
rect 115846 425983 115902 425992
rect 115860 425134 115888 425983
rect 115848 425128 115900 425134
rect 115848 425070 115900 425076
rect 115754 424960 115810 424969
rect 115754 424895 115810 424904
rect 115768 423706 115796 424895
rect 115848 424380 115900 424386
rect 115848 424322 115900 424328
rect 115860 424153 115888 424322
rect 115846 424144 115902 424153
rect 115846 424079 115902 424088
rect 115756 423700 115808 423706
rect 115756 423642 115808 423648
rect 115848 423632 115900 423638
rect 115848 423574 115900 423580
rect 115860 423065 115888 423574
rect 115846 423056 115902 423065
rect 115846 422991 115902 423000
rect 115754 420880 115810 420889
rect 115754 420815 115810 420824
rect 115768 419558 115796 420815
rect 115756 419552 115808 419558
rect 115756 419494 115808 419500
rect 115848 416832 115900 416838
rect 115846 416800 115848 416809
rect 115900 416800 115902 416809
rect 115846 416735 115902 416744
rect 115848 415744 115900 415750
rect 115846 415712 115848 415721
rect 115900 415712 115902 415721
rect 115846 415647 115902 415656
rect 115846 414896 115902 414905
rect 115846 414831 115848 414840
rect 115900 414831 115902 414840
rect 115848 414802 115900 414808
rect 115112 414044 115164 414050
rect 115112 413986 115164 413992
rect 115296 414044 115348 414050
rect 115296 413986 115348 413992
rect 115124 412729 115152 413986
rect 115846 413808 115902 413817
rect 115846 413743 115902 413752
rect 115110 412720 115166 412729
rect 115860 412690 115888 413743
rect 115110 412655 115166 412664
rect 115848 412684 115900 412690
rect 115848 412626 115900 412632
rect 115204 411936 115256 411942
rect 115204 411878 115256 411884
rect 115216 411641 115244 411878
rect 115202 411632 115258 411641
rect 115202 411567 115258 411576
rect 115848 411256 115900 411262
rect 115848 411198 115900 411204
rect 115860 410553 115888 411198
rect 115846 410544 115902 410553
rect 115846 410479 115902 410488
rect 115848 409828 115900 409834
rect 115848 409770 115900 409776
rect 115860 409737 115888 409770
rect 115846 409728 115902 409737
rect 115846 409663 115902 409672
rect 115018 407552 115074 407561
rect 115018 407487 115020 407496
rect 115072 407487 115074 407496
rect 115020 407458 115072 407464
rect 115848 405680 115900 405686
rect 115846 405648 115848 405657
rect 115900 405648 115902 405657
rect 115846 405583 115902 405592
rect 115848 404592 115900 404598
rect 115846 404560 115848 404569
rect 115900 404560 115902 404569
rect 115846 404495 115902 404504
rect 115846 403472 115902 403481
rect 115846 403407 115902 403416
rect 115860 403034 115888 403407
rect 115848 403028 115900 403034
rect 114664 402946 114784 402974
rect 115848 402970 115900 402976
rect 114558 399528 114614 399537
rect 114558 399463 114614 399472
rect 114572 398857 114600 399463
rect 114558 398848 114614 398857
rect 114558 398783 114614 398792
rect 114572 396409 114600 398783
rect 114558 396400 114614 396409
rect 114558 396335 114614 396344
rect 114558 392048 114614 392057
rect 114558 391983 114614 391992
rect 114008 325780 114060 325786
rect 114008 325722 114060 325728
rect 114020 325694 114048 325722
rect 113836 325666 114048 325694
rect 113824 323604 113876 323610
rect 113824 323546 113876 323552
rect 112536 288516 112588 288522
rect 112536 288458 112588 288464
rect 112444 241460 112496 241466
rect 112444 241402 112496 241408
rect 110616 238726 110736 238754
rect 110708 231810 110736 238726
rect 111708 236700 111760 236706
rect 111708 236642 111760 236648
rect 110696 231804 110748 231810
rect 110696 231746 110748 231752
rect 110708 231130 110736 231746
rect 110696 231124 110748 231130
rect 110696 231066 110748 231072
rect 111614 216064 111670 216073
rect 111614 215999 111670 216008
rect 110512 177336 110564 177342
rect 110512 177278 110564 177284
rect 110418 85504 110474 85513
rect 110418 85439 110474 85448
rect 109684 77172 109736 77178
rect 109684 77114 109736 77120
rect 106832 3528 106884 3534
rect 106832 3470 106884 3476
rect 106924 3528 106976 3534
rect 106924 3470 106976 3476
rect 107568 3528 107620 3534
rect 107568 3470 107620 3476
rect 108304 3528 108356 3534
rect 110512 3528 110564 3534
rect 108304 3470 108356 3476
rect 109314 3496 109370 3505
rect 106936 480 106964 3470
rect 108120 3460 108172 3466
rect 110512 3470 110564 3476
rect 109314 3431 109370 3440
rect 108120 3402 108172 3408
rect 108132 480 108160 3402
rect 109328 480 109356 3431
rect 110524 480 110552 3470
rect 111628 480 111656 215999
rect 111720 3534 111748 236642
rect 112548 222902 112576 288458
rect 113178 287192 113234 287201
rect 113178 287127 113234 287136
rect 112626 245712 112682 245721
rect 112626 245647 112682 245656
rect 112536 222896 112588 222902
rect 112536 222838 112588 222844
rect 112442 220280 112498 220289
rect 112442 220215 112498 220224
rect 112456 220114 112484 220215
rect 112444 220108 112496 220114
rect 112444 220050 112496 220056
rect 112456 89690 112484 220050
rect 112640 200802 112668 245647
rect 113088 225616 113140 225622
rect 113088 225558 113140 225564
rect 112628 200796 112680 200802
rect 112628 200738 112680 200744
rect 112536 147756 112588 147762
rect 112536 147698 112588 147704
rect 112548 119406 112576 147698
rect 112536 119400 112588 119406
rect 112536 119342 112588 119348
rect 111800 89684 111852 89690
rect 111800 89626 111852 89632
rect 112444 89684 112496 89690
rect 112444 89626 112496 89632
rect 111812 89457 111840 89626
rect 111798 89448 111854 89457
rect 111798 89383 111854 89392
rect 113100 6914 113128 225558
rect 113192 153785 113220 287127
rect 113836 268462 113864 323546
rect 113916 304360 113968 304366
rect 113916 304302 113968 304308
rect 113824 268456 113876 268462
rect 113824 268398 113876 268404
rect 113824 257440 113876 257446
rect 113824 257382 113876 257388
rect 113836 244934 113864 257382
rect 113928 255202 113956 304302
rect 114020 291854 114048 325666
rect 114100 304292 114152 304298
rect 114100 304234 114152 304240
rect 114112 294681 114140 304234
rect 114098 294672 114154 294681
rect 114098 294607 114154 294616
rect 114008 291848 114060 291854
rect 114008 291790 114060 291796
rect 113916 255196 113968 255202
rect 113916 255138 113968 255144
rect 114572 250510 114600 391983
rect 114756 388482 114784 402946
rect 115846 402384 115902 402393
rect 115846 402319 115902 402328
rect 115860 402014 115888 402319
rect 115848 402008 115900 402014
rect 115848 401950 115900 401956
rect 115848 401600 115900 401606
rect 115848 401542 115900 401548
rect 115202 401296 115258 401305
rect 115202 401231 115258 401240
rect 115018 391232 115074 391241
rect 115018 391167 115020 391176
rect 115072 391167 115074 391176
rect 115020 391138 115072 391144
rect 114744 388476 114796 388482
rect 114744 388418 114796 388424
rect 115216 335481 115244 401231
rect 115860 400489 115888 401542
rect 115846 400480 115902 400489
rect 115846 400415 115902 400424
rect 115386 399392 115442 399401
rect 115386 399327 115442 399336
rect 115400 399226 115428 399327
rect 115388 399220 115440 399226
rect 115388 399162 115440 399168
rect 115570 398304 115626 398313
rect 115570 398239 115626 398248
rect 115584 397526 115612 398239
rect 115572 397520 115624 397526
rect 115572 397462 115624 397468
rect 115846 397216 115902 397225
rect 115846 397151 115902 397160
rect 115860 396098 115888 397151
rect 115848 396092 115900 396098
rect 115848 396034 115900 396040
rect 115846 395312 115902 395321
rect 115846 395247 115902 395256
rect 115860 394738 115888 395247
rect 115848 394732 115900 394738
rect 115848 394674 115900 394680
rect 115386 394224 115442 394233
rect 115386 394159 115442 394168
rect 115202 335472 115258 335481
rect 115202 335407 115258 335416
rect 115216 335354 115244 335407
rect 115216 335326 115336 335354
rect 115204 331356 115256 331362
rect 115204 331298 115256 331304
rect 115216 251870 115244 331298
rect 115308 265674 115336 335326
rect 115400 331362 115428 394159
rect 115848 393304 115900 393310
rect 115848 393246 115900 393252
rect 115860 393145 115888 393246
rect 115846 393136 115902 393145
rect 115846 393071 115902 393080
rect 115952 386374 115980 550598
rect 116596 536761 116624 702714
rect 118700 576972 118752 576978
rect 118700 576914 118752 576920
rect 116582 536752 116638 536761
rect 116582 536687 116638 536696
rect 117320 529236 117372 529242
rect 117320 529178 117372 529184
rect 116124 472660 116176 472666
rect 116124 472602 116176 472608
rect 116032 444440 116084 444446
rect 116032 444382 116084 444388
rect 115940 386368 115992 386374
rect 115940 386310 115992 386316
rect 115940 380112 115992 380118
rect 115940 380054 115992 380060
rect 115388 331356 115440 331362
rect 115388 331298 115440 331304
rect 115952 268666 115980 380054
rect 116044 318209 116072 444382
rect 116136 411942 116164 472602
rect 116216 416764 116268 416770
rect 116216 416706 116268 416712
rect 116228 415750 116256 416706
rect 116216 415744 116268 415750
rect 116216 415686 116268 415692
rect 116124 411936 116176 411942
rect 116124 411878 116176 411884
rect 116228 380866 116256 415686
rect 117332 414866 117360 529178
rect 117504 449200 117556 449206
rect 117504 449142 117556 449148
rect 117412 434784 117464 434790
rect 117412 434726 117464 434732
rect 117320 414860 117372 414866
rect 117320 414802 117372 414808
rect 117320 405612 117372 405618
rect 117320 405554 117372 405560
rect 117332 404598 117360 405554
rect 117320 404592 117372 404598
rect 117320 404534 117372 404540
rect 117332 384305 117360 404534
rect 117318 384296 117374 384305
rect 117318 384231 117374 384240
rect 117320 381540 117372 381546
rect 117320 381482 117372 381488
rect 116216 380860 116268 380866
rect 116216 380802 116268 380808
rect 116228 380118 116256 380802
rect 116216 380112 116268 380118
rect 116216 380054 116268 380060
rect 116582 318336 116638 318345
rect 116582 318271 116638 318280
rect 116030 318200 116086 318209
rect 116030 318135 116086 318144
rect 116596 317490 116624 318271
rect 116584 317484 116636 317490
rect 116584 317426 116636 317432
rect 115940 268660 115992 268666
rect 115940 268602 115992 268608
rect 115952 268394 115980 268602
rect 115940 268388 115992 268394
rect 115940 268330 115992 268336
rect 115296 265668 115348 265674
rect 115296 265610 115348 265616
rect 115296 264240 115348 264246
rect 115296 264182 115348 264188
rect 115204 251864 115256 251870
rect 115204 251806 115256 251812
rect 114560 250504 114612 250510
rect 114560 250446 114612 250452
rect 113824 244928 113876 244934
rect 113824 244870 113876 244876
rect 115308 243545 115336 264182
rect 115388 249824 115440 249830
rect 115388 249766 115440 249772
rect 115294 243536 115350 243545
rect 115294 243471 115350 243480
rect 115202 241632 115258 241641
rect 115202 241567 115258 241576
rect 115216 228993 115244 241567
rect 115400 238649 115428 249766
rect 115386 238640 115442 238649
rect 115386 238575 115442 238584
rect 115940 234660 115992 234666
rect 115940 234602 115992 234608
rect 115202 228984 115258 228993
rect 115202 228919 115258 228928
rect 115754 225040 115810 225049
rect 115754 224975 115810 224984
rect 113272 218748 113324 218754
rect 113272 218690 113324 218696
rect 113284 218074 113312 218690
rect 113272 218068 113324 218074
rect 113272 218010 113324 218016
rect 113178 153776 113234 153785
rect 113178 153711 113234 153720
rect 113284 88097 113312 218010
rect 114560 211812 114612 211818
rect 114560 211754 114612 211760
rect 114572 211206 114600 211754
rect 114560 211200 114612 211206
rect 114560 211142 114612 211148
rect 114468 145580 114520 145586
rect 114468 145522 114520 145528
rect 113270 88088 113326 88097
rect 113270 88023 113326 88032
rect 112824 6886 113128 6914
rect 111708 3528 111760 3534
rect 111708 3470 111760 3476
rect 112824 480 112852 6886
rect 114480 3466 114508 145522
rect 114572 95198 114600 211142
rect 115768 150521 115796 224975
rect 115846 220144 115902 220153
rect 115846 220079 115902 220088
rect 115202 150512 115258 150521
rect 115202 150447 115258 150456
rect 115754 150512 115810 150521
rect 115754 150447 115810 150456
rect 115216 129674 115244 150447
rect 115204 129668 115256 129674
rect 115204 129610 115256 129616
rect 114560 95192 114612 95198
rect 114560 95134 114612 95140
rect 115860 3466 115888 220079
rect 115952 66162 115980 234602
rect 116596 146985 116624 317426
rect 117228 294092 117280 294098
rect 117228 294034 117280 294040
rect 116676 268660 116728 268666
rect 116676 268602 116728 268608
rect 116688 240786 116716 268602
rect 117240 249121 117268 294034
rect 117226 249112 117282 249121
rect 117226 249047 117282 249056
rect 117332 247722 117360 381482
rect 117424 316810 117452 434726
rect 117516 405618 117544 449142
rect 117596 432064 117648 432070
rect 117596 432006 117648 432012
rect 117608 407114 117636 432006
rect 117596 407108 117648 407114
rect 117596 407050 117648 407056
rect 117504 405612 117556 405618
rect 117504 405554 117556 405560
rect 117504 399220 117556 399226
rect 117504 399162 117556 399168
rect 117516 396778 117544 399162
rect 117504 396772 117556 396778
rect 117504 396714 117556 396720
rect 118712 389842 118740 576914
rect 119356 536790 119384 703122
rect 124220 589960 124272 589966
rect 124220 589902 124272 589908
rect 121736 585812 121788 585818
rect 121736 585754 121788 585760
rect 121748 585206 121776 585754
rect 121460 585200 121512 585206
rect 121460 585142 121512 585148
rect 121736 585200 121788 585206
rect 121736 585142 121788 585148
rect 120080 574796 120132 574802
rect 120080 574738 120132 574744
rect 119344 536784 119396 536790
rect 119344 536726 119396 536732
rect 118792 482316 118844 482322
rect 118792 482258 118844 482264
rect 118804 429146 118832 482258
rect 118884 446480 118936 446486
rect 118884 446422 118936 446428
rect 118792 429140 118844 429146
rect 118792 429082 118844 429088
rect 118792 426420 118844 426426
rect 118792 426362 118844 426368
rect 118804 425134 118832 426362
rect 118792 425128 118844 425134
rect 118792 425070 118844 425076
rect 118700 389836 118752 389842
rect 118700 389778 118752 389784
rect 118712 389230 118740 389778
rect 118700 389224 118752 389230
rect 118700 389166 118752 389172
rect 118700 377528 118752 377534
rect 118700 377470 118752 377476
rect 117412 316804 117464 316810
rect 117412 316746 117464 316752
rect 117412 309800 117464 309806
rect 117412 309742 117464 309748
rect 117320 247716 117372 247722
rect 117320 247658 117372 247664
rect 116676 240780 116728 240786
rect 116676 240722 116728 240728
rect 117320 222896 117372 222902
rect 117320 222838 117372 222844
rect 117226 214568 117282 214577
rect 117226 214503 117282 214512
rect 116674 153232 116730 153241
rect 116674 153167 116730 153176
rect 116582 146976 116638 146985
rect 116582 146911 116638 146920
rect 116688 122806 116716 153167
rect 116676 122800 116728 122806
rect 116676 122742 116728 122748
rect 116584 109744 116636 109750
rect 116584 109686 116636 109692
rect 116596 85542 116624 109686
rect 116584 85536 116636 85542
rect 116584 85478 116636 85484
rect 115940 66156 115992 66162
rect 115940 66098 115992 66104
rect 117240 3466 117268 214503
rect 117332 164966 117360 222838
rect 117424 215286 117452 309742
rect 117962 302560 118018 302569
rect 117962 302495 118018 302504
rect 117976 263566 118004 302495
rect 117964 263560 118016 263566
rect 117964 263502 118016 263508
rect 118712 233238 118740 377470
rect 118804 276690 118832 425070
rect 118896 391270 118924 446422
rect 118976 434036 119028 434042
rect 118976 433978 119028 433984
rect 118988 416770 119016 433978
rect 118976 416764 119028 416770
rect 118976 416706 119028 416712
rect 118976 402008 119028 402014
rect 118976 401950 119028 401956
rect 118884 391264 118936 391270
rect 118884 391206 118936 391212
rect 118896 390998 118924 391206
rect 118884 390992 118936 390998
rect 118884 390934 118936 390940
rect 118988 371210 119016 401950
rect 120092 383654 120120 574738
rect 120172 463004 120224 463010
rect 120172 462946 120224 462952
rect 120184 402014 120212 462946
rect 120264 442944 120316 442950
rect 120264 442886 120316 442892
rect 120276 409834 120304 442886
rect 120264 409828 120316 409834
rect 120264 409770 120316 409776
rect 120276 409154 120304 409770
rect 120264 409148 120316 409154
rect 120264 409090 120316 409096
rect 120172 402008 120224 402014
rect 120172 401950 120224 401956
rect 120172 391196 120224 391202
rect 120172 391138 120224 391144
rect 120080 383648 120132 383654
rect 120080 383590 120132 383596
rect 120092 382294 120120 383590
rect 120080 382288 120132 382294
rect 120080 382230 120132 382236
rect 118976 371204 119028 371210
rect 118976 371146 119028 371152
rect 119986 312216 120042 312225
rect 119986 312151 120042 312160
rect 118792 276684 118844 276690
rect 118792 276626 118844 276632
rect 118700 233232 118752 233238
rect 118698 233200 118700 233209
rect 118752 233200 118754 233209
rect 118698 233135 118754 233144
rect 118804 226273 118832 276626
rect 119344 233232 119396 233238
rect 119344 233174 119396 233180
rect 119356 232558 119384 233174
rect 119344 232552 119396 232558
rect 119344 232494 119396 232500
rect 118790 226264 118846 226273
rect 118790 226199 118846 226208
rect 118804 225049 118832 226199
rect 118790 225040 118846 225049
rect 118790 224975 118846 224984
rect 117412 215280 117464 215286
rect 117412 215222 117464 215228
rect 117424 214810 117452 215222
rect 117412 214804 117464 214810
rect 117412 214746 117464 214752
rect 118700 202224 118752 202230
rect 118700 202166 118752 202172
rect 117962 167240 118018 167249
rect 117962 167175 118018 167184
rect 117320 164960 117372 164966
rect 117320 164902 117372 164908
rect 117976 144129 118004 167175
rect 118056 150544 118108 150550
rect 118056 150486 118108 150492
rect 117962 144120 118018 144129
rect 117962 144055 118018 144064
rect 118068 129062 118096 150486
rect 118606 144120 118662 144129
rect 118606 144055 118662 144064
rect 118056 129056 118108 129062
rect 118056 128998 118108 129004
rect 118620 3466 118648 144055
rect 118712 57866 118740 202166
rect 119356 86737 119384 232494
rect 119342 86728 119398 86737
rect 119342 86663 119398 86672
rect 118700 57860 118752 57866
rect 118700 57802 118752 57808
rect 120000 6914 120028 312151
rect 120184 295322 120212 391138
rect 121472 387802 121500 585142
rect 122840 583772 122892 583778
rect 122840 583714 122892 583720
rect 121552 555484 121604 555490
rect 121552 555426 121604 555432
rect 121564 412690 121592 555426
rect 122196 438184 122248 438190
rect 122196 438126 122248 438132
rect 122208 437510 122236 438126
rect 122196 437504 122248 437510
rect 122196 437446 122248 437452
rect 122208 431954 122236 437446
rect 122116 431926 122236 431954
rect 121644 414860 121696 414866
rect 121644 414802 121696 414808
rect 121552 412684 121604 412690
rect 121552 412626 121604 412632
rect 121552 407516 121604 407522
rect 121552 407458 121604 407464
rect 120724 387796 120776 387802
rect 120724 387738 120776 387744
rect 121460 387796 121512 387802
rect 121460 387738 121512 387744
rect 120736 387122 120764 387738
rect 120724 387116 120776 387122
rect 120724 387058 120776 387064
rect 120172 295316 120224 295322
rect 120172 295258 120224 295264
rect 120184 294098 120212 295258
rect 120172 294092 120224 294098
rect 120172 294034 120224 294040
rect 120080 251864 120132 251870
rect 120080 251806 120132 251812
rect 120092 106282 120120 251806
rect 120736 220289 120764 387058
rect 121458 312080 121514 312089
rect 121458 312015 121514 312024
rect 121368 262676 121420 262682
rect 121368 262618 121420 262624
rect 121380 262274 121408 262618
rect 121368 262268 121420 262274
rect 121368 262210 121420 262216
rect 121380 254590 121408 262210
rect 121368 254584 121420 254590
rect 121368 254526 121420 254532
rect 121472 236774 121500 312015
rect 121564 262682 121592 407458
rect 121656 323610 121684 414802
rect 121644 323604 121696 323610
rect 121644 323546 121696 323552
rect 122116 318345 122144 431926
rect 122852 426426 122880 583714
rect 122932 485104 122984 485110
rect 122932 485046 122984 485052
rect 122840 426420 122892 426426
rect 122840 426362 122892 426368
rect 122944 423638 122972 485046
rect 123116 453348 123168 453354
rect 123116 453290 123168 453296
rect 123024 436212 123076 436218
rect 123024 436154 123076 436160
rect 122932 423632 122984 423638
rect 122932 423574 122984 423580
rect 122932 412684 122984 412690
rect 122932 412626 122984 412632
rect 122840 382288 122892 382294
rect 122840 382230 122892 382236
rect 122102 318336 122158 318345
rect 122102 318271 122158 318280
rect 122748 309188 122800 309194
rect 122748 309130 122800 309136
rect 122104 292596 122156 292602
rect 122104 292538 122156 292544
rect 122116 278730 122144 292538
rect 122104 278724 122156 278730
rect 122104 278666 122156 278672
rect 121552 262676 121604 262682
rect 121552 262618 121604 262624
rect 121460 236768 121512 236774
rect 121460 236710 121512 236716
rect 122656 227044 122708 227050
rect 122656 226986 122708 226992
rect 120722 220280 120778 220289
rect 120722 220215 120778 220224
rect 120172 214804 120224 214810
rect 120172 214746 120224 214752
rect 120080 106276 120132 106282
rect 120080 106218 120132 106224
rect 120184 88097 120212 214746
rect 122668 88233 122696 226986
rect 122102 88224 122158 88233
rect 122102 88159 122158 88168
rect 122654 88224 122710 88233
rect 122654 88159 122710 88168
rect 120170 88088 120226 88097
rect 120170 88023 120226 88032
rect 122116 82754 122144 88159
rect 122104 82748 122156 82754
rect 122104 82690 122156 82696
rect 121368 22772 121420 22778
rect 121368 22714 121420 22720
rect 121380 6914 121408 22714
rect 119908 6886 120028 6914
rect 121104 6886 121408 6914
rect 114008 3460 114060 3466
rect 114008 3402 114060 3408
rect 114468 3460 114520 3466
rect 114468 3402 114520 3408
rect 115204 3460 115256 3466
rect 115204 3402 115256 3408
rect 115848 3460 115900 3466
rect 115848 3402 115900 3408
rect 116400 3460 116452 3466
rect 116400 3402 116452 3408
rect 117228 3460 117280 3466
rect 117228 3402 117280 3408
rect 117596 3460 117648 3466
rect 117596 3402 117648 3408
rect 118608 3460 118660 3466
rect 118608 3402 118660 3408
rect 118792 3460 118844 3466
rect 118792 3402 118844 3408
rect 114020 480 114048 3402
rect 115216 480 115244 3402
rect 116412 480 116440 3402
rect 117608 480 117636 3402
rect 118804 480 118832 3402
rect 119908 480 119936 6886
rect 121104 480 121132 6886
rect 122760 3602 122788 309130
rect 122852 235929 122880 382230
rect 122944 267714 122972 412626
rect 123036 320958 123064 436154
rect 123128 422294 123156 453290
rect 124128 423632 124180 423638
rect 124128 423574 124180 423580
rect 124140 422958 124168 423574
rect 124128 422952 124180 422958
rect 124128 422894 124180 422900
rect 123128 422266 123248 422294
rect 123220 411262 123248 422266
rect 123208 411256 123260 411262
rect 123208 411198 123260 411204
rect 124128 411256 124180 411262
rect 124128 411198 124180 411204
rect 124140 410582 124168 411198
rect 124128 410576 124180 410582
rect 124128 410518 124180 410524
rect 124232 397526 124260 589902
rect 132590 582720 132646 582729
rect 132590 582655 132646 582664
rect 130384 578264 130436 578270
rect 130384 578206 130436 578212
rect 128360 576904 128412 576910
rect 128360 576846 128412 576852
rect 128372 527882 128400 576846
rect 128360 527876 128412 527882
rect 128360 527818 128412 527824
rect 124312 443012 124364 443018
rect 124312 442954 124364 442960
rect 124220 397520 124272 397526
rect 124140 397468 124220 397474
rect 124140 397462 124272 397468
rect 124140 397446 124260 397462
rect 124140 343670 124168 397446
rect 123484 343664 123536 343670
rect 123484 343606 123536 343612
rect 124128 343664 124180 343670
rect 124128 343606 124180 343612
rect 123024 320952 123076 320958
rect 123024 320894 123076 320900
rect 123496 304366 123524 343606
rect 124324 316742 124352 442954
rect 127072 439000 127124 439006
rect 127072 438942 127124 438948
rect 125600 437572 125652 437578
rect 125600 437514 125652 437520
rect 124864 429140 124916 429146
rect 124864 429082 124916 429088
rect 124772 389088 124824 389094
rect 124770 389056 124772 389065
rect 124824 389056 124826 389065
rect 124770 388991 124826 389000
rect 124876 340950 124904 429082
rect 124864 340944 124916 340950
rect 124864 340886 124916 340892
rect 125508 340944 125560 340950
rect 125508 340886 125560 340892
rect 125324 320952 125376 320958
rect 125324 320894 125376 320900
rect 125336 320210 125364 320894
rect 125324 320204 125376 320210
rect 125324 320146 125376 320152
rect 124312 316736 124364 316742
rect 124312 316678 124364 316684
rect 125336 316034 125364 320146
rect 125416 316736 125468 316742
rect 125414 316704 125416 316713
rect 125468 316704 125470 316713
rect 125414 316639 125470 316648
rect 125336 316006 125456 316034
rect 124218 307864 124274 307873
rect 124218 307799 124274 307808
rect 123484 304360 123536 304366
rect 123484 304302 123536 304308
rect 124128 295996 124180 296002
rect 124128 295938 124180 295944
rect 124140 293282 124168 295938
rect 124128 293276 124180 293282
rect 124128 293218 124180 293224
rect 124128 272536 124180 272542
rect 124128 272478 124180 272484
rect 122932 267708 122984 267714
rect 122932 267650 122984 267656
rect 122944 266422 122972 267650
rect 122932 266416 122984 266422
rect 122932 266358 122984 266364
rect 122930 243536 122986 243545
rect 122930 243471 122986 243480
rect 122838 235920 122894 235929
rect 122838 235855 122894 235864
rect 122840 199436 122892 199442
rect 122840 199378 122892 199384
rect 122852 85377 122880 199378
rect 122944 169046 122972 243471
rect 123668 169720 123720 169726
rect 123668 169662 123720 169668
rect 123680 169046 123708 169662
rect 122932 169040 122984 169046
rect 122932 168982 122984 168988
rect 123668 169040 123720 169046
rect 123668 168982 123720 168988
rect 124036 85536 124088 85542
rect 124036 85478 124088 85484
rect 124048 85377 124076 85478
rect 122838 85368 122894 85377
rect 122838 85303 122894 85312
rect 124034 85368 124090 85377
rect 124034 85303 124090 85312
rect 124140 3602 124168 272478
rect 124232 233238 124260 307799
rect 124220 233232 124272 233238
rect 124220 233174 124272 233180
rect 125428 149122 125456 316006
rect 125520 304298 125548 340886
rect 125612 325038 125640 437514
rect 126980 423700 127032 423706
rect 126980 423642 127032 423648
rect 126336 403028 126388 403034
rect 126336 402970 126388 402976
rect 125600 325032 125652 325038
rect 125600 324974 125652 324980
rect 125508 304292 125560 304298
rect 125508 304234 125560 304240
rect 126242 276040 126298 276049
rect 126242 275975 126298 275984
rect 125508 238128 125560 238134
rect 125508 238070 125560 238076
rect 125416 149116 125468 149122
rect 125416 149058 125468 149064
rect 125428 144906 125456 149058
rect 125416 144900 125468 144906
rect 125416 144842 125468 144848
rect 125520 3602 125548 238070
rect 125600 204944 125652 204950
rect 125600 204886 125652 204892
rect 125612 92585 125640 204886
rect 125598 92576 125654 92585
rect 125598 92511 125654 92520
rect 125600 33788 125652 33794
rect 125600 33730 125652 33736
rect 125612 16574 125640 33730
rect 126256 22778 126284 275975
rect 126348 262274 126376 402970
rect 126428 300144 126480 300150
rect 126428 300086 126480 300092
rect 126336 262268 126388 262274
rect 126336 262210 126388 262216
rect 126348 259418 126376 262210
rect 126336 259412 126388 259418
rect 126336 259354 126388 259360
rect 126440 253230 126468 300086
rect 126520 294024 126572 294030
rect 126520 293966 126572 293972
rect 126532 269822 126560 293966
rect 126992 280158 127020 423642
rect 127084 321570 127112 438942
rect 128372 393310 128400 527818
rect 128452 490612 128504 490618
rect 128452 490554 128504 490560
rect 128464 401606 128492 490554
rect 129740 487824 129792 487830
rect 129740 487766 129792 487772
rect 128452 401600 128504 401606
rect 128452 401542 128504 401548
rect 128464 400926 128492 401542
rect 128452 400920 128504 400926
rect 128452 400862 128504 400868
rect 128452 397452 128504 397458
rect 128452 397394 128504 397400
rect 128464 396098 128492 397394
rect 128452 396092 128504 396098
rect 128452 396034 128504 396040
rect 128360 393304 128412 393310
rect 128360 393246 128412 393252
rect 128372 392018 128400 393246
rect 128360 392012 128412 392018
rect 128360 391954 128412 391960
rect 128360 389836 128412 389842
rect 128360 389778 128412 389784
rect 127072 321564 127124 321570
rect 127072 321506 127124 321512
rect 127084 320890 127112 321506
rect 127072 320884 127124 320890
rect 127072 320826 127124 320832
rect 127624 287700 127676 287706
rect 127624 287642 127676 287648
rect 127636 287162 127664 287642
rect 127624 287156 127676 287162
rect 127624 287098 127676 287104
rect 126980 280152 127032 280158
rect 126980 280094 127032 280100
rect 127440 280152 127492 280158
rect 127440 280094 127492 280100
rect 127452 279478 127480 280094
rect 127440 279472 127492 279478
rect 127440 279414 127492 279420
rect 126520 269816 126572 269822
rect 126520 269758 126572 269764
rect 126428 253224 126480 253230
rect 126428 253166 126480 253172
rect 126334 249112 126390 249121
rect 126334 249047 126390 249056
rect 126348 201686 126376 249047
rect 126336 201680 126388 201686
rect 126336 201622 126388 201628
rect 127636 146946 127664 287098
rect 127714 282976 127770 282985
rect 127714 282911 127770 282920
rect 127728 241670 127756 282911
rect 127716 241664 127768 241670
rect 127716 241606 127768 241612
rect 128372 227730 128400 389778
rect 128464 262857 128492 396034
rect 129752 386306 129780 487766
rect 129832 419552 129884 419558
rect 129832 419494 129884 419500
rect 129740 386300 129792 386306
rect 129740 386242 129792 386248
rect 128544 380180 128596 380186
rect 128544 380122 128596 380128
rect 128450 262848 128506 262857
rect 128450 262783 128506 262792
rect 128452 246356 128504 246362
rect 128452 246298 128504 246304
rect 128360 227724 128412 227730
rect 128360 227666 128412 227672
rect 128372 227050 128400 227666
rect 128360 227044 128412 227050
rect 128360 226986 128412 226992
rect 127714 149152 127770 149161
rect 127714 149087 127770 149096
rect 127624 146940 127676 146946
rect 127624 146882 127676 146888
rect 127728 133890 127756 149087
rect 127716 133884 127768 133890
rect 127716 133826 127768 133832
rect 128464 103514 128492 246298
rect 128556 239873 128584 380122
rect 129740 378820 129792 378826
rect 129740 378762 129792 378768
rect 129752 258777 129780 378762
rect 129844 327758 129872 419494
rect 130292 386300 130344 386306
rect 130292 386242 130344 386248
rect 130304 385082 130332 386242
rect 130292 385076 130344 385082
rect 130292 385018 130344 385024
rect 129832 327752 129884 327758
rect 129832 327694 129884 327700
rect 129738 258768 129794 258777
rect 129738 258703 129794 258712
rect 128542 239864 128598 239873
rect 128542 239799 128598 239808
rect 129002 229936 129058 229945
rect 129002 229871 129058 229880
rect 128372 103486 128492 103514
rect 128372 99498 128400 103486
rect 128280 99482 128400 99498
rect 128268 99476 128400 99482
rect 128320 99470 128400 99476
rect 128268 99418 128320 99424
rect 128280 71738 128308 99418
rect 128268 71732 128320 71738
rect 128268 71674 128320 71680
rect 126244 22772 126296 22778
rect 126244 22714 126296 22720
rect 125612 16546 125916 16574
rect 122288 3596 122340 3602
rect 122288 3538 122340 3544
rect 122748 3596 122800 3602
rect 122748 3538 122800 3544
rect 123484 3596 123536 3602
rect 123484 3538 123536 3544
rect 124128 3596 124180 3602
rect 124128 3538 124180 3544
rect 124680 3596 124732 3602
rect 124680 3538 124732 3544
rect 125508 3596 125560 3602
rect 125508 3538 125560 3544
rect 122300 480 122328 3538
rect 123496 480 123524 3538
rect 124692 480 124720 3538
rect 125888 480 125916 16546
rect 129016 490 129044 229871
rect 130396 4826 130424 578206
rect 131120 441652 131172 441658
rect 131120 441594 131172 441600
rect 131028 316804 131080 316810
rect 131028 316746 131080 316752
rect 131040 316062 131068 316746
rect 131028 316056 131080 316062
rect 131028 315998 131080 316004
rect 131040 152658 131068 315998
rect 131132 286385 131160 441594
rect 132500 434852 132552 434858
rect 132500 434794 132552 434800
rect 131856 302252 131908 302258
rect 131856 302194 131908 302200
rect 131118 286376 131174 286385
rect 131118 286311 131174 286320
rect 131764 266416 131816 266422
rect 131764 266358 131816 266364
rect 131776 162994 131804 266358
rect 131868 261497 131896 302194
rect 131854 261488 131910 261497
rect 131854 261423 131910 261432
rect 131764 162988 131816 162994
rect 131764 162930 131816 162936
rect 130476 152652 130528 152658
rect 130476 152594 130528 152600
rect 131028 152652 131080 152658
rect 131028 152594 131080 152600
rect 130488 151842 130516 152594
rect 130476 151836 130528 151842
rect 130476 151778 130528 151784
rect 130488 134026 130516 151778
rect 130476 134020 130528 134026
rect 130476 133962 130528 133968
rect 131776 118969 131804 162930
rect 131762 118960 131818 118969
rect 131762 118895 131818 118904
rect 132512 16574 132540 434794
rect 132604 397458 132632 582655
rect 133880 569220 133932 569226
rect 133880 569162 133932 569168
rect 132592 397452 132644 397458
rect 132592 397394 132644 397400
rect 133892 385014 133920 569162
rect 136652 538218 136680 703582
rect 137664 703474 137692 703582
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 137848 703474 137876 703520
rect 137664 703446 137876 703474
rect 154132 703322 154160 703520
rect 154120 703316 154172 703322
rect 154120 703258 154172 703264
rect 170324 703050 170352 703520
rect 170312 703044 170364 703050
rect 170312 702986 170364 702992
rect 202800 702982 202828 703520
rect 218992 703186 219020 703520
rect 235184 703254 235212 703520
rect 264244 703384 264296 703390
rect 264244 703326 264296 703332
rect 235172 703248 235224 703254
rect 235172 703190 235224 703196
rect 218980 703180 219032 703186
rect 218980 703122 219032 703128
rect 202788 702976 202840 702982
rect 202788 702918 202840 702924
rect 140780 586560 140832 586566
rect 140780 586502 140832 586508
rect 136640 538212 136692 538218
rect 136640 538154 136692 538160
rect 136640 533384 136692 533390
rect 136640 533326 136692 533332
rect 133972 431996 134024 432002
rect 133972 431938 134024 431944
rect 133144 385008 133196 385014
rect 133144 384950 133196 384956
rect 133880 385008 133932 385014
rect 133880 384950 133932 384956
rect 133156 384334 133184 384950
rect 133144 384328 133196 384334
rect 133144 384270 133196 384276
rect 133156 204950 133184 384270
rect 133234 299568 133290 299577
rect 133234 299503 133290 299512
rect 133144 204944 133196 204950
rect 133144 204886 133196 204892
rect 133248 201414 133276 299503
rect 133984 281625 134012 431938
rect 135904 430636 135956 430642
rect 135904 430578 135956 430584
rect 134064 392012 134116 392018
rect 134064 391954 134116 391960
rect 134076 311166 134104 391954
rect 134156 385076 134208 385082
rect 134156 385018 134208 385024
rect 134064 311160 134116 311166
rect 134064 311102 134116 311108
rect 133970 281616 134026 281625
rect 133970 281551 134026 281560
rect 134168 206310 134196 385018
rect 135916 288561 135944 430578
rect 136652 430574 136680 533326
rect 137284 438932 137336 438938
rect 137284 438874 137336 438880
rect 136640 430568 136692 430574
rect 136640 430510 136692 430516
rect 136640 410576 136692 410582
rect 136640 410518 136692 410524
rect 135996 304292 136048 304298
rect 135996 304234 136048 304240
rect 135902 288552 135958 288561
rect 135902 288487 135958 288496
rect 134614 284336 134670 284345
rect 134614 284271 134670 284280
rect 134522 280800 134578 280809
rect 134522 280735 134578 280744
rect 134156 206304 134208 206310
rect 134156 206246 134208 206252
rect 133236 201408 133288 201414
rect 133236 201350 133288 201356
rect 132592 200796 132644 200802
rect 132592 200738 132644 200744
rect 132604 99346 132632 200738
rect 132592 99340 132644 99346
rect 132592 99282 132644 99288
rect 133788 99340 133840 99346
rect 133788 99282 133840 99288
rect 133800 98666 133828 99282
rect 133788 98660 133840 98666
rect 133788 98602 133840 98608
rect 132512 16546 133000 16574
rect 130384 4820 130436 4826
rect 130384 4762 130436 4768
rect 129200 598 129412 626
rect 129200 490 129228 598
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129016 462 129228 490
rect 129384 480 129412 598
rect 132972 480 133000 16546
rect 134536 11762 134564 280735
rect 134628 273970 134656 284271
rect 135916 281450 135944 288487
rect 135904 281444 135956 281450
rect 135904 281386 135956 281392
rect 134616 273964 134668 273970
rect 134616 273906 134668 273912
rect 135076 206984 135128 206990
rect 135076 206926 135128 206932
rect 135088 206310 135116 206926
rect 135076 206304 135128 206310
rect 135076 206246 135128 206252
rect 134616 201680 134668 201686
rect 134616 201622 134668 201628
rect 134628 103494 134656 201622
rect 136008 180794 136036 304234
rect 136652 267073 136680 410518
rect 137296 325694 137324 438874
rect 139400 409148 139452 409154
rect 139400 409090 139452 409096
rect 138020 391264 138072 391270
rect 138020 391206 138072 391212
rect 137296 325666 137416 325694
rect 137388 321638 137416 325666
rect 137376 321632 137428 321638
rect 137376 321574 137428 321580
rect 137282 308000 137338 308009
rect 137282 307935 137338 307944
rect 136638 267064 136694 267073
rect 136638 266999 136694 267008
rect 135916 180766 136036 180794
rect 135916 179450 135944 180766
rect 135904 179444 135956 179450
rect 135904 179386 135956 179392
rect 135916 131034 135944 179386
rect 135904 131028 135956 131034
rect 135904 130970 135956 130976
rect 134616 103488 134668 103494
rect 134616 103430 134668 103436
rect 134524 11756 134576 11762
rect 134524 11698 134576 11704
rect 136456 4820 136508 4826
rect 136456 4762 136508 4768
rect 136468 480 136496 4762
rect 137296 3534 137324 307935
rect 137388 287706 137416 321574
rect 137466 289912 137522 289921
rect 137466 289847 137522 289856
rect 137376 287700 137428 287706
rect 137376 287642 137428 287648
rect 137480 257378 137508 289847
rect 138032 257446 138060 391206
rect 138662 281616 138718 281625
rect 138662 281551 138718 281560
rect 138020 257440 138072 257446
rect 138020 257382 138072 257388
rect 137468 257372 137520 257378
rect 137468 257314 137520 257320
rect 138032 257281 138060 257382
rect 138018 257272 138074 257281
rect 138018 257207 138074 257216
rect 137376 256012 137428 256018
rect 137376 255954 137428 255960
rect 137388 53106 137416 255954
rect 138676 224330 138704 281551
rect 139412 264926 139440 409090
rect 140792 405686 140820 586502
rect 140872 436144 140924 436150
rect 140872 436086 140924 436092
rect 140780 405680 140832 405686
rect 140780 405622 140832 405628
rect 140778 398848 140834 398857
rect 140778 398783 140834 398792
rect 140134 304192 140190 304201
rect 140134 304127 140190 304136
rect 140044 265668 140096 265674
rect 140044 265610 140096 265616
rect 139400 264920 139452 264926
rect 139400 264862 139452 264868
rect 138664 224324 138716 224330
rect 138664 224266 138716 224272
rect 138664 202224 138716 202230
rect 138664 202166 138716 202172
rect 137376 53100 137428 53106
rect 137376 53042 137428 53048
rect 138676 42090 138704 202166
rect 138664 42084 138716 42090
rect 138664 42026 138716 42032
rect 140056 36582 140084 265610
rect 140148 228993 140176 304127
rect 140792 253910 140820 398783
rect 140884 277409 140912 436086
rect 142804 430568 142856 430574
rect 142804 430510 142856 430516
rect 142160 411936 142212 411942
rect 142160 411878 142212 411884
rect 141424 405680 141476 405686
rect 141424 405622 141476 405628
rect 141436 404394 141464 405622
rect 141424 404388 141476 404394
rect 141424 404330 141476 404336
rect 141608 302932 141660 302938
rect 141608 302874 141660 302880
rect 140870 277400 140926 277409
rect 140870 277335 140926 277344
rect 140884 276729 140912 277335
rect 140870 276720 140926 276729
rect 140870 276655 140926 276664
rect 141516 271176 141568 271182
rect 141516 271118 141568 271124
rect 141424 262880 141476 262886
rect 141424 262822 141476 262828
rect 140780 253904 140832 253910
rect 140780 253846 140832 253852
rect 141056 253904 141108 253910
rect 141056 253846 141108 253852
rect 141068 253201 141096 253846
rect 141054 253192 141110 253201
rect 141054 253127 141110 253136
rect 140780 249076 140832 249082
rect 140780 249018 140832 249024
rect 140792 246362 140820 249018
rect 140780 246356 140832 246362
rect 140780 246298 140832 246304
rect 140134 228984 140190 228993
rect 140134 228919 140190 228928
rect 140044 36576 140096 36582
rect 140044 36518 140096 36524
rect 141436 13122 141464 262822
rect 141528 50386 141556 271118
rect 141620 256698 141648 302874
rect 142172 266354 142200 411878
rect 142816 320249 142844 430510
rect 144920 424380 144972 424386
rect 144920 424322 144972 424328
rect 143540 416832 143592 416838
rect 143540 416774 143592 416780
rect 142802 320240 142858 320249
rect 142802 320175 142858 320184
rect 142816 316034 142844 320175
rect 142816 316006 142936 316034
rect 142804 303816 142856 303822
rect 142804 303758 142856 303764
rect 142160 266348 142212 266354
rect 142160 266290 142212 266296
rect 141608 256692 141660 256698
rect 141608 256634 141660 256640
rect 141516 50380 141568 50386
rect 141516 50322 141568 50328
rect 141424 13116 141476 13122
rect 141424 13058 141476 13064
rect 141148 7676 141200 7682
rect 141148 7618 141200 7624
rect 141160 3534 141188 7618
rect 142816 7614 142844 303758
rect 142908 280090 142936 316006
rect 142988 288516 143040 288522
rect 142988 288458 143040 288464
rect 142896 280084 142948 280090
rect 142896 280026 142948 280032
rect 143000 272610 143028 288458
rect 142988 272604 143040 272610
rect 142988 272546 143040 272552
rect 143552 269793 143580 416774
rect 143632 404388 143684 404394
rect 143632 404330 143684 404336
rect 143538 269784 143594 269793
rect 143538 269719 143594 269728
rect 142896 267028 142948 267034
rect 142896 266970 142948 266976
rect 142908 28286 142936 266970
rect 143448 266348 143500 266354
rect 143448 266290 143500 266296
rect 143460 265742 143488 266290
rect 143448 265736 143500 265742
rect 143448 265678 143500 265684
rect 143644 261526 143672 404330
rect 144932 274553 144960 424322
rect 148324 422952 148376 422958
rect 148324 422894 148376 422900
rect 146944 421592 146996 421598
rect 146944 421534 146996 421540
rect 146300 400920 146352 400926
rect 146300 400862 146352 400868
rect 145654 284880 145710 284889
rect 145654 284815 145710 284824
rect 144918 274544 144974 274553
rect 144918 274479 144974 274488
rect 145564 268388 145616 268394
rect 145564 268330 145616 268336
rect 144276 264920 144328 264926
rect 144276 264862 144328 264868
rect 143632 261520 143684 261526
rect 143632 261462 143684 261468
rect 144184 260160 144236 260166
rect 144184 260102 144236 260108
rect 142986 157448 143042 157457
rect 142986 157383 143042 157392
rect 143000 132394 143028 157383
rect 142988 132388 143040 132394
rect 142988 132330 143040 132336
rect 144196 44878 144224 260102
rect 144288 242185 144316 264862
rect 144274 242176 144330 242185
rect 144274 242111 144330 242120
rect 144826 202192 144882 202201
rect 144826 202127 144882 202136
rect 144184 44872 144236 44878
rect 144184 44814 144236 44820
rect 142896 28280 142948 28286
rect 142896 28222 142948 28228
rect 142804 7608 142856 7614
rect 142804 7550 142856 7556
rect 144840 3534 144868 202127
rect 145576 29646 145604 268330
rect 145668 215286 145696 284815
rect 146206 274544 146262 274553
rect 146206 274479 146262 274488
rect 146220 273873 146248 274479
rect 146206 273864 146262 273873
rect 146206 273799 146262 273808
rect 146312 255921 146340 400862
rect 146956 299470 146984 421534
rect 147680 414044 147732 414050
rect 147680 413986 147732 413992
rect 146944 299464 146996 299470
rect 146944 299406 146996 299412
rect 146956 274650 146984 299406
rect 146944 274644 146996 274650
rect 146944 274586 146996 274592
rect 146944 272604 146996 272610
rect 146944 272546 146996 272552
rect 146298 255912 146354 255921
rect 146298 255847 146354 255856
rect 146312 255377 146340 255847
rect 146298 255368 146354 255377
rect 146298 255303 146354 255312
rect 145656 215280 145708 215286
rect 145656 215222 145708 215228
rect 145654 160168 145710 160177
rect 145654 160103 145710 160112
rect 145668 135250 145696 160103
rect 145656 135244 145708 135250
rect 145656 135186 145708 135192
rect 145564 29640 145616 29646
rect 145564 29582 145616 29588
rect 146956 21418 146984 272546
rect 147128 264240 147180 264246
rect 147128 264182 147180 264188
rect 147036 198756 147088 198762
rect 147036 198698 147088 198704
rect 147048 25566 147076 198698
rect 147140 185638 147168 264182
rect 147692 260817 147720 413986
rect 148336 345014 148364 422894
rect 149060 396772 149112 396778
rect 149060 396714 149112 396720
rect 148336 344986 148456 345014
rect 148428 332722 148456 344986
rect 148416 332716 148468 332722
rect 148416 332658 148468 332664
rect 148324 309256 148376 309262
rect 148324 309198 148376 309204
rect 147678 260808 147734 260817
rect 147678 260743 147734 260752
rect 147692 260137 147720 260743
rect 147678 260128 147734 260137
rect 147678 260063 147734 260072
rect 147128 185632 147180 185638
rect 147128 185574 147180 185580
rect 147036 25560 147088 25566
rect 147036 25502 147088 25508
rect 146944 21412 146996 21418
rect 146944 21354 146996 21360
rect 137284 3528 137336 3534
rect 137284 3470 137336 3476
rect 140044 3528 140096 3534
rect 140044 3470 140096 3476
rect 141148 3528 141200 3534
rect 141148 3470 141200 3476
rect 143540 3528 143592 3534
rect 143540 3470 143592 3476
rect 144828 3528 144880 3534
rect 148336 3505 148364 309198
rect 148428 275398 148456 332658
rect 149072 303618 149100 396714
rect 190460 394732 190512 394738
rect 190460 394674 190512 394680
rect 153844 336864 153896 336870
rect 153844 336806 153896 336812
rect 151084 328500 151136 328506
rect 151084 328442 151136 328448
rect 149060 303612 149112 303618
rect 149060 303554 149112 303560
rect 149072 302938 149100 303554
rect 149060 302932 149112 302938
rect 149060 302874 149112 302880
rect 149794 288552 149850 288561
rect 149794 288487 149850 288496
rect 149704 281580 149756 281586
rect 149704 281522 149756 281528
rect 148416 275392 148468 275398
rect 148416 275334 148468 275340
rect 148416 271244 148468 271250
rect 148416 271186 148468 271192
rect 148428 202230 148456 271186
rect 148416 202224 148468 202230
rect 148416 202166 148468 202172
rect 149716 200122 149744 281522
rect 149808 218754 149836 288487
rect 149796 218748 149848 218754
rect 149796 218690 149848 218696
rect 149704 200116 149756 200122
rect 149704 200058 149756 200064
rect 149702 193896 149758 193905
rect 149702 193831 149758 193840
rect 148414 152416 148470 152425
rect 148414 152351 148470 152360
rect 148428 117230 148456 152351
rect 148416 117224 148468 117230
rect 148416 117166 148468 117172
rect 149716 49026 149744 193831
rect 149704 49020 149756 49026
rect 149704 48962 149756 48968
rect 151096 31074 151124 328442
rect 151268 314696 151320 314702
rect 151268 314638 151320 314644
rect 151280 305658 151308 314638
rect 151268 305652 151320 305658
rect 151268 305594 151320 305600
rect 152464 305040 152516 305046
rect 151174 305008 151230 305017
rect 152464 304982 152516 304988
rect 151174 304943 151230 304952
rect 151188 186998 151216 304943
rect 151268 253972 151320 253978
rect 151268 253914 151320 253920
rect 151280 209778 151308 253914
rect 151268 209772 151320 209778
rect 151268 209714 151320 209720
rect 151176 186992 151228 186998
rect 151176 186934 151228 186940
rect 151174 165744 151230 165753
rect 151174 165679 151230 165688
rect 151188 128246 151216 165679
rect 151176 128240 151228 128246
rect 151176 128182 151228 128188
rect 151084 31068 151136 31074
rect 151084 31010 151136 31016
rect 144828 3470 144880 3476
rect 148322 3496 148378 3505
rect 140056 480 140084 3470
rect 143552 480 143580 3470
rect 148322 3431 148378 3440
rect 152476 3369 152504 304982
rect 152648 278112 152700 278118
rect 152648 278054 152700 278060
rect 152556 265736 152608 265742
rect 152556 265678 152608 265684
rect 152568 257446 152596 265678
rect 152556 257440 152608 257446
rect 152556 257382 152608 257388
rect 152556 202836 152608 202842
rect 152556 202778 152608 202784
rect 152568 54534 152596 202778
rect 152660 192506 152688 278054
rect 153856 262886 153884 336806
rect 166356 329860 166408 329866
rect 166356 329802 166408 329808
rect 162124 327140 162176 327146
rect 162124 327082 162176 327088
rect 155222 308136 155278 308145
rect 155222 308071 155278 308080
rect 153934 267064 153990 267073
rect 153934 266999 153990 267008
rect 153844 262880 153896 262886
rect 153844 262822 153896 262828
rect 153844 250504 153896 250510
rect 153844 250446 153896 250452
rect 153200 231124 153252 231130
rect 153200 231066 153252 231072
rect 153212 223553 153240 231066
rect 153198 223544 153254 223553
rect 153198 223479 153254 223488
rect 153856 198762 153884 250446
rect 153948 242214 153976 266999
rect 153936 242208 153988 242214
rect 153936 242150 153988 242156
rect 154028 241596 154080 241602
rect 154028 241538 154080 241544
rect 154040 231742 154068 241538
rect 154028 231736 154080 231742
rect 154028 231678 154080 231684
rect 153844 198756 153896 198762
rect 153844 198698 153896 198704
rect 152648 192500 152700 192506
rect 152648 192442 152700 192448
rect 153842 161800 153898 161809
rect 153842 161735 153898 161744
rect 153856 131209 153884 161735
rect 154210 157448 154266 157457
rect 154210 157383 154266 157392
rect 154224 152522 154252 157383
rect 154212 152516 154264 152522
rect 154212 152458 154264 152464
rect 153936 133204 153988 133210
rect 153936 133146 153988 133152
rect 153842 131200 153898 131209
rect 153842 131135 153898 131144
rect 153948 121446 153976 133146
rect 153936 121440 153988 121446
rect 153936 121382 153988 121388
rect 153844 111920 153896 111926
rect 153844 111862 153896 111868
rect 153856 82822 153884 111862
rect 153844 82816 153896 82822
rect 153844 82758 153896 82764
rect 152556 54528 152608 54534
rect 152556 54470 152608 54476
rect 155236 3466 155264 308071
rect 159362 303920 159418 303929
rect 159362 303855 159418 303864
rect 156604 295384 156656 295390
rect 156604 295326 156656 295332
rect 155406 276720 155462 276729
rect 155406 276655 155462 276664
rect 155314 262848 155370 262857
rect 155314 262783 155370 262792
rect 155328 202842 155356 262783
rect 155420 249121 155448 276655
rect 155406 249112 155462 249121
rect 155406 249047 155462 249056
rect 155408 240780 155460 240786
rect 155408 240722 155460 240728
rect 155420 204270 155448 240722
rect 155408 204264 155460 204270
rect 155408 204206 155460 204212
rect 155316 202836 155368 202842
rect 155316 202778 155368 202784
rect 155316 153264 155368 153270
rect 155316 153206 155368 153212
rect 155328 126274 155356 153206
rect 156616 131102 156644 295326
rect 158074 284880 158130 284889
rect 158074 284815 158130 284824
rect 156696 273964 156748 273970
rect 156696 273906 156748 273912
rect 156708 238513 156736 273906
rect 157984 266416 158036 266422
rect 157984 266358 158036 266364
rect 156694 238504 156750 238513
rect 156694 238439 156750 238448
rect 156708 178158 156736 238439
rect 157246 237960 157302 237969
rect 157246 237895 157302 237904
rect 157260 230489 157288 237895
rect 157246 230480 157302 230489
rect 157246 230415 157302 230424
rect 156696 178152 156748 178158
rect 156696 178094 156748 178100
rect 156604 131096 156656 131102
rect 156604 131038 156656 131044
rect 155316 126268 155368 126274
rect 155316 126210 155368 126216
rect 156708 125526 156736 178094
rect 156696 125520 156748 125526
rect 156696 125462 156748 125468
rect 157260 112470 157288 230415
rect 157248 112464 157300 112470
rect 157248 112406 157300 112412
rect 157260 111926 157288 112406
rect 156604 111920 156656 111926
rect 156604 111862 156656 111868
rect 157248 111920 157300 111926
rect 157248 111862 157300 111868
rect 156616 84153 156644 111862
rect 156602 84144 156658 84153
rect 156602 84079 156658 84088
rect 157996 71058 158024 266358
rect 158088 153882 158116 284815
rect 158720 284436 158772 284442
rect 158720 284378 158772 284384
rect 158732 281518 158760 284378
rect 158720 281512 158772 281518
rect 158720 281454 158772 281460
rect 158076 153876 158128 153882
rect 158076 153818 158128 153824
rect 158088 120086 158116 153818
rect 158076 120080 158128 120086
rect 158076 120022 158128 120028
rect 158732 88330 158760 281454
rect 158720 88324 158772 88330
rect 158720 88266 158772 88272
rect 157984 71052 158036 71058
rect 157984 70994 158036 71000
rect 159376 6186 159404 303855
rect 159456 299532 159508 299538
rect 159456 299474 159508 299480
rect 159468 287706 159496 299474
rect 160098 298752 160154 298761
rect 160098 298687 160154 298696
rect 160112 298110 160140 298687
rect 160100 298104 160152 298110
rect 160100 298046 160152 298052
rect 161296 298104 161348 298110
rect 161296 298046 161348 298052
rect 159456 287700 159508 287706
rect 159456 287642 159508 287648
rect 160742 286376 160798 286385
rect 160742 286311 160798 286320
rect 159456 269816 159508 269822
rect 159456 269758 159508 269764
rect 159468 237153 159496 269758
rect 159548 249824 159600 249830
rect 159548 249766 159600 249772
rect 159454 237144 159510 237153
rect 159454 237079 159510 237088
rect 159560 227662 159588 249766
rect 159914 237144 159970 237153
rect 159914 237079 159970 237088
rect 159548 227656 159600 227662
rect 159548 227598 159600 227604
rect 159928 149734 159956 237079
rect 160100 229016 160152 229022
rect 160100 228958 160152 228964
rect 160008 227656 160060 227662
rect 160008 227598 160060 227604
rect 159916 149728 159968 149734
rect 159916 149670 159968 149676
rect 160020 109041 160048 227598
rect 159454 109032 159510 109041
rect 159454 108967 159510 108976
rect 160006 109032 160062 109041
rect 160006 108967 160062 108976
rect 159468 81394 159496 108967
rect 160112 101454 160140 228958
rect 160756 215966 160784 286311
rect 160836 249076 160888 249082
rect 160836 249018 160888 249024
rect 160848 229022 160876 249018
rect 160926 235376 160982 235385
rect 160926 235311 160982 235320
rect 160836 229016 160888 229022
rect 160836 228958 160888 228964
rect 160940 226302 160968 235311
rect 160928 226296 160980 226302
rect 160928 226238 160980 226244
rect 160744 215960 160796 215966
rect 160744 215902 160796 215908
rect 160836 156052 160888 156058
rect 160836 155994 160888 156000
rect 160848 144906 160876 155994
rect 161308 145042 161336 298046
rect 162136 250510 162164 327082
rect 162860 287088 162912 287094
rect 162860 287030 162912 287036
rect 162872 281518 162900 287030
rect 164976 284368 165028 284374
rect 164976 284310 165028 284316
rect 162860 281512 162912 281518
rect 162860 281454 162912 281460
rect 164148 281512 164200 281518
rect 164148 281454 164200 281460
rect 164160 280838 164188 281454
rect 164148 280832 164200 280838
rect 164148 280774 164200 280780
rect 162214 269784 162270 269793
rect 162214 269719 162270 269728
rect 162124 250504 162176 250510
rect 162124 250446 162176 250452
rect 161480 242956 161532 242962
rect 161480 242898 161532 242904
rect 161388 217320 161440 217326
rect 161388 217262 161440 217268
rect 161400 216646 161428 217262
rect 161388 216640 161440 216646
rect 161388 216582 161440 216588
rect 160928 145036 160980 145042
rect 160928 144978 160980 144984
rect 161296 145036 161348 145042
rect 161296 144978 161348 144984
rect 160836 144900 160888 144906
rect 160836 144842 160888 144848
rect 160742 143576 160798 143585
rect 160742 143511 160798 143520
rect 160756 109002 160784 143511
rect 160940 135930 160968 144978
rect 160928 135924 160980 135930
rect 160928 135866 160980 135872
rect 160836 109064 160888 109070
rect 160836 109006 160888 109012
rect 160744 108996 160796 109002
rect 160744 108938 160796 108944
rect 160100 101448 160152 101454
rect 160100 101390 160152 101396
rect 160848 84153 160876 109006
rect 160834 84144 160890 84153
rect 161492 84114 161520 242898
rect 162122 241632 162178 241641
rect 162122 241567 162178 241576
rect 162136 226137 162164 241567
rect 162228 232665 162256 269719
rect 163504 251252 163556 251258
rect 163504 251194 163556 251200
rect 162214 232656 162270 232665
rect 162214 232591 162270 232600
rect 162122 226128 162178 226137
rect 162122 226063 162178 226072
rect 162136 225049 162164 226063
rect 162122 225040 162178 225049
rect 162122 224975 162178 224984
rect 162766 225040 162822 225049
rect 162766 224975 162822 224984
rect 161572 216640 161624 216646
rect 161572 216582 161624 216588
rect 161584 144945 161612 216582
rect 161570 144936 161626 144945
rect 161570 144871 161626 144880
rect 162122 144936 162178 144945
rect 162122 144871 162178 144880
rect 162136 117201 162164 144871
rect 162122 117192 162178 117201
rect 162122 117127 162178 117136
rect 162780 107642 162808 224975
rect 162768 107636 162820 107642
rect 162768 107578 162820 107584
rect 162124 103556 162176 103562
rect 162124 103498 162176 103504
rect 160834 84079 160890 84088
rect 161480 84108 161532 84114
rect 161480 84050 161532 84056
rect 159456 81388 159508 81394
rect 159456 81330 159508 81336
rect 162136 70378 162164 103498
rect 162768 84108 162820 84114
rect 162768 84050 162820 84056
rect 162780 79966 162808 84050
rect 162768 79960 162820 79966
rect 162768 79902 162820 79908
rect 162124 70372 162176 70378
rect 162124 70314 162176 70320
rect 163516 39370 163544 251194
rect 164160 156466 164188 280774
rect 164884 267776 164936 267782
rect 164884 267718 164936 267724
rect 163596 156460 163648 156466
rect 163596 156402 163648 156408
rect 164148 156460 164200 156466
rect 164148 156402 164200 156408
rect 163608 138718 163636 156402
rect 164160 156058 164188 156402
rect 164148 156052 164200 156058
rect 164148 155994 164200 156000
rect 163596 138712 163648 138718
rect 163596 138654 163648 138660
rect 164896 69698 164924 267718
rect 164988 250510 165016 284310
rect 166264 269136 166316 269142
rect 166264 269078 166316 269084
rect 164976 250504 165028 250510
rect 164976 250446 165028 250452
rect 165528 244316 165580 244322
rect 165528 244258 165580 244264
rect 165540 241398 165568 244258
rect 165528 241392 165580 241398
rect 165528 241334 165580 241340
rect 165540 93158 165568 241334
rect 165528 93152 165580 93158
rect 165528 93094 165580 93100
rect 166170 92440 166226 92449
rect 166170 92375 166226 92384
rect 166184 91798 166212 92375
rect 166172 91792 166224 91798
rect 166172 91734 166224 91740
rect 164884 69692 164936 69698
rect 164884 69634 164936 69640
rect 163504 39364 163556 39370
rect 163504 39306 163556 39312
rect 166276 19990 166304 269078
rect 166368 268394 166396 329802
rect 190472 325694 190500 394674
rect 260840 343664 260892 343670
rect 260840 343606 260892 343612
rect 259828 339516 259880 339522
rect 259828 339458 259880 339464
rect 222200 338156 222252 338162
rect 222200 338098 222252 338104
rect 192484 328568 192536 328574
rect 192484 328510 192536 328516
rect 201498 328536 201554 328545
rect 190472 325666 190592 325694
rect 180064 321700 180116 321706
rect 180064 321642 180116 321648
rect 175924 306400 175976 306406
rect 175924 306342 175976 306348
rect 170404 303748 170456 303754
rect 170404 303690 170456 303696
rect 169024 293276 169076 293282
rect 169024 293218 169076 293224
rect 168288 288448 168340 288454
rect 168288 288390 168340 288396
rect 166908 287700 166960 287706
rect 166908 287642 166960 287648
rect 166920 287094 166948 287642
rect 166908 287088 166960 287094
rect 166908 287030 166960 287036
rect 166356 268388 166408 268394
rect 166356 268330 166408 268336
rect 166356 247784 166408 247790
rect 166356 247726 166408 247732
rect 166368 223582 166396 247726
rect 166356 223576 166408 223582
rect 166356 223518 166408 223524
rect 166356 192500 166408 192506
rect 166356 192442 166408 192448
rect 166368 136610 166396 192442
rect 166356 136604 166408 136610
rect 166356 136546 166408 136552
rect 166368 105670 166396 136546
rect 166356 105664 166408 105670
rect 166356 105606 166408 105612
rect 166920 93906 166948 287030
rect 167644 264988 167696 264994
rect 167644 264930 167696 264936
rect 166908 93900 166960 93906
rect 166908 93842 166960 93848
rect 166920 92410 166948 93842
rect 166908 92404 166960 92410
rect 166908 92346 166960 92352
rect 167656 26926 167684 264930
rect 167736 239420 167788 239426
rect 167736 239362 167788 239368
rect 167748 86970 167776 239362
rect 168300 147762 168328 288390
rect 169036 283626 169064 293218
rect 169024 283620 169076 283626
rect 169024 283562 169076 283568
rect 167828 147756 167880 147762
rect 167828 147698 167880 147704
rect 168288 147756 168340 147762
rect 168288 147698 168340 147704
rect 167840 138689 167868 147698
rect 169036 147014 169064 283562
rect 169208 276684 169260 276690
rect 169208 276626 169260 276632
rect 169116 253972 169168 253978
rect 169116 253914 169168 253920
rect 169128 149705 169156 253914
rect 169220 249082 169248 276626
rect 169298 255912 169354 255921
rect 169298 255847 169354 255856
rect 169208 249076 169260 249082
rect 169208 249018 169260 249024
rect 169208 243568 169260 243574
rect 169208 243510 169260 243516
rect 169220 220726 169248 243510
rect 169312 242282 169340 255847
rect 169300 242276 169352 242282
rect 169300 242218 169352 242224
rect 169208 220720 169260 220726
rect 169208 220662 169260 220668
rect 169668 220720 169720 220726
rect 169668 220662 169720 220668
rect 169114 149696 169170 149705
rect 169114 149631 169170 149640
rect 169298 149152 169354 149161
rect 169298 149087 169354 149096
rect 169024 147008 169076 147014
rect 169024 146950 169076 146956
rect 167826 138680 167882 138689
rect 167826 138615 167882 138624
rect 169312 117298 169340 149087
rect 169300 117292 169352 117298
rect 169300 117234 169352 117240
rect 169024 100768 169076 100774
rect 169024 100710 169076 100716
rect 167736 86964 167788 86970
rect 167736 86906 167788 86912
rect 169036 73166 169064 100710
rect 169680 95946 169708 220662
rect 169760 129056 169812 129062
rect 169760 128998 169812 129004
rect 169772 128382 169800 128998
rect 169760 128376 169812 128382
rect 169760 128318 169812 128324
rect 169668 95940 169720 95946
rect 169668 95882 169720 95888
rect 169024 73160 169076 73166
rect 169024 73102 169076 73108
rect 170416 72486 170444 303690
rect 173254 293176 173310 293185
rect 173254 293111 173310 293120
rect 172426 287736 172482 287745
rect 172426 287671 172482 287680
rect 170586 273864 170642 273873
rect 170586 273799 170642 273808
rect 170496 249824 170548 249830
rect 170496 249766 170548 249772
rect 170404 72480 170456 72486
rect 170404 72422 170456 72428
rect 167644 26920 167696 26926
rect 167644 26862 167696 26868
rect 170508 24138 170536 249766
rect 170600 235958 170628 273799
rect 171784 260908 171836 260914
rect 171784 260850 171836 260856
rect 170588 235952 170640 235958
rect 170588 235894 170640 235900
rect 170586 233336 170642 233345
rect 170586 233271 170642 233280
rect 170600 209774 170628 233271
rect 170600 209746 170996 209774
rect 170968 200054 170996 209746
rect 170956 200048 171008 200054
rect 170956 199990 171008 199996
rect 170968 120834 170996 199990
rect 171048 128376 171100 128382
rect 171048 128318 171100 128324
rect 170956 120828 171008 120834
rect 170956 120770 171008 120776
rect 171060 44878 171088 128318
rect 171796 75206 171824 260850
rect 171874 226400 171930 226409
rect 171874 226335 171930 226344
rect 171888 201482 171916 226335
rect 171876 201476 171928 201482
rect 171876 201418 171928 201424
rect 172336 201476 172388 201482
rect 172336 201418 172388 201424
rect 172348 114617 172376 201418
rect 172334 114608 172390 114617
rect 172334 114543 172390 114552
rect 172440 90982 172468 287671
rect 173268 267034 173296 293111
rect 175936 272542 175964 306342
rect 177302 305144 177358 305153
rect 177302 305079 177358 305088
rect 176108 286408 176160 286414
rect 176108 286350 176160 286356
rect 175924 272536 175976 272542
rect 175924 272478 175976 272484
rect 176014 268424 176070 268433
rect 176014 268359 176070 268368
rect 173256 267028 173308 267034
rect 173256 266970 173308 266976
rect 173164 266484 173216 266490
rect 173164 266426 173216 266432
rect 172428 90976 172480 90982
rect 172428 90918 172480 90924
rect 171784 75200 171836 75206
rect 171784 75142 171836 75148
rect 173176 73846 173204 266426
rect 173346 260128 173402 260137
rect 173346 260063 173402 260072
rect 173256 257372 173308 257378
rect 173256 257314 173308 257320
rect 173268 226302 173296 257314
rect 173360 247625 173388 260063
rect 174544 259480 174596 259486
rect 174544 259422 174596 259428
rect 173346 247616 173402 247625
rect 173346 247551 173402 247560
rect 173256 226296 173308 226302
rect 173256 226238 173308 226244
rect 173268 225010 173296 226238
rect 173256 225004 173308 225010
rect 173256 224946 173308 224952
rect 173808 225004 173860 225010
rect 173808 224946 173860 224952
rect 173254 158808 173310 158817
rect 173254 158743 173310 158752
rect 173268 125594 173296 158743
rect 173348 144152 173400 144158
rect 173348 144094 173400 144100
rect 173256 125588 173308 125594
rect 173256 125530 173308 125536
rect 173360 115870 173388 144094
rect 173820 141545 173848 224946
rect 173806 141536 173862 141545
rect 173806 141471 173862 141480
rect 173820 141438 173848 141471
rect 173808 141432 173860 141438
rect 173808 141374 173860 141380
rect 173348 115864 173400 115870
rect 173348 115806 173400 115812
rect 173256 108316 173308 108322
rect 173256 108258 173308 108264
rect 173268 85474 173296 108258
rect 173348 99408 173400 99414
rect 173348 99350 173400 99356
rect 173256 85468 173308 85474
rect 173256 85410 173308 85416
rect 173360 81394 173388 99350
rect 173348 81388 173400 81394
rect 173348 81330 173400 81336
rect 174556 76537 174584 259422
rect 175924 258120 175976 258126
rect 175924 258062 175976 258068
rect 174634 251288 174690 251297
rect 174634 251223 174690 251232
rect 174648 224942 174676 251223
rect 174636 224936 174688 224942
rect 174636 224878 174688 224884
rect 174728 224256 174780 224262
rect 174728 224198 174780 224204
rect 174740 214606 174768 224198
rect 175186 217424 175242 217433
rect 175186 217359 175242 217368
rect 175200 216753 175228 217359
rect 175186 216744 175242 216753
rect 175186 216679 175242 216688
rect 174728 214600 174780 214606
rect 174728 214542 174780 214548
rect 175200 100706 175228 216679
rect 175832 153332 175884 153338
rect 175832 153274 175884 153280
rect 175844 147121 175872 153274
rect 175830 147112 175886 147121
rect 175830 147047 175886 147056
rect 175188 100700 175240 100706
rect 175188 100642 175240 100648
rect 174542 76528 174598 76537
rect 174542 76463 174598 76472
rect 173164 73840 173216 73846
rect 173164 73782 173216 73788
rect 175936 47598 175964 258062
rect 176028 234598 176056 268359
rect 176120 264246 176148 286350
rect 177316 280809 177344 305079
rect 178684 300892 178736 300898
rect 178684 300834 178736 300840
rect 178038 282976 178094 282985
rect 178038 282911 178040 282920
rect 178092 282911 178094 282920
rect 178040 282882 178092 282888
rect 177302 280800 177358 280809
rect 177302 280735 177358 280744
rect 177856 278044 177908 278050
rect 177856 277986 177908 277992
rect 177868 277394 177896 277986
rect 177868 277370 177988 277394
rect 177868 277366 178000 277370
rect 176108 264240 176160 264246
rect 176108 264182 176160 264188
rect 177304 262336 177356 262342
rect 177304 262278 177356 262284
rect 176566 240816 176622 240825
rect 176566 240751 176622 240760
rect 176016 234592 176068 234598
rect 176016 234534 176068 234540
rect 176580 92449 176608 240751
rect 176566 92440 176622 92449
rect 176566 92375 176622 92384
rect 175924 47592 175976 47598
rect 175924 47534 175976 47540
rect 171048 44872 171100 44878
rect 171048 44814 171100 44820
rect 170496 24132 170548 24138
rect 170496 24074 170548 24080
rect 166264 19984 166316 19990
rect 166264 19926 166316 19932
rect 177316 18630 177344 262278
rect 177396 247716 177448 247722
rect 177396 247658 177448 247664
rect 177408 233238 177436 247658
rect 177396 233232 177448 233238
rect 177396 233174 177448 233180
rect 177868 171222 177896 277366
rect 177948 277364 178000 277366
rect 177948 277306 178000 277312
rect 178696 260166 178724 300834
rect 179328 300212 179380 300218
rect 179328 300154 179380 300160
rect 179236 282940 179288 282946
rect 179236 282882 179288 282888
rect 178684 260160 178736 260166
rect 178684 260102 178736 260108
rect 178684 257440 178736 257446
rect 178684 257382 178736 257388
rect 178696 238649 178724 257382
rect 178682 238640 178738 238649
rect 178682 238575 178738 238584
rect 177948 233232 178000 233238
rect 177948 233174 178000 233180
rect 177856 171216 177908 171222
rect 177856 171158 177908 171164
rect 177868 170474 177896 171158
rect 177856 170468 177908 170474
rect 177856 170410 177908 170416
rect 177396 155236 177448 155242
rect 177396 155178 177448 155184
rect 177408 129742 177436 155178
rect 177396 129736 177448 129742
rect 177396 129678 177448 129684
rect 177396 111852 177448 111858
rect 177396 111794 177448 111800
rect 177408 75818 177436 111794
rect 177960 78606 177988 233174
rect 178684 214600 178736 214606
rect 178684 214542 178736 214548
rect 178696 191826 178724 214542
rect 178684 191820 178736 191826
rect 178684 191762 178736 191768
rect 178696 147801 178724 191762
rect 178776 154624 178828 154630
rect 178776 154566 178828 154572
rect 178682 147792 178738 147801
rect 178682 147727 178738 147736
rect 178696 124098 178724 147727
rect 178788 145625 178816 154566
rect 178774 145616 178830 145625
rect 178774 145551 178830 145560
rect 178684 124092 178736 124098
rect 178684 124034 178736 124040
rect 178776 98660 178828 98666
rect 178776 98602 178828 98608
rect 178684 93152 178736 93158
rect 178684 93094 178736 93100
rect 177948 78600 178000 78606
rect 177948 78542 178000 78548
rect 177396 75812 177448 75818
rect 177396 75754 177448 75760
rect 178696 73098 178724 93094
rect 178788 88262 178816 98602
rect 179248 92546 179276 282882
rect 179236 92540 179288 92546
rect 179236 92482 179288 92488
rect 179340 91050 179368 300154
rect 180076 288386 180104 321642
rect 185584 316124 185636 316130
rect 185584 316066 185636 316072
rect 182916 306468 182968 306474
rect 182916 306410 182968 306416
rect 180154 305280 180210 305289
rect 180154 305215 180210 305224
rect 180064 288380 180116 288386
rect 180064 288322 180116 288328
rect 180064 273284 180116 273290
rect 180064 273226 180116 273232
rect 179420 235952 179472 235958
rect 179420 235894 179472 235900
rect 179432 235521 179460 235894
rect 179418 235512 179474 235521
rect 179418 235447 179474 235456
rect 180076 145586 180104 273226
rect 180168 272610 180196 305215
rect 182822 303784 182878 303793
rect 182822 303719 182878 303728
rect 180248 294636 180300 294642
rect 180248 294578 180300 294584
rect 180156 272604 180208 272610
rect 180156 272546 180208 272552
rect 180260 262857 180288 294578
rect 181628 275324 181680 275330
rect 181628 275266 181680 275272
rect 181536 271924 181588 271930
rect 181536 271866 181588 271872
rect 180246 262848 180302 262857
rect 180246 262783 180302 262792
rect 180248 261520 180300 261526
rect 180248 261462 180300 261468
rect 180154 235648 180210 235657
rect 180154 235583 180210 235592
rect 180168 202842 180196 235583
rect 180260 231810 180288 261462
rect 180338 257272 180394 257281
rect 180338 257207 180394 257216
rect 180352 234025 180380 257207
rect 181444 255332 181496 255338
rect 181444 255274 181496 255280
rect 180338 234016 180394 234025
rect 180338 233951 180394 233960
rect 180248 231804 180300 231810
rect 180248 231746 180300 231752
rect 180156 202836 180208 202842
rect 180156 202778 180208 202784
rect 180708 202836 180760 202842
rect 180708 202778 180760 202784
rect 180154 178664 180210 178673
rect 180154 178599 180210 178608
rect 180064 145580 180116 145586
rect 180064 145522 180116 145528
rect 180064 135312 180116 135318
rect 180064 135254 180116 135260
rect 179328 91044 179380 91050
rect 179328 90986 179380 90992
rect 178776 88256 178828 88262
rect 178776 88198 178828 88204
rect 178684 73092 178736 73098
rect 178684 73034 178736 73040
rect 177304 18624 177356 18630
rect 177304 18566 177356 18572
rect 180076 7682 180104 135254
rect 180168 126954 180196 178599
rect 180248 151904 180300 151910
rect 180248 151846 180300 151852
rect 180260 144158 180288 151846
rect 180248 144152 180300 144158
rect 180248 144094 180300 144100
rect 180156 126948 180208 126954
rect 180156 126890 180208 126896
rect 180168 118017 180196 126890
rect 180154 118008 180210 118017
rect 180154 117943 180210 117952
rect 180156 105596 180208 105602
rect 180156 105538 180208 105544
rect 180168 74458 180196 105538
rect 180248 104168 180300 104174
rect 180248 104110 180300 104116
rect 180260 75886 180288 104110
rect 180720 81433 180748 202778
rect 180800 161492 180852 161498
rect 180800 161434 180852 161440
rect 180812 159390 180840 161434
rect 180800 159384 180852 159390
rect 180800 159326 180852 159332
rect 180706 81424 180762 81433
rect 180706 81359 180762 81368
rect 180248 75880 180300 75886
rect 180248 75822 180300 75828
rect 180156 74452 180208 74458
rect 180156 74394 180208 74400
rect 180260 50386 180288 75822
rect 181456 58682 181484 255274
rect 181548 236706 181576 271866
rect 181640 241466 181668 275266
rect 181628 241460 181680 241466
rect 181628 241402 181680 241408
rect 181640 238754 181668 241402
rect 181640 238726 182036 238754
rect 181536 236700 181588 236706
rect 181536 236642 181588 236648
rect 181534 214024 181590 214033
rect 181534 213959 181590 213968
rect 181548 209681 181576 213959
rect 181534 209672 181590 209681
rect 181534 209607 181590 209616
rect 182008 161498 182036 238726
rect 182086 209672 182142 209681
rect 182086 209607 182142 209616
rect 181996 161492 182048 161498
rect 181996 161434 182048 161440
rect 181536 133952 181588 133958
rect 181536 133894 181588 133900
rect 181548 128314 181576 133894
rect 181536 128308 181588 128314
rect 181536 128250 181588 128256
rect 181444 58676 181496 58682
rect 181444 58618 181496 58624
rect 180248 50380 180300 50386
rect 180248 50322 180300 50328
rect 181548 43450 181576 128250
rect 182100 109177 182128 209607
rect 182178 144800 182234 144809
rect 182178 144735 182234 144744
rect 182192 135969 182220 144735
rect 182178 135960 182234 135969
rect 182178 135895 182234 135904
rect 182086 109168 182142 109177
rect 182086 109103 182142 109112
rect 182836 82113 182864 303719
rect 182928 265674 182956 306410
rect 184204 296744 184256 296750
rect 184204 296686 184256 296692
rect 182916 265668 182968 265674
rect 182916 265610 182968 265616
rect 182914 261488 182970 261497
rect 182914 261423 182970 261432
rect 182928 219337 182956 261423
rect 184216 233889 184244 296686
rect 185596 280158 185624 316066
rect 186320 313404 186372 313410
rect 186320 313346 186372 313352
rect 186332 309126 186360 313346
rect 187148 311908 187200 311914
rect 187148 311850 187200 311856
rect 187054 309496 187110 309505
rect 187054 309431 187110 309440
rect 186320 309120 186372 309126
rect 186320 309062 186372 309068
rect 186962 296712 187018 296721
rect 186962 296647 187018 296656
rect 186228 288516 186280 288522
rect 186228 288458 186280 288464
rect 185584 280152 185636 280158
rect 185584 280094 185636 280100
rect 185766 258768 185822 258777
rect 185766 258703 185822 258712
rect 185584 256760 185636 256766
rect 185584 256702 185636 256708
rect 184388 254584 184440 254590
rect 184388 254526 184440 254532
rect 184296 247104 184348 247110
rect 184296 247046 184348 247052
rect 184202 233880 184258 233889
rect 184202 233815 184258 233824
rect 182914 219328 182970 219337
rect 182914 219263 182970 219272
rect 182928 218113 182956 219263
rect 182914 218104 182970 218113
rect 182914 218039 182970 218048
rect 183466 218104 183522 218113
rect 183466 218039 183522 218048
rect 182916 169040 182968 169046
rect 182916 168982 182968 168988
rect 182928 133890 182956 168982
rect 183480 144809 183508 218039
rect 184308 209098 184336 247046
rect 184400 237386 184428 254526
rect 184388 237380 184440 237386
rect 184388 237322 184440 237328
rect 184296 209092 184348 209098
rect 184296 209034 184348 209040
rect 184478 161664 184534 161673
rect 184478 161599 184534 161608
rect 184202 149696 184258 149705
rect 184202 149631 184258 149640
rect 183466 144800 183522 144809
rect 183466 144735 183522 144744
rect 183480 143585 183508 144735
rect 183466 143576 183522 143585
rect 183466 143511 183522 143520
rect 182916 133884 182968 133890
rect 182916 133826 182968 133832
rect 182928 122126 182956 133826
rect 184216 124166 184244 149631
rect 184294 147248 184350 147257
rect 184294 147183 184350 147192
rect 184308 144906 184336 147183
rect 184388 147008 184440 147014
rect 184388 146950 184440 146956
rect 184296 144900 184348 144906
rect 184296 144842 184348 144848
rect 184308 124273 184336 144842
rect 184400 136610 184428 146950
rect 184492 145761 184520 161599
rect 185492 149728 185544 149734
rect 185492 149670 185544 149676
rect 184478 145752 184534 145761
rect 184478 145687 184534 145696
rect 185504 144226 185532 149670
rect 185492 144220 185544 144226
rect 185492 144162 185544 144168
rect 184848 139596 184900 139602
rect 184848 139538 184900 139544
rect 184860 137970 184888 139538
rect 184848 137964 184900 137970
rect 184848 137906 184900 137912
rect 184388 136604 184440 136610
rect 184388 136546 184440 136552
rect 184294 124264 184350 124273
rect 184294 124199 184350 124208
rect 184204 124160 184256 124166
rect 184204 124102 184256 124108
rect 182916 122120 182968 122126
rect 182916 122062 182968 122068
rect 183468 122120 183520 122126
rect 183468 122062 183520 122068
rect 183376 120760 183428 120766
rect 183376 120702 183428 120708
rect 183388 120154 183416 120702
rect 183376 120148 183428 120154
rect 183376 120090 183428 120096
rect 182822 82104 182878 82113
rect 182822 82039 182878 82048
rect 183388 71058 183416 120090
rect 183376 71052 183428 71058
rect 183376 70994 183428 71000
rect 181536 43444 181588 43450
rect 181536 43386 181588 43392
rect 183480 29646 183508 122062
rect 184848 120828 184900 120834
rect 184848 120770 184900 120776
rect 184296 119400 184348 119406
rect 184296 119342 184348 119348
rect 184204 106344 184256 106350
rect 184204 106286 184256 106292
rect 184216 82657 184244 106286
rect 184308 105942 184336 119342
rect 184860 117298 184888 120770
rect 184848 117292 184900 117298
rect 184848 117234 184900 117240
rect 184756 110900 184808 110906
rect 184756 110842 184808 110848
rect 184296 105936 184348 105942
rect 184296 105878 184348 105884
rect 184296 96688 184348 96694
rect 184296 96630 184348 96636
rect 184308 85377 184336 96630
rect 184294 85368 184350 85377
rect 184294 85303 184350 85312
rect 184202 82648 184258 82657
rect 184202 82583 184258 82592
rect 184768 74497 184796 110842
rect 184848 93900 184900 93906
rect 184848 93842 184900 93848
rect 184754 74488 184810 74497
rect 184754 74423 184810 74432
rect 184860 53106 184888 93842
rect 185596 77897 185624 256702
rect 185676 251320 185728 251326
rect 185676 251262 185728 251268
rect 185688 207670 185716 251262
rect 185780 229094 185808 258703
rect 186240 235278 186268 288458
rect 186976 256018 187004 296647
rect 187068 271182 187096 309431
rect 187160 277370 187188 311850
rect 189816 310548 189868 310554
rect 189816 310490 189868 310496
rect 189722 309360 189778 309369
rect 189722 309295 189778 309304
rect 188436 307896 188488 307902
rect 188436 307838 188488 307844
rect 188342 306640 188398 306649
rect 188342 306575 188398 306584
rect 187148 277364 187200 277370
rect 187148 277306 187200 277312
rect 187148 271992 187200 271998
rect 187148 271934 187200 271940
rect 187056 271176 187108 271182
rect 187056 271118 187108 271124
rect 186964 256012 187016 256018
rect 186964 255954 187016 255960
rect 186964 252612 187016 252618
rect 186964 252554 187016 252560
rect 186228 235272 186280 235278
rect 186228 235214 186280 235220
rect 185780 229066 186268 229094
rect 186240 227633 186268 229066
rect 186226 227624 186282 227633
rect 186226 227559 186282 227568
rect 186134 223000 186190 223009
rect 186134 222935 186190 222944
rect 186148 222329 186176 222935
rect 186134 222320 186190 222329
rect 186134 222255 186190 222264
rect 185676 207664 185728 207670
rect 185676 207606 185728 207612
rect 186148 108225 186176 222255
rect 186134 108216 186190 108225
rect 186134 108151 186190 108160
rect 186136 95940 186188 95946
rect 186136 95882 186188 95888
rect 185676 92608 185728 92614
rect 185676 92550 185728 92556
rect 185688 82754 185716 92550
rect 185676 82748 185728 82754
rect 185676 82690 185728 82696
rect 185582 77888 185638 77897
rect 185582 77823 185638 77832
rect 184848 53100 184900 53106
rect 184848 53042 184900 53048
rect 186148 51746 186176 95882
rect 186240 89593 186268 227559
rect 186320 218068 186372 218074
rect 186320 218010 186372 218016
rect 186332 211070 186360 218010
rect 186320 211064 186372 211070
rect 186320 211006 186372 211012
rect 186976 148345 187004 252554
rect 187054 249112 187110 249121
rect 187054 249047 187110 249056
rect 187068 221610 187096 249047
rect 187160 238066 187188 271934
rect 188356 271250 188384 306575
rect 188448 291145 188476 307838
rect 188710 301336 188766 301345
rect 188710 301271 188766 301280
rect 188526 301200 188582 301209
rect 188526 301135 188582 301144
rect 188434 291136 188490 291145
rect 188434 291071 188490 291080
rect 188436 286340 188488 286346
rect 188436 286282 188488 286288
rect 188344 271244 188396 271250
rect 188344 271186 188396 271192
rect 187240 245676 187292 245682
rect 187240 245618 187292 245624
rect 187148 238060 187200 238066
rect 187148 238002 187200 238008
rect 187252 232529 187280 245618
rect 188342 241632 188398 241641
rect 188342 241567 188398 241576
rect 187238 232520 187294 232529
rect 187238 232455 187294 232464
rect 187056 221604 187108 221610
rect 187056 221546 187108 221552
rect 187608 189780 187660 189786
rect 187608 189722 187660 189728
rect 187054 156088 187110 156097
rect 187054 156023 187110 156032
rect 186962 148336 187018 148345
rect 186962 148271 187018 148280
rect 186964 143676 187016 143682
rect 186964 143618 187016 143624
rect 186976 132462 187004 143618
rect 186964 132456 187016 132462
rect 186964 132398 187016 132404
rect 186964 118720 187016 118726
rect 186964 118662 187016 118668
rect 186226 89584 186282 89593
rect 186226 89519 186282 89528
rect 186136 51740 186188 51746
rect 186136 51682 186188 51688
rect 186976 40730 187004 118662
rect 187068 115938 187096 156023
rect 187146 150512 187202 150521
rect 187146 150447 187202 150456
rect 187160 133210 187188 150447
rect 187148 133204 187200 133210
rect 187148 133146 187200 133152
rect 187516 122868 187568 122874
rect 187516 122810 187568 122816
rect 187528 120086 187556 122810
rect 187516 120080 187568 120086
rect 187516 120022 187568 120028
rect 187528 118726 187556 120022
rect 187516 118720 187568 118726
rect 187516 118662 187568 118668
rect 187056 115932 187108 115938
rect 187056 115874 187108 115880
rect 187148 113212 187200 113218
rect 187148 113154 187200 113160
rect 187056 109064 187108 109070
rect 187056 109006 187108 109012
rect 187068 74526 187096 109006
rect 187160 78577 187188 113154
rect 187620 107846 187648 189722
rect 188356 182850 188384 241567
rect 188448 238746 188476 286282
rect 188540 278118 188568 301135
rect 188724 286414 188752 301271
rect 189736 289785 189764 309295
rect 189828 301510 189856 310490
rect 189906 302424 189962 302433
rect 189906 302359 189962 302368
rect 189816 301504 189868 301510
rect 189816 301446 189868 301452
rect 189920 294545 189948 302359
rect 190458 300928 190514 300937
rect 190458 300863 190514 300872
rect 190368 300824 190420 300830
rect 190368 300766 190420 300772
rect 190380 297401 190408 300766
rect 190472 300218 190500 300863
rect 190460 300212 190512 300218
rect 190460 300154 190512 300160
rect 190564 300150 190592 325666
rect 191102 310856 191158 310865
rect 191102 310791 191158 310800
rect 191116 302234 191144 310791
rect 191024 302206 191144 302234
rect 191380 302252 191432 302258
rect 190552 300144 190604 300150
rect 190552 300086 190604 300092
rect 190564 299849 190592 300086
rect 190550 299840 190606 299849
rect 190550 299775 190606 299784
rect 191024 299470 191052 302206
rect 191380 302194 191432 302200
rect 191102 300656 191158 300665
rect 191102 300591 191158 300600
rect 191012 299464 191064 299470
rect 191012 299406 191064 299412
rect 191116 298110 191144 300591
rect 191286 298616 191342 298625
rect 191286 298551 191342 298560
rect 191104 298104 191156 298110
rect 191104 298046 191156 298052
rect 191194 297528 191250 297537
rect 191194 297463 191250 297472
rect 190366 297392 190422 297401
rect 190366 297327 190422 297336
rect 190458 296304 190514 296313
rect 190458 296239 190514 296248
rect 190472 295390 190500 296239
rect 190460 295384 190512 295390
rect 190460 295326 190512 295332
rect 190552 295316 190604 295322
rect 190552 295258 190604 295264
rect 189906 294536 189962 294545
rect 189906 294471 189962 294480
rect 190564 294001 190592 295258
rect 190550 293992 190606 294001
rect 190550 293927 190606 293936
rect 191102 291680 191158 291689
rect 191102 291615 191158 291624
rect 189722 289776 189778 289785
rect 189722 289711 189778 289720
rect 191010 289368 191066 289377
rect 191010 289303 191066 289312
rect 191024 288522 191052 289303
rect 191012 288516 191064 288522
rect 191012 288458 191064 288464
rect 188712 286408 188764 286414
rect 188712 286350 188764 286356
rect 191010 283656 191066 283665
rect 191010 283591 191066 283600
rect 191024 282946 191052 283591
rect 191012 282940 191064 282946
rect 191012 282882 191064 282888
rect 190458 280120 190514 280129
rect 190458 280055 190514 280064
rect 190366 279032 190422 279041
rect 190366 278967 190422 278976
rect 188528 278112 188580 278118
rect 188528 278054 188580 278060
rect 188620 277432 188672 277438
rect 188620 277374 188672 277380
rect 188528 248464 188580 248470
rect 188528 248406 188580 248412
rect 188436 238740 188488 238746
rect 188436 238682 188488 238688
rect 188540 202162 188568 248406
rect 188632 238134 188660 277374
rect 189722 270600 189778 270609
rect 189722 270535 189778 270544
rect 188620 238128 188672 238134
rect 188620 238070 188672 238076
rect 188528 202156 188580 202162
rect 188528 202098 188580 202104
rect 188344 182844 188396 182850
rect 188344 182786 188396 182792
rect 188344 171216 188396 171222
rect 188344 171158 188396 171164
rect 188356 159458 188384 171158
rect 188986 160712 189042 160721
rect 188986 160647 189042 160656
rect 188344 159452 188396 159458
rect 188344 159394 188396 159400
rect 188434 159352 188490 159361
rect 188434 159287 188490 159296
rect 188066 153776 188122 153785
rect 188066 153711 188122 153720
rect 188080 145897 188108 153711
rect 188342 150784 188398 150793
rect 188342 150719 188398 150728
rect 188066 145888 188122 145897
rect 188066 145823 188122 145832
rect 187698 139496 187754 139505
rect 187698 139431 187754 139440
rect 187712 135153 187740 139431
rect 187698 135144 187754 135153
rect 187698 135079 187754 135088
rect 188356 120086 188384 150719
rect 188448 144265 188476 159287
rect 188894 145616 188950 145625
rect 188894 145551 188950 145560
rect 188434 144256 188490 144265
rect 188434 144191 188490 144200
rect 188436 135244 188488 135250
rect 188436 135186 188488 135192
rect 188448 131102 188476 135186
rect 188436 131096 188488 131102
rect 188436 131038 188488 131044
rect 188908 126954 188936 145551
rect 189000 139505 189028 160647
rect 189736 156641 189764 270535
rect 189814 244624 189870 244633
rect 189814 244559 189870 244568
rect 189828 221513 189856 244559
rect 189906 242992 189962 243001
rect 189906 242927 189962 242936
rect 189920 235249 189948 242927
rect 189906 235240 189962 235249
rect 189906 235175 189962 235184
rect 190380 232529 190408 278967
rect 190472 276690 190500 280055
rect 190460 276684 190512 276690
rect 190460 276626 190512 276632
rect 191012 266484 191064 266490
rect 191012 266426 191064 266432
rect 191024 266393 191052 266426
rect 191010 266384 191066 266393
rect 191010 266319 191066 266328
rect 190460 258120 190512 258126
rect 190512 258068 190592 258074
rect 190460 258062 190592 258068
rect 190472 258058 190592 258062
rect 190472 258052 190604 258058
rect 190472 258046 190552 258052
rect 190552 257994 190604 258000
rect 190642 255912 190698 255921
rect 190642 255847 190698 255856
rect 190656 255338 190684 255847
rect 190644 255332 190696 255338
rect 190644 255274 190696 255280
rect 190828 251320 190880 251326
rect 190826 251288 190828 251297
rect 190880 251288 190882 251297
rect 190826 251223 190882 251232
rect 190642 246664 190698 246673
rect 190642 246599 190698 246608
rect 190656 245682 190684 246599
rect 190644 245676 190696 245682
rect 190644 245618 190696 245624
rect 190366 232520 190422 232529
rect 190366 232455 190422 232464
rect 189814 221504 189870 221513
rect 189814 221439 189870 221448
rect 189816 160132 189868 160138
rect 189816 160074 189868 160080
rect 189722 156632 189778 156641
rect 189722 156567 189778 156576
rect 189722 151872 189778 151881
rect 189722 151807 189778 151816
rect 189078 142352 189134 142361
rect 189078 142287 189134 142296
rect 189092 140758 189120 142287
rect 189080 140752 189132 140758
rect 189080 140694 189132 140700
rect 188986 139496 189042 139505
rect 188986 139431 189042 139440
rect 189736 138553 189764 151807
rect 189722 138544 189778 138553
rect 189722 138479 189778 138488
rect 189828 133929 189856 160074
rect 190368 158024 190420 158030
rect 190368 157966 190420 157972
rect 189908 157480 189960 157486
rect 189908 157422 189960 157428
rect 189920 148617 189948 157422
rect 189906 148608 189962 148617
rect 189906 148543 189962 148552
rect 189814 133920 189870 133929
rect 189814 133855 189870 133864
rect 190380 133793 190408 157966
rect 190366 133784 190422 133793
rect 190366 133719 190422 133728
rect 190380 132569 190408 133719
rect 190366 132560 190422 132569
rect 190366 132495 190422 132504
rect 191116 132494 191144 291615
rect 191208 284889 191236 297463
rect 191300 287745 191328 298551
rect 191392 293185 191420 302194
rect 192496 296585 192524 328510
rect 201498 328471 201554 328480
rect 212540 328500 212592 328506
rect 196990 306776 197046 306785
rect 196990 306711 197046 306720
rect 192576 305108 192628 305114
rect 192576 305050 192628 305056
rect 192482 296576 192538 296585
rect 192482 296511 192538 296520
rect 192496 296002 192524 296511
rect 192484 295996 192536 296002
rect 192484 295938 192536 295944
rect 192588 293282 192616 305050
rect 195978 302832 196034 302841
rect 195978 302767 196034 302776
rect 195992 301594 196020 302767
rect 195992 301566 196374 301594
rect 197004 301580 197032 306711
rect 200210 302424 200266 302433
rect 200210 302359 200266 302368
rect 198278 302288 198334 302297
rect 198278 302223 198334 302232
rect 198292 301580 198320 302223
rect 200224 301580 200252 302359
rect 201512 301580 201540 328471
rect 212540 328442 212592 328448
rect 203614 311944 203670 311953
rect 203614 311879 203670 311888
rect 201774 309224 201830 309233
rect 201774 309159 201830 309168
rect 201788 301594 201816 309159
rect 202510 308272 202566 308281
rect 202510 308207 202566 308216
rect 202524 307834 202552 308207
rect 202420 307828 202472 307834
rect 202420 307770 202472 307776
rect 202512 307828 202564 307834
rect 202512 307770 202564 307776
rect 202432 301594 202460 307770
rect 203430 305008 203486 305017
rect 203430 304943 203486 304952
rect 201788 301566 202170 301594
rect 202432 301566 202814 301594
rect 203444 301580 203472 304943
rect 203628 301594 203656 311879
rect 204902 310720 204958 310729
rect 204902 310655 204958 310664
rect 204258 310584 204314 310593
rect 204258 310519 204314 310528
rect 204272 301594 204300 310519
rect 204916 301594 204944 310655
rect 208398 309496 208454 309505
rect 208398 309431 208454 309440
rect 207846 301880 207902 301889
rect 207846 301815 207902 301824
rect 203628 301566 204010 301594
rect 204272 301566 204654 301594
rect 204916 301566 205298 301594
rect 207860 301580 207888 301815
rect 208412 301594 208440 309431
rect 209778 306640 209834 306649
rect 209778 306575 209834 306584
rect 208412 301566 208518 301594
rect 209792 301580 209820 306575
rect 210424 306468 210476 306474
rect 210424 306410 210476 306416
rect 210436 301580 210464 306410
rect 212552 306374 212580 328442
rect 212632 327140 212684 327146
rect 212632 327082 212684 327088
rect 212644 325694 212672 327082
rect 222212 325694 222240 338098
rect 233884 336864 233936 336870
rect 233884 336806 233936 336812
rect 227812 329860 227864 329866
rect 227812 329802 227864 329808
rect 227824 325694 227852 329802
rect 212644 325666 213224 325694
rect 222212 325666 222792 325694
rect 227824 325666 227944 325694
rect 212552 306346 212672 306374
rect 211068 302252 211120 302258
rect 211068 302194 211120 302200
rect 211080 301580 211108 302194
rect 212644 301594 212672 306346
rect 213196 301594 213224 325666
rect 220910 313440 220966 313449
rect 220910 313375 220966 313384
rect 220176 309188 220228 309194
rect 220176 309130 220228 309136
rect 219990 308136 220046 308145
rect 219990 308071 220046 308080
rect 218058 308000 218114 308009
rect 218058 307935 218114 307944
rect 214838 305280 214894 305289
rect 214838 305215 214894 305224
rect 214196 303748 214248 303754
rect 214196 303690 214248 303696
rect 213920 303680 213972 303686
rect 213918 303648 213920 303657
rect 213972 303648 213974 303657
rect 213918 303583 213974 303592
rect 212644 301566 213026 301594
rect 213196 301566 213670 301594
rect 214208 301580 214236 303690
rect 214852 301580 214880 305215
rect 215482 305144 215538 305153
rect 215482 305079 215538 305088
rect 215298 303920 215354 303929
rect 215298 303855 215354 303864
rect 215312 303754 215340 303855
rect 215300 303748 215352 303754
rect 215300 303690 215352 303696
rect 215496 301580 215524 305079
rect 216772 305040 216824 305046
rect 216772 304982 216824 304988
rect 216128 303816 216180 303822
rect 216128 303758 216180 303764
rect 216140 301580 216168 303758
rect 216784 301580 216812 304982
rect 218072 301580 218100 307935
rect 220004 301580 220032 308071
rect 220188 301594 220216 309130
rect 220924 301594 220952 313375
rect 222764 301594 222792 325666
rect 224038 314800 224094 314809
rect 224038 314735 224094 314744
rect 224052 301594 224080 314735
rect 226982 303648 227038 303657
rect 226982 303583 227038 303592
rect 220188 301566 220662 301594
rect 220924 301566 221306 301594
rect 222764 301566 223238 301594
rect 224052 301566 224434 301594
rect 226996 301580 227024 303583
rect 227916 301594 227944 325666
rect 232502 318880 232558 318889
rect 232502 318815 232558 318824
rect 232516 305658 232544 318815
rect 232504 305652 232556 305658
rect 232504 305594 232556 305600
rect 228916 303748 228968 303754
rect 228916 303690 228968 303696
rect 227916 301566 228298 301594
rect 228928 301580 228956 303690
rect 233896 303686 233924 336806
rect 255964 336796 256016 336802
rect 255964 336738 256016 336744
rect 246304 334008 246356 334014
rect 246304 333950 246356 333956
rect 244924 332648 244976 332654
rect 244924 332590 244976 332596
rect 244188 331356 244240 331362
rect 244188 331298 244240 331304
rect 240138 312216 240194 312225
rect 240138 312151 240194 312160
rect 238024 309256 238076 309262
rect 238024 309198 238076 309204
rect 234618 303784 234674 303793
rect 234618 303719 234674 303728
rect 229560 303680 229612 303686
rect 229560 303622 229612 303628
rect 233884 303680 233936 303686
rect 233884 303622 233936 303628
rect 229572 301580 229600 303622
rect 234632 301580 234660 303719
rect 237840 303680 237892 303686
rect 237840 303622 237892 303628
rect 237852 301580 237880 303622
rect 238036 301594 238064 309198
rect 240048 303680 240100 303686
rect 240046 303648 240048 303657
rect 240100 303648 240102 303657
rect 240046 303583 240102 303592
rect 240152 301594 240180 312151
rect 241060 306400 241112 306406
rect 241060 306342 241112 306348
rect 240690 303648 240746 303657
rect 240690 303583 240692 303592
rect 240744 303583 240746 303592
rect 240692 303554 240744 303560
rect 238036 301566 238510 301594
rect 240152 301566 240442 301594
rect 241072 301580 241100 306342
rect 242990 303648 243046 303657
rect 242990 303583 243046 303592
rect 243004 301580 243032 303583
rect 198738 301472 198794 301481
rect 198794 301430 198950 301458
rect 198738 301407 198794 301416
rect 224774 301336 224830 301345
rect 233790 301336 233846 301345
rect 224830 301294 225078 301322
rect 224774 301271 224830 301280
rect 235630 301336 235686 301345
rect 233846 301294 234002 301322
rect 233790 301271 233846 301280
rect 236918 301336 236974 301345
rect 235686 301294 235934 301322
rect 235630 301271 235686 301280
rect 239494 301336 239550 301345
rect 236974 301294 237222 301322
rect 236918 301271 236974 301280
rect 239550 301294 239798 301322
rect 239494 301271 239550 301280
rect 194230 301200 194286 301209
rect 193312 301164 193364 301170
rect 200578 301200 200634 301209
rect 194286 301158 194442 301186
rect 194230 301135 194286 301144
rect 200634 301158 200882 301186
rect 200578 301135 200634 301144
rect 193312 301106 193364 301112
rect 193324 294642 193352 301106
rect 218426 301064 218482 301073
rect 195440 301034 195730 301050
rect 212000 301034 212382 301050
rect 195428 301028 195730 301034
rect 195480 301022 195730 301028
rect 211988 301028 212382 301034
rect 195428 300970 195480 300976
rect 212040 301022 212382 301028
rect 218482 301022 218730 301050
rect 218426 300999 218482 301008
rect 211988 300970 212040 300976
rect 208860 300960 208912 300966
rect 194690 300928 194746 300937
rect 193416 300886 193890 300914
rect 193312 294636 193364 294642
rect 193312 294578 193364 294584
rect 193416 294522 193444 300886
rect 197358 300928 197414 300937
rect 194746 300886 195086 300914
rect 194690 300863 194746 300872
rect 199290 300928 199346 300937
rect 197414 300886 197662 300914
rect 197358 300863 197414 300872
rect 205638 300928 205694 300937
rect 199346 300886 199594 300914
rect 199290 300863 199346 300872
rect 206282 300928 206338 300937
rect 205694 300886 205942 300914
rect 205638 300863 205694 300872
rect 207110 300928 207166 300937
rect 206338 300886 206586 300914
rect 206282 300863 206338 300872
rect 207166 300886 207230 300914
rect 219440 300960 219492 300966
rect 211526 300928 211582 300937
rect 208912 300908 209162 300914
rect 208860 300902 209162 300908
rect 208872 300886 209162 300902
rect 207110 300863 207166 300872
rect 217046 300928 217102 300937
rect 211582 300886 211738 300914
rect 211526 300863 211582 300872
rect 218978 300928 219034 300937
rect 217102 300886 217442 300914
rect 217046 300863 217102 300872
rect 219438 300928 219440 300937
rect 219492 300928 219494 300937
rect 219034 300886 219374 300914
rect 218978 300863 219034 300872
rect 219438 300863 219494 300872
rect 221646 300928 221702 300937
rect 222382 300928 222438 300937
rect 221702 300886 221950 300914
rect 221646 300863 221702 300872
rect 224130 300928 224186 300937
rect 222438 300886 222594 300914
rect 223882 300886 224130 300914
rect 222382 300863 222438 300872
rect 225970 300928 226026 300937
rect 225722 300886 225970 300914
rect 224130 300863 224186 300872
rect 226522 300928 226578 300937
rect 226366 300886 226522 300914
rect 225970 300863 226026 300872
rect 226522 300863 226578 300872
rect 227258 300928 227314 300937
rect 229834 300928 229890 300937
rect 227314 300886 227654 300914
rect 227258 300863 227314 300872
rect 230570 300928 230626 300937
rect 229890 300886 230230 300914
rect 229834 300863 229890 300872
rect 231214 300928 231270 300937
rect 230626 300886 230874 300914
rect 230570 300863 230626 300872
rect 232042 300928 232098 300937
rect 231270 300886 231518 300914
rect 231214 300863 231270 300872
rect 232502 300928 232558 300937
rect 232098 300886 232162 300914
rect 232042 300863 232098 300872
rect 233330 300928 233386 300937
rect 232558 300886 232806 300914
rect 232502 300863 232558 300872
rect 234986 300928 235042 300937
rect 233386 300886 233450 300914
rect 233330 300863 233386 300872
rect 236642 300928 236698 300937
rect 235042 300886 235290 300914
rect 236578 300886 236642 300914
rect 234986 300863 235042 300872
rect 236642 300863 236698 300872
rect 238850 300928 238906 300937
rect 241426 300928 241482 300937
rect 238906 300886 239154 300914
rect 238850 300863 238906 300872
rect 241978 300928 242034 300937
rect 241482 300886 241730 300914
rect 241426 300863 241482 300872
rect 243266 300928 243322 300937
rect 242034 300886 242374 300914
rect 241978 300863 242034 300872
rect 244200 300914 244228 331298
rect 244936 307057 244964 332590
rect 245016 321700 245068 321706
rect 245016 321642 245068 321648
rect 244922 307048 244978 307057
rect 244922 306983 244978 306992
rect 245028 302938 245056 321642
rect 246316 304298 246344 333950
rect 250444 328568 250496 328574
rect 250444 328510 250496 328516
rect 249064 325780 249116 325786
rect 249064 325722 249116 325728
rect 247684 314696 247736 314702
rect 247684 314638 247736 314644
rect 246304 304292 246356 304298
rect 246304 304234 246356 304240
rect 246118 304056 246174 304065
rect 246118 303991 246174 304000
rect 245016 302932 245068 302938
rect 245016 302874 245068 302880
rect 246132 301580 246160 303991
rect 247408 303612 247460 303618
rect 247408 303554 247460 303560
rect 247420 301580 247448 303554
rect 247696 302841 247724 314638
rect 247682 302832 247738 302841
rect 247682 302767 247738 302776
rect 248510 302560 248566 302569
rect 248510 302495 248566 302504
rect 244554 301064 244610 301073
rect 244610 301022 244858 301050
rect 244554 300999 244610 301008
rect 244280 300960 244332 300966
rect 243322 300886 243662 300914
rect 244200 300908 244280 300914
rect 248524 300937 248552 302495
rect 249076 301918 249104 325722
rect 249154 316704 249210 316713
rect 249154 316639 249210 316648
rect 249168 304201 249196 316639
rect 249154 304192 249210 304201
rect 249154 304127 249210 304136
rect 250456 304094 250484 328510
rect 251824 327752 251876 327758
rect 251824 327694 251876 327700
rect 250536 316056 250588 316062
rect 250536 315998 250588 316004
rect 250444 304088 250496 304094
rect 250444 304030 250496 304036
rect 249338 303920 249394 303929
rect 249338 303855 249394 303864
rect 249064 301912 249116 301918
rect 249064 301854 249116 301860
rect 249352 301580 249380 303855
rect 249982 303648 250038 303657
rect 249982 303583 250038 303592
rect 249996 301580 250024 303583
rect 250548 302462 250576 315998
rect 251272 304292 251324 304298
rect 251272 304234 251324 304240
rect 250628 303680 250680 303686
rect 250628 303622 250680 303628
rect 250536 302456 250588 302462
rect 250536 302398 250588 302404
rect 250640 301580 250668 303622
rect 251284 301580 251312 304234
rect 251836 301753 251864 327694
rect 252744 324964 252796 324970
rect 252744 324906 252796 324912
rect 251916 319456 251968 319462
rect 251916 319398 251968 319404
rect 251928 302297 251956 319398
rect 252756 303090 252784 324906
rect 254216 321632 254268 321638
rect 254216 321574 254268 321580
rect 252836 313336 252888 313342
rect 252836 313278 252888 313284
rect 252848 303226 252876 313278
rect 254030 312080 254086 312089
rect 254030 312015 254086 312024
rect 253940 304088 253992 304094
rect 253940 304030 253992 304036
rect 252848 303198 253152 303226
rect 252756 303062 253060 303090
rect 252744 302932 252796 302938
rect 252744 302874 252796 302880
rect 251914 302288 251970 302297
rect 251914 302223 251970 302232
rect 251822 301744 251878 301753
rect 251822 301679 251878 301688
rect 244200 300902 244332 300908
rect 245106 300928 245162 300937
rect 244200 300900 244320 300902
rect 244214 300886 244320 300900
rect 243266 300863 243322 300872
rect 246394 300928 246450 300937
rect 245162 300886 245502 300914
rect 245106 300863 245162 300872
rect 247774 300928 247830 300937
rect 246450 300886 246790 300914
rect 246394 300863 246450 300872
rect 248510 300928 248566 300937
rect 247830 300886 248078 300914
rect 247774 300863 247830 300872
rect 251546 300928 251602 300937
rect 248566 300886 248722 300914
rect 248510 300863 248566 300872
rect 252466 300928 252522 300937
rect 251602 300886 251942 300914
rect 251546 300863 251602 300872
rect 252522 300886 252586 300914
rect 252466 300863 252522 300872
rect 252756 299962 252784 302874
rect 252926 300656 252982 300665
rect 252926 300591 252982 300600
rect 252940 300150 252968 300591
rect 252928 300144 252980 300150
rect 252928 300086 252980 300092
rect 252756 299934 252968 299962
rect 252836 299872 252888 299878
rect 252836 299814 252888 299820
rect 193232 294494 193444 294522
rect 192576 293276 192628 293282
rect 192576 293218 192628 293224
rect 191378 293176 191434 293185
rect 191378 293111 191434 293120
rect 193126 292904 193182 292913
rect 193126 292839 193182 292848
rect 193140 292602 193168 292839
rect 193128 292596 193180 292602
rect 193128 292538 193180 292544
rect 191746 288280 191802 288289
rect 191746 288215 191802 288224
rect 191286 287736 191342 287745
rect 191286 287671 191342 287680
rect 191760 287094 191788 288215
rect 191748 287088 191800 287094
rect 191748 287030 191800 287036
rect 191654 285968 191710 285977
rect 191654 285903 191710 285912
rect 191194 284880 191250 284889
rect 191194 284815 191250 284824
rect 191562 284744 191618 284753
rect 191562 284679 191618 284688
rect 191576 284442 191604 284679
rect 191564 284436 191616 284442
rect 191564 284378 191616 284384
rect 191668 280650 191696 285903
rect 192392 282872 192444 282878
rect 192392 282814 192444 282820
rect 192404 282441 192432 282814
rect 192390 282432 192446 282441
rect 192390 282367 192446 282376
rect 193034 282432 193090 282441
rect 193034 282367 193090 282376
rect 191746 281344 191802 281353
rect 191746 281279 191802 281288
rect 191760 280838 191788 281279
rect 191748 280832 191800 280838
rect 191748 280774 191800 280780
rect 191668 280622 191788 280650
rect 191654 277808 191710 277817
rect 191654 277743 191710 277752
rect 191668 277438 191696 277743
rect 191656 277432 191708 277438
rect 191656 277374 191708 277380
rect 191654 274408 191710 274417
rect 191654 274343 191710 274352
rect 191668 273290 191696 274343
rect 191656 273284 191708 273290
rect 191656 273226 191708 273232
rect 191562 273184 191618 273193
rect 191562 273119 191618 273128
rect 191576 271930 191604 273119
rect 191654 272096 191710 272105
rect 191654 272031 191710 272040
rect 191668 271998 191696 272031
rect 191656 271992 191708 271998
rect 191656 271934 191708 271940
rect 191564 271924 191616 271930
rect 191564 271866 191616 271872
rect 191654 269784 191710 269793
rect 191654 269719 191710 269728
rect 191668 269142 191696 269719
rect 191656 269136 191708 269142
rect 191656 269078 191708 269084
rect 191654 268696 191710 268705
rect 191654 268631 191710 268640
rect 191668 267782 191696 268631
rect 191656 267776 191708 267782
rect 191656 267718 191708 267724
rect 191286 267472 191342 267481
rect 191286 267407 191342 267416
rect 191300 266422 191328 267407
rect 191288 266416 191340 266422
rect 191288 266358 191340 266364
rect 191562 265160 191618 265169
rect 191562 265095 191618 265104
rect 191576 264994 191604 265095
rect 191564 264988 191616 264994
rect 191564 264930 191616 264936
rect 191654 262848 191710 262857
rect 191654 262783 191710 262792
rect 191668 262342 191696 262783
rect 191656 262336 191708 262342
rect 191656 262278 191708 262284
rect 191196 262268 191248 262274
rect 191196 262210 191248 262216
rect 191208 230450 191236 262210
rect 191654 261760 191710 261769
rect 191654 261695 191710 261704
rect 191668 260914 191696 261695
rect 191656 260908 191708 260914
rect 191656 260850 191708 260856
rect 191286 260536 191342 260545
rect 191286 260471 191342 260480
rect 191300 259486 191328 260471
rect 191288 259480 191340 259486
rect 191288 259422 191340 259428
rect 191654 257136 191710 257145
rect 191654 257071 191710 257080
rect 191668 256766 191696 257071
rect 191656 256760 191708 256766
rect 191656 256702 191708 256708
rect 191654 254824 191710 254833
rect 191654 254759 191710 254768
rect 191668 253978 191696 254759
rect 191656 253972 191708 253978
rect 191656 253914 191708 253920
rect 191654 253600 191710 253609
rect 191654 253535 191710 253544
rect 191668 252618 191696 253535
rect 191656 252612 191708 252618
rect 191656 252554 191708 252560
rect 191654 252512 191710 252521
rect 191654 252447 191710 252456
rect 191668 251258 191696 252447
rect 191656 251252 191708 251258
rect 191656 251194 191708 251200
rect 191654 250200 191710 250209
rect 191654 250135 191710 250144
rect 191668 249830 191696 250135
rect 191656 249824 191708 249830
rect 191656 249766 191708 249772
rect 191654 248976 191710 248985
rect 191654 248911 191710 248920
rect 191668 248470 191696 248911
rect 191656 248464 191708 248470
rect 191656 248406 191708 248412
rect 191654 247888 191710 247897
rect 191654 247823 191710 247832
rect 191668 247110 191696 247823
rect 191656 247104 191708 247110
rect 191656 247046 191708 247052
rect 191196 230444 191248 230450
rect 191196 230386 191248 230392
rect 191562 148472 191618 148481
rect 191562 148407 191618 148416
rect 191576 138281 191604 148407
rect 191654 148336 191710 148345
rect 191654 148271 191710 148280
rect 191562 138272 191618 138281
rect 191562 138207 191618 138216
rect 191564 136604 191616 136610
rect 191564 136546 191616 136552
rect 191576 136377 191604 136546
rect 191562 136368 191618 136377
rect 191562 136303 191618 136312
rect 191562 135552 191618 135561
rect 191562 135487 191618 135496
rect 191576 135318 191604 135487
rect 191564 135312 191616 135318
rect 191564 135254 191616 135260
rect 191116 132466 191236 132494
rect 190366 129840 190422 129849
rect 190366 129775 190422 129784
rect 188896 126948 188948 126954
rect 188896 126890 188948 126896
rect 190380 125526 190408 129775
rect 190368 125520 190420 125526
rect 190368 125462 190420 125468
rect 190644 124092 190696 124098
rect 190644 124034 190696 124040
rect 190656 123049 190684 124034
rect 190642 123040 190698 123049
rect 190642 122975 190698 122984
rect 191102 120320 191158 120329
rect 191102 120255 191158 120264
rect 190366 120184 190422 120193
rect 188988 120148 189040 120154
rect 190366 120119 190422 120128
rect 188988 120090 189040 120096
rect 188344 120080 188396 120086
rect 188344 120022 188396 120028
rect 189000 117473 189028 120090
rect 188986 117464 189042 117473
rect 188986 117399 189042 117408
rect 190380 117201 190408 120119
rect 191116 118697 191144 120255
rect 191102 118688 191158 118697
rect 191102 118623 191158 118632
rect 190366 117192 190422 117201
rect 190366 117127 190422 117136
rect 190642 116784 190698 116793
rect 190642 116719 190698 116728
rect 190656 116074 190684 116719
rect 188436 116068 188488 116074
rect 188436 116010 188488 116016
rect 190644 116068 190696 116074
rect 190644 116010 190696 116016
rect 188252 113212 188304 113218
rect 188252 113154 188304 113160
rect 187700 110492 187752 110498
rect 187700 110434 187752 110440
rect 187712 109002 187740 110434
rect 188264 109750 188292 113154
rect 188252 109744 188304 109750
rect 188252 109686 188304 109692
rect 187700 108996 187752 109002
rect 187700 108938 187752 108944
rect 187608 107840 187660 107846
rect 187608 107782 187660 107788
rect 188344 102196 188396 102202
rect 188344 102138 188396 102144
rect 187700 101448 187752 101454
rect 187700 101390 187752 101396
rect 187712 101046 187740 101390
rect 187700 101040 187752 101046
rect 187700 100982 187752 100988
rect 187146 78568 187202 78577
rect 187146 78503 187202 78512
rect 187056 74520 187108 74526
rect 187056 74462 187108 74468
rect 188356 73137 188384 102138
rect 188448 97306 188476 116010
rect 190366 113520 190422 113529
rect 190366 113455 190422 113464
rect 190380 110906 190408 113455
rect 191010 113248 191066 113257
rect 191010 113183 191012 113192
rect 191064 113183 191066 113192
rect 191012 113154 191064 113160
rect 190368 110900 190420 110906
rect 190368 110842 190420 110848
rect 190366 110800 190422 110809
rect 190366 110735 190422 110744
rect 190380 109041 190408 110735
rect 190366 109032 190422 109041
rect 190366 108967 190422 108976
rect 189080 107840 189132 107846
rect 189080 107782 189132 107788
rect 188988 101040 189040 101046
rect 188988 100982 189040 100988
rect 188528 98116 188580 98122
rect 188528 98058 188580 98064
rect 188436 97300 188488 97306
rect 188436 97242 188488 97248
rect 188436 94512 188488 94518
rect 188436 94454 188488 94460
rect 188448 86970 188476 94454
rect 188540 92478 188568 98058
rect 188528 92472 188580 92478
rect 188528 92414 188580 92420
rect 188436 86964 188488 86970
rect 188436 86906 188488 86912
rect 188342 73128 188398 73137
rect 188342 73063 188398 73072
rect 189000 49026 189028 100982
rect 189092 82793 189120 107782
rect 190460 105664 190512 105670
rect 190460 105606 190512 105612
rect 190472 105097 190500 105606
rect 190458 105088 190514 105097
rect 190458 105023 190514 105032
rect 190472 104802 190500 105023
rect 190380 104774 190500 104802
rect 189078 82784 189134 82793
rect 189078 82719 189134 82728
rect 189092 81569 189120 82719
rect 189078 81560 189134 81569
rect 189078 81495 189134 81504
rect 189722 81560 189778 81569
rect 189722 81495 189778 81504
rect 188988 49020 189040 49026
rect 188988 48962 189040 48968
rect 189736 46918 189764 81495
rect 190380 69698 190408 104774
rect 191010 103456 191066 103465
rect 191010 103391 191066 103400
rect 191024 102202 191052 103391
rect 191012 102196 191064 102202
rect 191012 102138 191064 102144
rect 190642 101552 190698 101561
rect 190642 101487 190698 101496
rect 190656 101046 190684 101487
rect 190644 101040 190696 101046
rect 190644 100982 190696 100988
rect 190644 100700 190696 100706
rect 190644 100642 190696 100648
rect 190656 99929 190684 100642
rect 190642 99920 190698 99929
rect 190642 99855 190698 99864
rect 190826 98832 190882 98841
rect 190826 98767 190882 98776
rect 190840 98054 190868 98767
rect 190828 98048 190880 98054
rect 190828 97990 190880 97996
rect 191116 80714 191144 118623
rect 191208 117473 191236 132466
rect 191668 132394 191696 148271
rect 191656 132388 191708 132394
rect 191656 132330 191708 132336
rect 191668 132025 191696 132330
rect 191654 132016 191710 132025
rect 191654 131951 191710 131960
rect 191654 129296 191710 129305
rect 191654 129231 191710 129240
rect 191668 128382 191696 129231
rect 191656 128376 191708 128382
rect 191656 128318 191708 128324
rect 191656 126948 191708 126954
rect 191656 126890 191708 126896
rect 191668 126585 191696 126890
rect 191654 126576 191710 126585
rect 191654 126511 191710 126520
rect 191654 123856 191710 123865
rect 191654 123791 191710 123800
rect 191668 122874 191696 123791
rect 191656 122868 191708 122874
rect 191656 122810 191708 122816
rect 191654 122224 191710 122233
rect 191654 122159 191710 122168
rect 191668 122126 191696 122159
rect 191656 122120 191708 122126
rect 191656 122062 191708 122068
rect 191562 121408 191618 121417
rect 191562 121343 191618 121352
rect 191576 120193 191604 121343
rect 191562 120184 191618 120193
rect 191562 120119 191618 120128
rect 191656 120080 191708 120086
rect 191656 120022 191708 120028
rect 191668 119513 191696 120022
rect 191654 119504 191710 119513
rect 191654 119439 191710 119448
rect 191194 117464 191250 117473
rect 191194 117399 191250 117408
rect 191656 117292 191708 117298
rect 191656 117234 191708 117240
rect 191668 115977 191696 117234
rect 191654 115968 191710 115977
rect 191654 115903 191710 115912
rect 191760 113174 191788 280622
rect 192576 250504 192628 250510
rect 192576 250446 192628 250452
rect 192484 248532 192536 248538
rect 192484 248474 192536 248480
rect 192496 228857 192524 248474
rect 192588 235958 192616 250446
rect 193048 238202 193076 282367
rect 193036 238196 193088 238202
rect 193036 238138 193088 238144
rect 192576 235952 192628 235958
rect 192576 235894 192628 235900
rect 192482 228848 192538 228857
rect 192482 228783 192538 228792
rect 191838 211168 191894 211177
rect 191838 211103 191894 211112
rect 191852 209710 191880 211103
rect 191840 209704 191892 209710
rect 191840 209646 191892 209652
rect 193140 206310 193168 292538
rect 193232 292534 193260 294494
rect 193220 292528 193272 292534
rect 193220 292470 193272 292476
rect 193218 290592 193274 290601
rect 193218 290527 193274 290536
rect 193232 289882 193260 290527
rect 193220 289876 193272 289882
rect 193220 289818 193272 289824
rect 193232 236706 193260 289818
rect 252848 281353 252876 299814
rect 252940 289785 252968 299934
rect 253032 290193 253060 303062
rect 253124 299878 253152 303198
rect 253478 301064 253534 301073
rect 253230 301022 253478 301050
rect 253478 300999 253534 301008
rect 253112 299872 253164 299878
rect 253112 299814 253164 299820
rect 253952 296449 253980 304030
rect 253938 296440 253994 296449
rect 253938 296375 253994 296384
rect 253938 293856 253994 293865
rect 253938 293791 253994 293800
rect 253018 290184 253074 290193
rect 253018 290119 253074 290128
rect 252926 289776 252982 289785
rect 252926 289711 252982 289720
rect 252834 281344 252890 281353
rect 252834 281279 252890 281288
rect 252834 274816 252890 274825
rect 252834 274751 252890 274760
rect 252848 267734 252876 274751
rect 252848 267706 253060 267734
rect 252926 267336 252982 267345
rect 252926 267271 252982 267280
rect 252940 264330 252968 267271
rect 252756 264302 252968 264330
rect 193402 258904 193458 258913
rect 193402 258839 193458 258848
rect 193416 258058 193444 258839
rect 193404 258052 193456 258058
rect 193404 257994 193456 258000
rect 193680 246356 193732 246362
rect 193680 246298 193732 246304
rect 193586 242856 193642 242865
rect 193586 242791 193642 242800
rect 193600 241670 193628 242791
rect 193692 241754 193720 246298
rect 193692 241726 194350 241754
rect 193588 241664 193640 241670
rect 193588 241606 193640 241612
rect 193692 238754 193720 241726
rect 193772 241664 193824 241670
rect 193772 241606 193824 241612
rect 195244 241664 195296 241670
rect 195244 241606 195296 241612
rect 195612 241664 195664 241670
rect 249064 241664 249116 241670
rect 195664 241612 195914 241618
rect 195612 241606 195914 241612
rect 193324 238726 193720 238754
rect 193220 236700 193272 236706
rect 193220 236642 193272 236648
rect 193128 206304 193180 206310
rect 193128 206246 193180 206252
rect 193324 195362 193352 238726
rect 193784 224369 193812 241606
rect 195256 237969 195284 241606
rect 195624 241590 195914 241606
rect 196624 241596 196676 241602
rect 196624 241538 196676 241544
rect 195978 241496 196034 241505
rect 195978 241431 196034 241440
rect 195242 237960 195298 237969
rect 195242 237895 195298 237904
rect 195242 235512 195298 235521
rect 195242 235447 195298 235456
rect 195152 235272 195204 235278
rect 195152 235214 195204 235220
rect 195164 229094 195192 235214
rect 195256 234666 195284 235447
rect 195244 234660 195296 234666
rect 195244 234602 195296 234608
rect 195164 229066 195284 229094
rect 193770 224360 193826 224369
rect 193770 224295 193826 224304
rect 193312 195356 193364 195362
rect 193312 195298 193364 195304
rect 192484 182844 192536 182850
rect 192484 182786 192536 182792
rect 192496 164898 192524 182786
rect 193862 181384 193918 181393
rect 193862 181319 193918 181328
rect 193036 167748 193088 167754
rect 193036 167690 193088 167696
rect 192484 164892 192536 164898
rect 192484 164834 192536 164840
rect 192496 127673 192524 164834
rect 192576 144968 192628 144974
rect 192576 144910 192628 144916
rect 192588 137902 192616 144910
rect 192576 137896 192628 137902
rect 192576 137838 192628 137844
rect 192850 137456 192906 137465
rect 192850 137391 192906 137400
rect 192864 135250 192892 137391
rect 192852 135244 192904 135250
rect 192852 135186 192904 135192
rect 192482 127664 192538 127673
rect 192482 127599 192538 127608
rect 191668 113146 191788 113174
rect 191562 109712 191618 109721
rect 191562 109647 191618 109656
rect 191576 109070 191604 109647
rect 191564 109064 191616 109070
rect 191564 109006 191616 109012
rect 191564 107636 191616 107642
rect 191564 107578 191616 107584
rect 191576 107001 191604 107578
rect 191562 106992 191618 107001
rect 191562 106927 191618 106936
rect 191668 104281 191696 113146
rect 191748 112464 191800 112470
rect 191746 112432 191748 112441
rect 191800 112432 191802 112441
rect 191746 112367 191802 112376
rect 191746 110528 191802 110537
rect 191746 110463 191748 110472
rect 191800 110463 191802 110472
rect 191748 110434 191800 110440
rect 191748 107840 191800 107846
rect 191746 107808 191748 107817
rect 191800 107808 191802 107817
rect 191746 107743 191802 107752
rect 191746 106176 191802 106185
rect 191746 106111 191802 106120
rect 191760 105942 191788 106111
rect 191748 105936 191800 105942
rect 191748 105878 191800 105884
rect 191654 104272 191710 104281
rect 191654 104207 191710 104216
rect 191668 104174 191696 104207
rect 191656 104168 191708 104174
rect 191656 104110 191708 104116
rect 191654 100736 191710 100745
rect 191654 100671 191710 100680
rect 191668 97866 191696 100671
rect 191748 98116 191800 98122
rect 191748 98058 191800 98064
rect 191760 98025 191788 98058
rect 191746 98016 191802 98025
rect 191746 97951 191802 97960
rect 191668 97838 191788 97866
rect 191562 96384 191618 96393
rect 191562 96319 191618 96328
rect 191576 95946 191604 96319
rect 191564 95940 191616 95946
rect 191564 95882 191616 95888
rect 191654 94480 191710 94489
rect 191654 94415 191710 94424
rect 191668 93906 191696 94415
rect 191656 93900 191708 93906
rect 191656 93842 191708 93848
rect 191760 82890 191788 97838
rect 191840 95260 191892 95266
rect 191840 95202 191892 95208
rect 191852 92177 191880 95202
rect 191838 92168 191894 92177
rect 191838 92103 191894 92112
rect 192864 83473 192892 135186
rect 193048 134745 193076 167690
rect 193876 161474 193904 181319
rect 195256 180130 195284 229066
rect 195888 188352 195940 188358
rect 195888 188294 195940 188300
rect 195244 180124 195296 180130
rect 195244 180066 195296 180072
rect 195900 175370 195928 188294
rect 195244 175364 195296 175370
rect 195244 175306 195296 175312
rect 195888 175364 195940 175370
rect 195888 175306 195940 175312
rect 195060 166388 195112 166394
rect 195060 166330 195112 166336
rect 195072 165646 195100 166330
rect 194600 165640 194652 165646
rect 194600 165582 194652 165588
rect 195060 165640 195112 165646
rect 195060 165582 195112 165588
rect 193416 161446 193904 161474
rect 193416 160857 193444 161446
rect 193402 160848 193458 160857
rect 193402 160783 193458 160792
rect 193126 144120 193182 144129
rect 193126 144055 193182 144064
rect 193034 134736 193090 134745
rect 193034 134671 193090 134680
rect 193048 133958 193076 134671
rect 193036 133952 193088 133958
rect 193036 133894 193088 133900
rect 193140 128489 193168 144055
rect 193416 139641 193444 160783
rect 194612 151814 194640 165582
rect 194612 151786 195008 151814
rect 193496 147008 193548 147014
rect 193496 146950 193548 146956
rect 193402 139632 193458 139641
rect 193402 139567 193458 139576
rect 193126 128480 193182 128489
rect 193126 128415 193182 128424
rect 192942 127664 192998 127673
rect 192942 127599 192998 127608
rect 192850 83464 192906 83473
rect 192850 83399 192906 83408
rect 191748 82884 191800 82890
rect 191748 82826 191800 82832
rect 191104 80708 191156 80714
rect 191104 80650 191156 80656
rect 191760 80034 191788 82826
rect 191748 80028 191800 80034
rect 191748 79970 191800 79976
rect 190460 75200 190512 75206
rect 190460 75142 190512 75148
rect 190368 69692 190420 69698
rect 190368 69634 190420 69640
rect 190472 68950 190500 75142
rect 192956 71058 192984 127599
rect 193036 92472 193088 92478
rect 193036 92414 193088 92420
rect 193048 92313 193076 92414
rect 193034 92304 193090 92313
rect 193034 92239 193090 92248
rect 193034 91216 193090 91225
rect 193034 91151 193090 91160
rect 191104 71052 191156 71058
rect 191104 70994 191156 71000
rect 192944 71052 192996 71058
rect 192944 70994 192996 71000
rect 190460 68944 190512 68950
rect 190460 68886 190512 68892
rect 189724 46912 189776 46918
rect 189724 46854 189776 46860
rect 186964 40724 187016 40730
rect 186964 40666 187016 40672
rect 183468 29640 183520 29646
rect 183468 29582 183520 29588
rect 191116 21418 191144 70994
rect 193048 33794 193076 91151
rect 193140 68338 193168 128415
rect 193508 103514 193536 146950
rect 193772 145036 193824 145042
rect 193772 144978 193824 144984
rect 193588 144220 193640 144226
rect 193588 144162 193640 144168
rect 193600 140964 193628 144162
rect 193784 140978 193812 144978
rect 194690 143440 194746 143449
rect 194690 143375 194746 143384
rect 194704 142225 194732 143375
rect 194690 142216 194746 142225
rect 194690 142151 194746 142160
rect 193784 140950 194166 140978
rect 194704 140964 194732 142151
rect 194980 140978 195008 151786
rect 195256 143449 195284 175306
rect 195992 172378 196020 241431
rect 196636 235249 196664 241538
rect 197556 240106 197584 241604
rect 199120 241398 199148 241604
rect 199108 241392 199160 241398
rect 199108 241334 199160 241340
rect 198646 240272 198702 240281
rect 198646 240207 198702 240216
rect 197544 240100 197596 240106
rect 197544 240042 197596 240048
rect 198004 240100 198056 240106
rect 198004 240042 198056 240048
rect 196622 235240 196678 235249
rect 196622 235175 196678 235184
rect 196622 221504 196678 221513
rect 196622 221439 196678 221448
rect 195980 172372 196032 172378
rect 195980 172314 196032 172320
rect 196636 164937 196664 221439
rect 198016 185638 198044 240042
rect 198096 216028 198148 216034
rect 198096 215970 198148 215976
rect 198004 185632 198056 185638
rect 198004 185574 198056 185580
rect 198002 175400 198058 175409
rect 198002 175335 198058 175344
rect 196808 172372 196860 172378
rect 196808 172314 196860 172320
rect 196820 171154 196848 172314
rect 196808 171148 196860 171154
rect 196808 171090 196860 171096
rect 196716 170468 196768 170474
rect 196716 170410 196768 170416
rect 196622 164928 196678 164937
rect 196622 164863 196678 164872
rect 196070 159352 196126 159361
rect 196070 159287 196126 159296
rect 196084 158778 196112 159287
rect 196072 158772 196124 158778
rect 196072 158714 196124 158720
rect 196728 147257 196756 170410
rect 196820 149734 196848 171090
rect 197360 166116 197412 166122
rect 197360 166058 197412 166064
rect 197372 165714 197400 166058
rect 197360 165708 197412 165714
rect 197360 165650 197412 165656
rect 196898 159352 196954 159361
rect 196898 159287 196954 159296
rect 196808 149728 196860 149734
rect 196808 149670 196860 149676
rect 196714 147248 196770 147257
rect 196714 147183 196770 147192
rect 196530 145752 196586 145761
rect 196530 145687 196586 145696
rect 195242 143440 195298 143449
rect 195242 143375 195298 143384
rect 195978 142216 196034 142225
rect 195978 142151 196034 142160
rect 194980 140950 195454 140978
rect 195992 140964 196020 142151
rect 196544 140964 196572 145687
rect 196912 142225 196940 159287
rect 197084 145648 197136 145654
rect 197084 145590 197136 145596
rect 197096 142361 197124 145590
rect 197082 142352 197138 142361
rect 197082 142287 197138 142296
rect 196898 142216 196954 142225
rect 196898 142151 196954 142160
rect 197096 140964 197124 142287
rect 197372 140978 197400 165650
rect 197910 148608 197966 148617
rect 197910 148543 197966 148552
rect 197924 140978 197952 148543
rect 198016 143449 198044 175335
rect 198108 166122 198136 215970
rect 198096 166116 198148 166122
rect 198096 166058 198148 166064
rect 198660 154737 198688 240207
rect 198832 238196 198884 238202
rect 198832 238138 198884 238144
rect 198740 164892 198792 164898
rect 198740 164834 198792 164840
rect 198752 162926 198780 164834
rect 198740 162920 198792 162926
rect 198740 162862 198792 162868
rect 198094 154728 198150 154737
rect 198094 154663 198150 154672
rect 198646 154728 198702 154737
rect 198646 154663 198702 154672
rect 198108 149705 198136 154663
rect 198094 149696 198150 149705
rect 198094 149631 198150 149640
rect 198752 143562 198780 162862
rect 198844 143721 198872 238138
rect 200776 235958 200804 241604
rect 202432 239426 202460 241604
rect 202420 239420 202472 239426
rect 202420 239362 202472 239368
rect 203996 236609 204024 241604
rect 204904 238060 204956 238066
rect 204904 238002 204956 238008
rect 203982 236600 204038 236609
rect 203982 236535 204038 236544
rect 200120 235952 200172 235958
rect 200120 235894 200172 235900
rect 200764 235952 200816 235958
rect 200764 235894 200816 235900
rect 200132 167754 200160 235894
rect 200764 235272 200816 235278
rect 200764 235214 200816 235220
rect 200776 208457 200804 235214
rect 202788 228404 202840 228410
rect 202788 228346 202840 228352
rect 202800 223553 202828 228346
rect 202786 223544 202842 223553
rect 202786 223479 202842 223488
rect 202144 221536 202196 221542
rect 202144 221478 202196 221484
rect 200762 208448 200818 208457
rect 200762 208383 200818 208392
rect 202156 168473 202184 221478
rect 202236 221468 202288 221474
rect 202236 221410 202288 221416
rect 202248 211818 202276 221410
rect 202236 211812 202288 211818
rect 202236 211754 202288 211760
rect 202880 174548 202932 174554
rect 202880 174490 202932 174496
rect 202892 173194 202920 174490
rect 202880 173188 202932 173194
rect 202880 173130 202932 173136
rect 201498 168464 201554 168473
rect 201498 168399 201554 168408
rect 202142 168464 202198 168473
rect 202142 168399 202198 168408
rect 200120 167748 200172 167754
rect 200120 167690 200172 167696
rect 201512 151814 201540 168399
rect 201512 151786 201632 151814
rect 201406 145752 201462 145761
rect 201406 145687 201462 145696
rect 200210 144256 200266 144265
rect 200210 144191 200266 144200
rect 198830 143712 198886 143721
rect 198830 143647 198886 143656
rect 198752 143534 199240 143562
rect 198002 143440 198058 143449
rect 198002 143375 198058 143384
rect 198922 143440 198978 143449
rect 198922 143375 198978 143384
rect 198646 141128 198702 141137
rect 198646 141063 198702 141072
rect 197372 140950 197846 140978
rect 197924 140950 198398 140978
rect 198660 140554 198688 141063
rect 198936 140964 198964 143375
rect 199212 140978 199240 143534
rect 199212 140950 199686 140978
rect 200224 140964 200252 144191
rect 201314 143576 201370 143585
rect 201314 143511 201370 143520
rect 200764 141432 200816 141438
rect 200764 141374 200816 141380
rect 200776 140964 200804 141374
rect 201328 140964 201356 143511
rect 201420 142225 201448 145687
rect 201406 142216 201462 142225
rect 201406 142151 201462 142160
rect 201604 140978 201632 151786
rect 202144 147756 202196 147762
rect 202144 147698 202196 147704
rect 202156 140978 202184 147698
rect 202892 140978 202920 173130
rect 204916 170406 204944 238002
rect 205546 235920 205602 235929
rect 205546 235855 205602 235864
rect 205454 171728 205510 171737
rect 205454 171663 205510 171672
rect 204904 170400 204956 170406
rect 204904 170342 204956 170348
rect 204168 163532 204220 163538
rect 204168 163474 204220 163480
rect 201604 140950 202078 140978
rect 202156 140950 202630 140978
rect 202892 140950 203472 140978
rect 203444 140894 203472 140950
rect 203432 140888 203484 140894
rect 203432 140830 203484 140836
rect 198648 140548 198700 140554
rect 198648 140490 198700 140496
rect 203522 140448 203578 140457
rect 204180 140434 204208 163474
rect 204442 145888 204498 145897
rect 204442 145823 204498 145832
rect 204456 140964 204484 145823
rect 204916 143585 204944 170342
rect 205086 156224 205142 156233
rect 205086 156159 205142 156168
rect 205100 155242 205128 156159
rect 205088 155236 205140 155242
rect 205088 155178 205140 155184
rect 204902 143576 204958 143585
rect 204902 143511 204958 143520
rect 205468 141409 205496 171663
rect 205560 156233 205588 235855
rect 205652 231742 205680 241604
rect 206284 236700 206336 236706
rect 206284 236642 206336 236648
rect 205640 231736 205692 231742
rect 205640 231678 205692 231684
rect 205652 230994 205680 231678
rect 205640 230988 205692 230994
rect 205640 230930 205692 230936
rect 205640 170400 205692 170406
rect 205640 170342 205692 170348
rect 205652 169833 205680 170342
rect 205638 169824 205694 169833
rect 205638 169759 205694 169768
rect 205546 156224 205602 156233
rect 205546 156159 205602 156168
rect 205652 144129 205680 169759
rect 206296 151814 206324 236642
rect 207110 233880 207166 233889
rect 207110 233815 207166 233824
rect 206928 232552 206980 232558
rect 206928 232494 206980 232500
rect 206376 230988 206428 230994
rect 206376 230930 206428 230936
rect 206388 173913 206416 230930
rect 206374 173904 206430 173913
rect 206374 173839 206430 173848
rect 206296 151786 206416 151814
rect 206388 150550 206416 151786
rect 206376 150544 206428 150550
rect 206376 150486 206428 150492
rect 205638 144120 205694 144129
rect 205638 144055 205694 144064
rect 205546 143576 205602 143585
rect 205546 143511 205602 143520
rect 204994 141400 205050 141409
rect 204994 141335 205050 141344
rect 205454 141400 205510 141409
rect 205454 141335 205510 141344
rect 205008 140978 205036 141335
rect 205086 140992 205142 141001
rect 205008 140964 205086 140978
rect 205022 140950 205086 140964
rect 205560 140964 205588 143511
rect 206388 142186 206416 150486
rect 206940 147762 206968 232494
rect 207124 175302 207152 233815
rect 207112 175296 207164 175302
rect 207112 175238 207164 175244
rect 206928 147756 206980 147762
rect 206928 147698 206980 147704
rect 206376 142180 206428 142186
rect 206376 142122 206428 142128
rect 206388 140978 206416 142122
rect 206388 140950 206862 140978
rect 205086 140927 205142 140936
rect 206940 140486 206968 147698
rect 207124 140978 207152 175238
rect 207216 147014 207244 241604
rect 208872 237386 208900 241604
rect 208860 237380 208912 237386
rect 208860 237322 208912 237328
rect 208872 236026 208900 237322
rect 208400 236020 208452 236026
rect 208400 235962 208452 235968
rect 208860 236020 208912 236026
rect 208860 235962 208912 235968
rect 208412 151910 208440 235962
rect 208492 231124 208544 231130
rect 208492 231066 208544 231072
rect 208504 228857 208532 231066
rect 208490 228848 208546 228857
rect 208490 228783 208546 228792
rect 208504 227769 208532 228783
rect 208490 227760 208546 227769
rect 208490 227695 208546 227704
rect 210528 171134 210556 241604
rect 211068 236700 211120 236706
rect 211068 236642 211120 236648
rect 211080 233209 211108 236642
rect 211066 233200 211122 233209
rect 211066 233135 211122 233144
rect 212092 230450 212120 241604
rect 212080 230444 212132 230450
rect 212080 230386 212132 230392
rect 212092 227089 212120 230386
rect 212078 227080 212134 227089
rect 212078 227015 212134 227024
rect 213182 206272 213238 206281
rect 213182 206207 213238 206216
rect 213196 177313 213224 206207
rect 213182 177304 213238 177313
rect 213182 177239 213238 177248
rect 211804 173936 211856 173942
rect 211804 173878 211856 173884
rect 210436 171106 210556 171134
rect 210436 167686 210464 171106
rect 210424 167680 210476 167686
rect 210424 167622 210476 167628
rect 208584 159384 208636 159390
rect 208584 159326 208636 159332
rect 208596 157418 208624 159326
rect 208584 157412 208636 157418
rect 208584 157354 208636 157360
rect 208400 151904 208452 151910
rect 208400 151846 208452 151852
rect 208412 151094 208440 151846
rect 208596 151814 208624 157354
rect 209044 152516 209096 152522
rect 209044 152458 209096 152464
rect 208596 151786 208808 151814
rect 208400 151088 208452 151094
rect 208400 151030 208452 151036
rect 208400 150476 208452 150482
rect 208400 150418 208452 150424
rect 208412 150385 208440 150418
rect 208398 150376 208454 150385
rect 208398 150311 208454 150320
rect 207204 147008 207256 147014
rect 207204 146950 207256 146956
rect 208124 143540 208176 143546
rect 208124 143482 208176 143488
rect 207124 140950 207414 140978
rect 208136 140842 208164 143482
rect 208412 142154 208440 150311
rect 208412 142126 208532 142154
rect 208504 140978 208532 142126
rect 208780 140978 208808 151786
rect 209056 143546 209084 152458
rect 209780 149728 209832 149734
rect 209780 149670 209832 149676
rect 209044 143540 209096 143546
rect 209044 143482 209096 143488
rect 208504 140950 208702 140978
rect 208780 140950 209254 140978
rect 207768 140828 208164 140842
rect 207768 140826 208150 140828
rect 207756 140820 208150 140826
rect 207808 140814 208150 140820
rect 207756 140762 207808 140768
rect 209792 140570 209820 149670
rect 210436 149190 210464 167622
rect 211160 159452 211212 159458
rect 211160 159394 211212 159400
rect 210240 149184 210292 149190
rect 210240 149126 210292 149132
rect 210424 149184 210476 149190
rect 210424 149126 210476 149132
rect 210252 148481 210280 149126
rect 210238 148472 210294 148481
rect 210238 148407 210294 148416
rect 210700 147212 210752 147218
rect 210700 147154 210752 147160
rect 210054 146976 210110 146985
rect 210054 146911 210110 146920
rect 210068 140978 210096 146911
rect 210712 140978 210740 147154
rect 211172 140978 211200 159394
rect 211816 155922 211844 173878
rect 211252 155916 211304 155922
rect 211252 155858 211304 155864
rect 211804 155916 211856 155922
rect 211804 155858 211856 155864
rect 211264 151814 211292 155858
rect 211264 151786 211936 151814
rect 211908 140978 211936 151786
rect 213196 142186 213224 177239
rect 213276 161492 213328 161498
rect 213276 161434 213328 161440
rect 213288 146266 213316 161434
rect 213276 146260 213328 146266
rect 213276 146202 213328 146208
rect 213748 145654 213776 241604
rect 215404 240145 215432 241604
rect 215942 240952 215998 240961
rect 215942 240887 215998 240896
rect 215390 240136 215446 240145
rect 215390 240071 215446 240080
rect 214564 203584 214616 203590
rect 214564 203526 214616 203532
rect 214012 177336 214064 177342
rect 214012 177278 214064 177284
rect 213920 162852 213972 162858
rect 213920 162794 213972 162800
rect 213932 161498 213960 162794
rect 213920 161492 213972 161498
rect 213920 161434 213972 161440
rect 213736 145648 213788 145654
rect 213736 145590 213788 145596
rect 213458 142760 213514 142769
rect 213458 142695 213514 142704
rect 213472 142225 213500 142695
rect 213458 142216 213514 142225
rect 213184 142180 213236 142186
rect 212920 142128 213184 142154
rect 213458 142151 213514 142160
rect 212920 142126 213236 142128
rect 210068 140950 210542 140978
rect 210712 140950 211094 140978
rect 211172 140950 211646 140978
rect 211908 140950 212382 140978
rect 212920 140964 212948 142126
rect 213184 142122 213236 142126
rect 213472 140964 213500 142151
rect 213932 140978 213960 161434
rect 214024 147626 214052 177278
rect 214576 174049 214604 203526
rect 214562 174040 214618 174049
rect 214562 173975 214618 173984
rect 214576 162858 214604 173975
rect 215482 167104 215538 167113
rect 215482 167039 215538 167048
rect 214564 162852 214616 162858
rect 214564 162794 214616 162800
rect 214012 147620 214064 147626
rect 214012 147562 214064 147568
rect 214024 147218 214052 147562
rect 214012 147212 214064 147218
rect 214012 147154 214064 147160
rect 215300 142860 215352 142866
rect 215300 142802 215352 142808
rect 214746 141128 214802 141137
rect 214746 141063 214802 141072
rect 214760 140978 214788 141063
rect 213932 140950 214038 140978
rect 214760 140964 215064 140978
rect 215312 140964 215340 142802
rect 215496 140978 215524 167039
rect 215956 152425 215984 240887
rect 216968 233238 216996 241604
rect 216956 233232 217008 233238
rect 216956 233174 217008 233180
rect 217324 232620 217376 232626
rect 217324 232562 217376 232568
rect 216036 222896 216088 222902
rect 216036 222838 216088 222844
rect 216048 167113 216076 222838
rect 217336 192506 217364 232562
rect 218624 231130 218652 241604
rect 218612 231124 218664 231130
rect 218612 231066 218664 231072
rect 217416 196648 217468 196654
rect 217416 196590 217468 196596
rect 217324 192500 217376 192506
rect 217324 192442 217376 192448
rect 217324 178084 217376 178090
rect 217324 178026 217376 178032
rect 216128 176724 216180 176730
rect 216128 176666 216180 176672
rect 216034 167104 216090 167113
rect 216034 167039 216090 167048
rect 215942 152416 215998 152425
rect 215942 152351 215998 152360
rect 216140 142866 216168 176666
rect 216678 157448 216734 157457
rect 216678 157383 216734 157392
rect 216692 151814 216720 157383
rect 216692 151786 216996 151814
rect 216772 149116 216824 149122
rect 216772 149058 216824 149064
rect 216588 146260 216640 146266
rect 216588 146202 216640 146208
rect 216128 142860 216180 142866
rect 216128 142802 216180 142808
rect 214774 140950 215064 140964
rect 215496 140950 215878 140978
rect 216600 140964 216628 146202
rect 216784 140978 216812 149058
rect 216968 147674 216996 151786
rect 216968 147646 217272 147674
rect 217244 140978 217272 147646
rect 217336 142458 217364 178026
rect 217428 170406 217456 196590
rect 220188 182850 220216 241604
rect 221476 241590 221858 241618
rect 221476 238746 221504 241590
rect 223500 240145 223528 241604
rect 224132 240780 224184 240786
rect 224132 240722 224184 240728
rect 222382 240136 222438 240145
rect 222382 240071 222438 240080
rect 223486 240136 223542 240145
rect 223486 240071 223542 240080
rect 221464 238740 221516 238746
rect 221464 238682 221516 238688
rect 221002 234016 221058 234025
rect 221002 233951 221058 233960
rect 220728 233912 220780 233918
rect 220728 233854 220780 233860
rect 220176 182844 220228 182850
rect 220176 182786 220228 182792
rect 218704 180872 218756 180878
rect 218704 180814 218756 180820
rect 217416 170400 217468 170406
rect 217416 170342 217468 170348
rect 217416 166320 217468 166326
rect 217416 166262 217468 166268
rect 217428 157457 217456 166262
rect 217414 157448 217470 157457
rect 217414 157383 217470 157392
rect 217324 142452 217376 142458
rect 217324 142394 217376 142400
rect 218244 142452 218296 142458
rect 218244 142394 218296 142400
rect 218256 140978 218284 142394
rect 216784 140950 217166 140978
rect 217244 140950 217718 140978
rect 218256 140964 218560 140978
rect 218270 140950 218560 140964
rect 215036 140826 215064 140950
rect 215024 140820 215076 140826
rect 215024 140762 215076 140768
rect 209792 140556 210096 140570
rect 209806 140554 210096 140556
rect 209806 140548 210108 140554
rect 209806 140542 210056 140548
rect 210056 140490 210108 140496
rect 218532 140486 218560 140950
rect 218716 140758 218744 180814
rect 218796 179444 218848 179450
rect 218796 179386 218848 179392
rect 218808 141409 218836 179386
rect 220084 156052 220136 156058
rect 220084 155994 220136 156000
rect 218980 145580 219032 145586
rect 218980 145522 219032 145528
rect 218794 141400 218850 141409
rect 218794 141335 218850 141344
rect 218886 140856 218942 140865
rect 218992 140842 219020 145522
rect 219530 142760 219586 142769
rect 219530 142695 219586 142704
rect 219544 140964 219572 142695
rect 220096 142254 220124 155994
rect 220740 152522 220768 233854
rect 221016 230450 221044 233951
rect 221004 230444 221056 230450
rect 221004 230386 221056 230392
rect 220820 215960 220872 215966
rect 220820 215902 220872 215908
rect 220832 172582 220860 215902
rect 220820 172576 220872 172582
rect 220820 172518 220872 172524
rect 220832 171134 220860 172518
rect 220832 171106 221044 171134
rect 220820 164960 220872 164966
rect 220820 164902 220872 164908
rect 220728 152516 220780 152522
rect 220728 152458 220780 152464
rect 220832 147674 220860 164902
rect 220832 147646 220952 147674
rect 220820 146940 220872 146946
rect 220820 146882 220872 146888
rect 220084 142248 220136 142254
rect 220084 142190 220136 142196
rect 220096 140964 220124 142190
rect 220832 140964 220860 146882
rect 220924 140978 220952 147646
rect 221016 142769 221044 171106
rect 221476 167074 221504 238682
rect 222106 238640 222162 238649
rect 222106 238575 222162 238584
rect 222120 237454 222148 238575
rect 222108 237448 222160 237454
rect 222108 237390 222160 237396
rect 222198 172408 222254 172417
rect 222198 172343 222254 172352
rect 222212 171193 222240 172343
rect 222198 171184 222254 171193
rect 222198 171119 222254 171128
rect 221464 167068 221516 167074
rect 221464 167010 221516 167016
rect 222108 167068 222160 167074
rect 222108 167010 222160 167016
rect 222120 166394 222148 167010
rect 222108 166388 222160 166394
rect 222108 166330 222160 166336
rect 221002 142760 221058 142769
rect 221002 142695 221058 142704
rect 222212 140978 222240 171119
rect 222290 162752 222346 162761
rect 222290 162687 222346 162696
rect 222304 161537 222332 162687
rect 222290 161528 222346 161537
rect 222290 161463 222346 161472
rect 222304 156058 222332 161463
rect 222292 156052 222344 156058
rect 222292 155994 222344 156000
rect 222304 147674 222332 155994
rect 222396 148481 222424 240071
rect 222842 238096 222898 238105
rect 222842 238031 222898 238040
rect 222856 162761 222884 238031
rect 224144 229770 224172 240722
rect 224224 234660 224276 234666
rect 224224 234602 224276 234608
rect 224236 229770 224264 234602
rect 225064 232626 225092 241604
rect 225052 232620 225104 232626
rect 225052 232562 225104 232568
rect 224132 229764 224184 229770
rect 224132 229706 224184 229712
rect 224224 229764 224276 229770
rect 224224 229706 224276 229712
rect 223578 226536 223634 226545
rect 223578 226471 223634 226480
rect 223592 224233 223620 226471
rect 223578 224224 223634 224233
rect 223578 224159 223634 224168
rect 224224 221604 224276 221610
rect 224224 221546 224276 221552
rect 224236 219434 224264 221546
rect 224224 219428 224276 219434
rect 224224 219370 224276 219376
rect 222936 195288 222988 195294
rect 222936 195230 222988 195236
rect 222948 172417 222976 195230
rect 222934 172408 222990 172417
rect 222934 172343 222990 172352
rect 224236 167249 224264 219370
rect 224958 207088 225014 207097
rect 224958 207023 225014 207032
rect 224972 198014 225000 207023
rect 226524 206304 226576 206310
rect 226524 206246 226576 206252
rect 224960 198008 225012 198014
rect 224960 197950 225012 197956
rect 224960 195356 225012 195362
rect 224960 195298 225012 195304
rect 224866 173224 224922 173233
rect 224866 173159 224922 173168
rect 224880 169726 224908 173159
rect 224868 169720 224920 169726
rect 224868 169662 224920 169668
rect 224880 168434 224908 169662
rect 224316 168428 224368 168434
rect 224316 168370 224368 168376
rect 224868 168428 224920 168434
rect 224868 168370 224920 168376
rect 223578 167240 223634 167249
rect 223578 167175 223634 167184
rect 224222 167240 224278 167249
rect 224222 167175 224278 167184
rect 222842 162752 222898 162761
rect 222842 162687 222898 162696
rect 222934 156224 222990 156233
rect 222934 156159 222990 156168
rect 222382 148472 222438 148481
rect 222382 148407 222438 148416
rect 222304 147646 222792 147674
rect 222764 140978 222792 147646
rect 222948 142089 222976 156159
rect 222934 142080 222990 142089
rect 222934 142015 222990 142024
rect 223592 140978 223620 167175
rect 223672 151836 223724 151842
rect 223672 151778 223724 151784
rect 223684 147674 223712 151778
rect 223684 147646 224264 147674
rect 224132 143608 224184 143614
rect 224132 143550 224184 143556
rect 224144 140978 224172 143550
rect 224236 143426 224264 147646
rect 224328 143614 224356 168370
rect 224316 143608 224368 143614
rect 224316 143550 224368 143556
rect 224236 143398 224448 143426
rect 224420 140978 224448 143398
rect 220924 140950 221398 140978
rect 222212 140950 222502 140978
rect 222764 140950 223238 140978
rect 223592 140950 223790 140978
rect 224144 140950 224342 140978
rect 224420 140950 224894 140978
rect 218942 140828 219020 140842
rect 218942 140814 219006 140828
rect 218886 140791 218942 140800
rect 218704 140752 218756 140758
rect 218704 140694 218756 140700
rect 221832 140752 221884 140758
rect 221884 140700 222056 140706
rect 221832 140694 222056 140700
rect 221844 140678 222056 140694
rect 222028 140486 222056 140678
rect 203578 140406 204208 140434
rect 205916 140480 205968 140486
rect 206928 140480 206980 140486
rect 205968 140428 206310 140434
rect 205916 140422 206310 140428
rect 206928 140422 206980 140428
rect 218520 140480 218572 140486
rect 218520 140422 218572 140428
rect 222016 140480 222068 140486
rect 222016 140422 222068 140428
rect 205928 140406 206310 140422
rect 203522 140383 203578 140392
rect 224972 113174 225000 195298
rect 226432 185632 226484 185638
rect 226432 185574 226484 185580
rect 225144 155984 225196 155990
rect 225144 155926 225196 155932
rect 225052 151088 225104 151094
rect 225052 151030 225104 151036
rect 225064 118153 225092 151030
rect 225156 123865 225184 155926
rect 226340 143676 226392 143682
rect 226340 143618 226392 143624
rect 225326 141400 225382 141409
rect 225326 141335 225382 141344
rect 225236 140480 225288 140486
rect 225236 140422 225288 140428
rect 225248 139466 225276 140422
rect 225236 139460 225288 139466
rect 225236 139402 225288 139408
rect 225340 135561 225368 141335
rect 226352 137193 226380 143618
rect 226338 137184 226394 137193
rect 226338 137119 226394 137128
rect 225326 135552 225382 135561
rect 225326 135487 225382 135496
rect 226352 133958 226380 137119
rect 226340 133952 226392 133958
rect 226340 133894 226392 133900
rect 226340 126948 226392 126954
rect 226340 126890 226392 126896
rect 226352 126585 226380 126890
rect 226338 126576 226394 126585
rect 226338 126511 226394 126520
rect 225142 123856 225198 123865
rect 225142 123791 225198 123800
rect 226340 122800 226392 122806
rect 226340 122742 226392 122748
rect 226352 122233 226380 122742
rect 226338 122224 226394 122233
rect 226338 122159 226394 122168
rect 225050 118144 225106 118153
rect 225050 118079 225106 118088
rect 226338 117600 226394 117609
rect 226338 117535 226394 117544
rect 225142 116784 225198 116793
rect 225142 116719 225198 116728
rect 224972 113146 225092 113174
rect 225064 108390 225092 113146
rect 225052 108384 225104 108390
rect 225052 108326 225104 108332
rect 225052 108248 225104 108254
rect 225052 108190 225104 108196
rect 193416 103486 193536 103514
rect 193416 100745 193444 103486
rect 193402 100736 193458 100745
rect 193402 100671 193458 100680
rect 225064 98122 225092 108190
rect 225156 98138 225184 116719
rect 226352 116618 226380 117535
rect 226340 116612 226392 116618
rect 226340 116554 226392 116560
rect 225328 111784 225380 111790
rect 225328 111726 225380 111732
rect 225340 111353 225368 111726
rect 225326 111344 225382 111353
rect 225326 111279 225382 111288
rect 225236 108384 225288 108390
rect 225236 108326 225288 108332
rect 225248 102377 225276 108326
rect 225340 108254 225368 111279
rect 225328 108248 225380 108254
rect 225328 108190 225380 108196
rect 226338 105904 226394 105913
rect 226338 105839 226394 105848
rect 226352 105602 226380 105839
rect 226340 105596 226392 105602
rect 226340 105538 226392 105544
rect 226246 102776 226302 102785
rect 226246 102711 226302 102720
rect 225234 102368 225290 102377
rect 225234 102303 225290 102312
rect 226260 100745 226288 102711
rect 226246 100736 226302 100745
rect 226302 100694 226380 100722
rect 226246 100671 226302 100680
rect 226156 99340 226208 99346
rect 226156 99282 226208 99288
rect 225052 98116 225104 98122
rect 225156 98110 225368 98138
rect 225052 98058 225104 98064
rect 225142 98016 225198 98025
rect 224972 97974 225142 98002
rect 216126 93392 216182 93401
rect 224498 93392 224554 93401
rect 216182 93350 216628 93378
rect 224342 93350 224498 93378
rect 216126 93327 216182 93336
rect 201406 92984 201462 92993
rect 201406 92919 201462 92928
rect 193862 92848 193918 92857
rect 193324 92806 193862 92834
rect 193128 68332 193180 68338
rect 193128 68274 193180 68280
rect 193324 59362 193352 92806
rect 195518 92848 195574 92857
rect 193862 92783 193918 92792
rect 194152 88330 194180 92820
rect 194612 92806 194718 92834
rect 194796 92806 195518 92834
rect 194612 90982 194640 92806
rect 194600 90976 194652 90982
rect 194600 90918 194652 90924
rect 193864 88324 193916 88330
rect 193864 88266 193916 88272
rect 194140 88324 194192 88330
rect 194140 88266 194192 88272
rect 193876 60042 193904 88266
rect 194612 70281 194640 90918
rect 194796 84194 194824 92806
rect 200486 92848 200542 92857
rect 195518 92783 195574 92792
rect 195992 92546 196020 92820
rect 195980 92540 196032 92546
rect 195980 92482 196032 92488
rect 194704 84166 194824 84194
rect 194704 71777 194732 84166
rect 194690 71768 194746 71777
rect 194690 71703 194746 71712
rect 194704 70417 194732 71703
rect 194690 70408 194746 70417
rect 194690 70343 194746 70352
rect 195242 70408 195298 70417
rect 195242 70343 195298 70352
rect 194598 70272 194654 70281
rect 194598 70207 194654 70216
rect 194612 69873 194640 70207
rect 194598 69864 194654 69873
rect 194598 69799 194654 69808
rect 193864 60036 193916 60042
rect 193864 59978 193916 59984
rect 193312 59356 193364 59362
rect 193312 59298 193364 59304
rect 193864 59356 193916 59362
rect 193864 59298 193916 59304
rect 193876 54534 193904 59298
rect 193864 54528 193916 54534
rect 193864 54470 193916 54476
rect 193036 33788 193088 33794
rect 193036 33730 193088 33736
rect 191104 21412 191156 21418
rect 191104 21354 191156 21360
rect 195256 11762 195284 70343
rect 195334 69864 195390 69873
rect 195334 69799 195390 69808
rect 195348 64161 195376 69799
rect 195334 64152 195390 64161
rect 195334 64087 195390 64096
rect 195244 11756 195296 11762
rect 195244 11698 195296 11704
rect 180064 7676 180116 7682
rect 180064 7618 180116 7624
rect 195992 7614 196020 92482
rect 196544 92449 196572 92820
rect 196636 92806 197110 92834
rect 197662 92806 198044 92834
rect 196530 92440 196586 92449
rect 196530 92375 196586 92384
rect 196636 84194 196664 92806
rect 198016 92041 198044 92806
rect 198002 92032 198058 92041
rect 198002 91967 198058 91976
rect 196084 84182 196664 84194
rect 196072 84176 196664 84182
rect 196124 84166 196664 84176
rect 196072 84118 196124 84124
rect 198016 63510 198044 91967
rect 198384 89729 198412 92820
rect 198844 92806 198950 92834
rect 199396 92806 199502 92834
rect 200132 92806 200486 92834
rect 198370 89720 198426 89729
rect 198370 89655 198426 89664
rect 198844 79966 198872 92806
rect 199396 86902 199424 92806
rect 199384 86896 199436 86902
rect 199384 86838 199436 86844
rect 198832 79960 198884 79966
rect 198832 79902 198884 79908
rect 198844 79422 198872 79902
rect 198832 79416 198884 79422
rect 198832 79358 198884 79364
rect 198004 63504 198056 63510
rect 198004 63446 198056 63452
rect 198016 10334 198044 63446
rect 199396 28286 199424 86838
rect 200132 56574 200160 92806
rect 201420 92834 201448 92919
rect 201590 92848 201646 92857
rect 200486 92783 200542 92792
rect 200776 91905 200804 92820
rect 201342 92806 201448 92834
rect 200762 91896 200818 91905
rect 200762 91831 200818 91840
rect 201420 85474 201448 92806
rect 201512 92806 201590 92834
rect 201408 85468 201460 85474
rect 201408 85410 201460 85416
rect 201420 84862 201448 85410
rect 201408 84856 201460 84862
rect 201408 84798 201460 84804
rect 201512 64802 201540 92806
rect 207110 92848 207166 92857
rect 201646 92806 201894 92834
rect 201590 92783 201646 92792
rect 201604 92723 201632 92783
rect 202616 92478 202644 92820
rect 203182 92806 203564 92834
rect 202604 92472 202656 92478
rect 202604 92414 202656 92420
rect 203536 92313 203564 92806
rect 203628 92806 203734 92834
rect 203522 92304 203578 92313
rect 203522 92239 203578 92248
rect 203536 82754 203564 92239
rect 203628 90409 203656 92806
rect 204168 92472 204220 92478
rect 204166 92440 204168 92449
rect 204220 92440 204222 92449
rect 204166 92375 204222 92384
rect 203614 90400 203670 90409
rect 203614 90335 203670 90344
rect 203628 82754 203656 90335
rect 204456 89865 204484 92820
rect 204626 92712 204682 92721
rect 204626 92647 204682 92656
rect 204442 89856 204498 89865
rect 204442 89791 204498 89800
rect 204456 88330 204484 89791
rect 204444 88324 204496 88330
rect 204444 88266 204496 88272
rect 203524 82748 203576 82754
rect 203524 82690 203576 82696
rect 203616 82748 203668 82754
rect 203616 82690 203668 82696
rect 201500 64796 201552 64802
rect 201500 64738 201552 64744
rect 201512 63578 201540 64738
rect 201500 63572 201552 63578
rect 201500 63514 201552 63520
rect 202144 63572 202196 63578
rect 202144 63514 202196 63520
rect 200120 56568 200172 56574
rect 200120 56510 200172 56516
rect 200764 56568 200816 56574
rect 200764 56510 200816 56516
rect 200776 32434 200804 56510
rect 200764 32428 200816 32434
rect 200764 32370 200816 32376
rect 199384 28280 199436 28286
rect 199384 28222 199436 28228
rect 202156 22778 202184 63514
rect 203536 36582 203564 82690
rect 204640 60625 204668 92647
rect 205008 85513 205036 92820
rect 205100 92806 205574 92834
rect 205100 92721 205128 92806
rect 205086 92712 205142 92721
rect 205086 92647 205142 92656
rect 205100 90953 205128 92647
rect 206112 92478 206140 92820
rect 206204 92806 206862 92834
rect 206100 92472 206152 92478
rect 206100 92414 206152 92420
rect 205086 90944 205142 90953
rect 205086 90879 205142 90888
rect 204994 85504 205050 85513
rect 204994 85439 205050 85448
rect 205100 84194 205128 90879
rect 206204 84194 206232 92806
rect 208766 92848 208822 92857
rect 207166 92820 207414 92834
rect 207166 92806 207428 92820
rect 207110 92783 207166 92792
rect 207400 90273 207428 92806
rect 207386 90264 207442 90273
rect 207386 90199 207442 90208
rect 207952 89758 207980 92820
rect 208504 92806 208766 92834
rect 208306 90264 208362 90273
rect 208306 90199 208362 90208
rect 206284 89752 206336 89758
rect 206284 89694 206336 89700
rect 207940 89752 207992 89758
rect 207940 89694 207992 89700
rect 204916 84166 205128 84194
rect 205744 84166 206232 84194
rect 204626 60616 204682 60625
rect 204626 60551 204682 60560
rect 204640 60217 204668 60551
rect 204626 60208 204682 60217
rect 204626 60143 204682 60152
rect 204916 47598 204944 84166
rect 205744 73098 205772 84166
rect 206296 78606 206324 89694
rect 206284 78600 206336 78606
rect 206284 78542 206336 78548
rect 205732 73092 205784 73098
rect 205732 73034 205784 73040
rect 205744 71806 205772 73034
rect 205732 71800 205784 71806
rect 205732 71742 205784 71748
rect 204994 60208 205050 60217
rect 204994 60143 205050 60152
rect 204904 47592 204956 47598
rect 204904 47534 204956 47540
rect 203524 36576 203576 36582
rect 203524 36518 203576 36524
rect 202144 22772 202196 22778
rect 202144 22714 202196 22720
rect 205008 19990 205036 60143
rect 204996 19984 205048 19990
rect 204996 19926 205048 19932
rect 206296 13122 206324 78542
rect 208320 77314 208348 90199
rect 208400 88324 208452 88330
rect 208400 88266 208452 88272
rect 208412 86873 208440 88266
rect 208398 86864 208454 86873
rect 208398 86799 208454 86808
rect 207020 77308 207072 77314
rect 207020 77250 207072 77256
rect 208308 77308 208360 77314
rect 208308 77250 208360 77256
rect 207032 75206 207060 77250
rect 207020 75200 207072 75206
rect 207020 75142 207072 75148
rect 206376 71800 206428 71806
rect 206376 71742 206428 71748
rect 206388 38078 206416 71742
rect 208504 66230 208532 92806
rect 210054 92848 210110 92857
rect 208766 92783 208822 92792
rect 209240 89690 209268 92820
rect 209806 92806 210004 92834
rect 209228 89684 209280 89690
rect 209228 89626 209280 89632
rect 209872 88528 209924 88534
rect 209872 88470 209924 88476
rect 209884 81433 209912 88470
rect 209870 81424 209926 81433
rect 209870 81359 209926 81368
rect 209976 77217 210004 92806
rect 213642 92848 213698 92857
rect 210110 92820 210358 92834
rect 210110 92806 210372 92820
rect 210054 92783 210110 92792
rect 210344 89321 210372 92806
rect 210712 92806 211094 92834
rect 210330 89312 210386 89321
rect 210330 89247 210386 89256
rect 210712 88534 210740 92806
rect 210700 88528 210752 88534
rect 210700 88470 210752 88476
rect 211632 88330 211660 92820
rect 211816 92806 212198 92834
rect 212552 92806 212934 92834
rect 213012 92806 213642 92834
rect 211816 91050 211844 92806
rect 211804 91044 211856 91050
rect 211804 90986 211856 90992
rect 211620 88324 211672 88330
rect 211620 88266 211672 88272
rect 211066 81424 211122 81433
rect 211066 81359 211122 81368
rect 211080 79354 211108 81359
rect 211068 79348 211120 79354
rect 211068 79290 211120 79296
rect 209962 77208 210018 77217
rect 209962 77143 210018 77152
rect 209976 74534 210004 77143
rect 209976 74506 210464 74534
rect 208492 66224 208544 66230
rect 208492 66166 208544 66172
rect 209044 66224 209096 66230
rect 209044 66166 209096 66172
rect 206376 38072 206428 38078
rect 206376 38014 206428 38020
rect 206284 13116 206336 13122
rect 206284 13058 206336 13064
rect 198004 10328 198056 10334
rect 198004 10270 198056 10276
rect 209056 8974 209084 66166
rect 210436 57934 210464 74506
rect 211816 72486 211844 90986
rect 212552 81433 212580 92806
rect 213012 84194 213040 92806
rect 213642 92783 213698 92792
rect 214024 86601 214052 92820
rect 214576 89690 214604 92820
rect 214564 89684 214616 89690
rect 214564 89626 214616 89632
rect 214010 86592 214066 86601
rect 214010 86527 214066 86536
rect 215312 85542 215340 92820
rect 215864 89554 215892 92820
rect 215852 89548 215904 89554
rect 215852 89490 215904 89496
rect 215300 85536 215352 85542
rect 215300 85478 215352 85484
rect 214564 84856 214616 84862
rect 214564 84798 214616 84804
rect 212644 84166 213040 84194
rect 212538 81424 212594 81433
rect 212538 81359 212594 81368
rect 212552 80209 212580 81359
rect 212538 80200 212594 80209
rect 212538 80135 212594 80144
rect 211804 72480 211856 72486
rect 211804 72422 211856 72428
rect 212644 62082 212672 84166
rect 213182 80200 213238 80209
rect 213182 80135 213238 80144
rect 212632 62076 212684 62082
rect 212632 62018 212684 62024
rect 212644 60790 212672 62018
rect 212632 60784 212684 60790
rect 212632 60726 212684 60732
rect 210424 57928 210476 57934
rect 210424 57870 210476 57876
rect 210436 31074 210464 57870
rect 213196 57866 213224 80135
rect 213276 60784 213328 60790
rect 213276 60726 213328 60732
rect 213184 57860 213236 57866
rect 213184 57802 213236 57808
rect 213196 37942 213224 57802
rect 213184 37936 213236 37942
rect 213184 37878 213236 37884
rect 213288 35222 213316 60726
rect 213368 38072 213420 38078
rect 213368 38014 213420 38020
rect 213276 35216 213328 35222
rect 213276 35158 213328 35164
rect 210424 31068 210476 31074
rect 210424 31010 210476 31016
rect 209044 8968 209096 8974
rect 209044 8910 209096 8916
rect 195980 7608 196032 7614
rect 195980 7550 196032 7556
rect 159364 6180 159416 6186
rect 159364 6122 159416 6128
rect 213380 3466 213408 38014
rect 155224 3460 155276 3466
rect 155224 3402 155276 3408
rect 213368 3460 213420 3466
rect 213368 3402 213420 3408
rect 214576 3369 214604 84798
rect 215864 84194 215892 89490
rect 216600 84318 216628 93350
rect 224498 93327 224554 93336
rect 217152 90914 217180 92820
rect 217140 90908 217192 90914
rect 217140 90850 217192 90856
rect 217704 88097 217732 92820
rect 217690 88088 217746 88097
rect 217690 88023 217746 88032
rect 218256 86737 218284 92820
rect 218348 92806 218822 92834
rect 219558 92806 219940 92834
rect 218242 86728 218298 86737
rect 218242 86663 218298 86672
rect 216588 84312 216640 84318
rect 216588 84254 216640 84260
rect 215864 84166 215984 84194
rect 215956 66162 215984 84166
rect 216600 78674 216628 84254
rect 218348 84194 218376 92806
rect 219912 90409 219940 92806
rect 219898 90400 219954 90409
rect 219898 90335 219954 90344
rect 218072 84166 218376 84194
rect 219912 84194 219940 90335
rect 220096 89593 220124 92820
rect 220082 89584 220138 89593
rect 220082 89519 220138 89528
rect 220648 86902 220676 92820
rect 221384 90982 221412 92820
rect 221372 90976 221424 90982
rect 221372 90918 221424 90924
rect 221936 88233 221964 92820
rect 222384 91180 222436 91186
rect 222384 91122 222436 91128
rect 221922 88224 221978 88233
rect 221922 88159 221978 88168
rect 220636 86896 220688 86902
rect 220636 86838 220688 86844
rect 219912 84166 220124 84194
rect 216588 78668 216640 78674
rect 216588 78610 216640 78616
rect 218072 67590 218100 84166
rect 220096 69018 220124 84166
rect 220084 69012 220136 69018
rect 220084 68954 220136 68960
rect 218060 67584 218112 67590
rect 218060 67526 218112 67532
rect 215944 66156 215996 66162
rect 215944 66098 215996 66104
rect 215956 18630 215984 66098
rect 218072 63510 218100 67526
rect 218060 63504 218112 63510
rect 218060 63446 218112 63452
rect 222396 60722 222424 91122
rect 222488 91050 222516 92820
rect 222856 92806 223054 92834
rect 222476 91044 222528 91050
rect 222476 90986 222528 90992
rect 222856 84250 222884 92806
rect 223578 92440 223634 92449
rect 223578 92375 223634 92384
rect 223592 91798 223620 92375
rect 223580 91792 223632 91798
rect 223580 91734 223632 91740
rect 223776 91089 223804 92820
rect 224880 92546 224908 92820
rect 224868 92540 224920 92546
rect 224868 92482 224920 92488
rect 224224 91112 224276 91118
rect 223762 91080 223818 91089
rect 224224 91054 224276 91060
rect 224866 91080 224922 91089
rect 223762 91015 223818 91024
rect 222844 84244 222896 84250
rect 222844 84186 222896 84192
rect 222856 77246 222884 84186
rect 222844 77240 222896 77246
rect 222844 77182 222896 77188
rect 224236 73001 224264 91054
rect 224866 91015 224922 91024
rect 224222 72992 224278 73001
rect 224222 72927 224278 72936
rect 222384 60716 222436 60722
rect 222384 60658 222436 60664
rect 222936 60716 222988 60722
rect 222936 60658 222988 60664
rect 222844 43444 222896 43450
rect 222844 43386 222896 43392
rect 215944 18624 215996 18630
rect 215944 18566 215996 18572
rect 222856 6254 222884 43386
rect 222948 42090 222976 60658
rect 222936 42084 222988 42090
rect 222936 42026 222988 42032
rect 224880 7682 224908 91015
rect 224972 88262 225000 97974
rect 225142 97951 225198 97960
rect 225052 97912 225104 97918
rect 225052 97854 225104 97860
rect 224960 88256 225012 88262
rect 224960 88198 225012 88204
rect 225064 84153 225092 97854
rect 225340 93922 225368 98110
rect 226168 98025 226196 99282
rect 226154 98016 226210 98025
rect 226154 97951 226210 97960
rect 226248 94512 226300 94518
rect 226248 94454 226300 94460
rect 225156 93894 225368 93922
rect 225156 91118 225184 93894
rect 225144 91112 225196 91118
rect 225144 91054 225196 91060
rect 226260 90982 226288 94454
rect 226248 90976 226300 90982
rect 226248 90918 226300 90924
rect 225050 84144 225106 84153
rect 225050 84079 225106 84088
rect 226352 71738 226380 100694
rect 226444 96762 226472 185574
rect 226536 134745 226564 206246
rect 226616 180124 226668 180130
rect 226616 180066 226668 180072
rect 226522 134736 226578 134745
rect 226522 134671 226578 134680
rect 226628 129146 226656 180066
rect 226720 174554 226748 241604
rect 228376 239737 228404 241604
rect 227718 239728 227774 239737
rect 227718 239663 227774 239672
rect 228362 239728 228418 239737
rect 228362 239663 228418 239672
rect 226984 238808 227036 238814
rect 226984 238750 227036 238756
rect 226996 188358 227024 238750
rect 226984 188352 227036 188358
rect 226984 188294 227036 188300
rect 226708 174548 226760 174554
rect 226708 174490 226760 174496
rect 227076 135244 227128 135250
rect 227076 135186 227128 135192
rect 226706 134736 226762 134745
rect 226706 134671 226762 134680
rect 226720 134570 226748 134671
rect 226708 134564 226760 134570
rect 226708 134506 226760 134512
rect 226708 133884 226760 133890
rect 226708 133826 226760 133832
rect 226720 133657 226748 133826
rect 226706 133648 226762 133657
rect 226706 133583 226762 133592
rect 227088 132841 227116 135186
rect 227074 132832 227130 132841
rect 227074 132767 227130 132776
rect 226708 132456 226760 132462
rect 226708 132398 226760 132404
rect 226720 132025 226748 132398
rect 226706 132016 226762 132025
rect 226706 131951 226762 131960
rect 226708 131096 226760 131102
rect 226708 131038 226760 131044
rect 226720 130937 226748 131038
rect 226706 130928 226762 130937
rect 226706 130863 226762 130872
rect 226708 129736 226760 129742
rect 226708 129678 226760 129684
rect 226720 129305 226748 129678
rect 226706 129296 226762 129305
rect 226706 129231 226762 129240
rect 226628 129118 226748 129146
rect 226720 129062 226748 129118
rect 226708 129056 226760 129062
rect 226708 128998 226760 129004
rect 226720 128489 226748 128998
rect 226706 128480 226762 128489
rect 226706 128415 226762 128424
rect 226616 128308 226668 128314
rect 226616 128250 226668 128256
rect 226628 127401 226656 128250
rect 226614 127392 226670 127401
rect 226614 127327 226670 127336
rect 226708 126880 226760 126886
rect 226708 126822 226760 126828
rect 226720 125769 226748 126822
rect 226706 125760 226762 125769
rect 226706 125695 226762 125704
rect 226708 125520 226760 125526
rect 226708 125462 226760 125468
rect 226720 124681 226748 125462
rect 226706 124672 226762 124681
rect 226706 124607 226762 124616
rect 226708 124160 226760 124166
rect 226708 124102 226760 124108
rect 226720 123049 226748 124102
rect 226706 123040 226762 123049
rect 226706 122975 226762 122984
rect 226708 121440 226760 121446
rect 226708 121382 226760 121388
rect 226720 120329 226748 121382
rect 226706 120320 226762 120329
rect 226706 120255 226762 120264
rect 226524 119876 226576 119882
rect 226524 119818 226576 119824
rect 226536 119513 226564 119818
rect 226522 119504 226578 119513
rect 226522 119439 226578 119448
rect 226616 118652 226668 118658
rect 226616 118594 226668 118600
rect 226628 118425 226656 118594
rect 226614 118416 226670 118425
rect 226614 118351 226670 118360
rect 226708 116680 226760 116686
rect 226708 116622 226760 116628
rect 226720 115977 226748 116622
rect 226706 115968 226762 115977
rect 226706 115903 226762 115912
rect 226524 115252 226576 115258
rect 226524 115194 226576 115200
rect 226536 114889 226564 115194
rect 226522 114880 226578 114889
rect 226522 114815 226578 114824
rect 227350 114064 227406 114073
rect 227350 113999 227406 114008
rect 227364 113218 227392 113999
rect 227352 113212 227404 113218
rect 227352 113154 227404 113160
rect 226524 111104 226576 111110
rect 226524 111046 226576 111052
rect 226536 110537 226564 111046
rect 226522 110528 226578 110537
rect 226522 110463 226578 110472
rect 226984 109744 227036 109750
rect 226984 109686 227036 109692
rect 226614 108624 226670 108633
rect 226614 108559 226670 108568
rect 226628 107778 226656 108559
rect 226706 107808 226762 107817
rect 226616 107772 226668 107778
rect 226706 107743 226762 107752
rect 226616 107714 226668 107720
rect 226720 107710 226748 107743
rect 226708 107704 226760 107710
rect 226708 107646 226760 107652
rect 226706 106992 226762 107001
rect 226706 106927 226762 106936
rect 226720 106350 226748 106927
rect 226708 106344 226760 106350
rect 226708 106286 226760 106292
rect 226614 105088 226670 105097
rect 226614 105023 226670 105032
rect 226524 104848 226576 104854
rect 226524 104790 226576 104796
rect 226536 104281 226564 104790
rect 226522 104272 226578 104281
rect 226522 104207 226578 104216
rect 226628 104122 226656 105023
rect 226536 104094 226656 104122
rect 226432 96756 226484 96762
rect 226432 96698 226484 96704
rect 226432 96620 226484 96626
rect 226432 96562 226484 96568
rect 226444 96121 226472 96562
rect 226430 96112 226486 96121
rect 226430 96047 226486 96056
rect 226536 86970 226564 104094
rect 226614 103456 226670 103465
rect 226614 103391 226670 103400
rect 226628 102202 226656 103391
rect 226616 102196 226668 102202
rect 226616 102138 226668 102144
rect 226708 102128 226760 102134
rect 226708 102070 226760 102076
rect 226720 101561 226748 102070
rect 226706 101552 226762 101561
rect 226706 101487 226762 101496
rect 226616 97980 226668 97986
rect 226616 97922 226668 97928
rect 226628 97209 226656 97922
rect 226614 97200 226670 97209
rect 226614 97135 226670 97144
rect 226708 96756 226760 96762
rect 226708 96698 226760 96704
rect 226616 96552 226668 96558
rect 226616 96494 226668 96500
rect 226628 95305 226656 96494
rect 226614 95296 226670 95305
rect 226614 95231 226670 95240
rect 226720 94586 226748 96698
rect 226708 94580 226760 94586
rect 226708 94522 226760 94528
rect 226720 94489 226748 94522
rect 226706 94480 226762 94489
rect 226706 94415 226762 94424
rect 226996 93673 227024 109686
rect 227536 100020 227588 100026
rect 227536 99962 227588 99968
rect 227548 99657 227576 99962
rect 227534 99648 227590 99657
rect 227534 99583 227590 99592
rect 226982 93664 227038 93673
rect 226982 93599 227038 93608
rect 227732 91186 227760 239663
rect 227812 237448 227864 237454
rect 227812 237390 227864 237396
rect 227824 234433 227852 237390
rect 227810 234424 227866 234433
rect 227810 234359 227866 234368
rect 229940 233918 229968 241604
rect 231122 239456 231178 239465
rect 231122 239391 231178 239400
rect 229928 233912 229980 233918
rect 229928 233854 229980 233860
rect 227812 224324 227864 224330
rect 227812 224266 227864 224272
rect 227824 164257 227852 224266
rect 230388 218748 230440 218754
rect 230388 218690 230440 218696
rect 230400 218006 230428 218690
rect 229744 218000 229796 218006
rect 229744 217942 229796 217948
rect 230388 218000 230440 218006
rect 230388 217942 230440 217948
rect 227810 164248 227866 164257
rect 227810 164183 227866 164192
rect 229756 162761 229784 217942
rect 231136 211177 231164 239391
rect 231596 238814 231624 241604
rect 231584 238808 231636 238814
rect 231584 238750 231636 238756
rect 232502 213480 232558 213489
rect 232502 213415 232558 213424
rect 230478 211168 230534 211177
rect 230478 211103 230534 211112
rect 231122 211168 231178 211177
rect 231122 211103 231178 211112
rect 229190 162752 229246 162761
rect 229190 162687 229246 162696
rect 229742 162752 229798 162761
rect 229742 162687 229798 162696
rect 229204 161537 229232 162687
rect 229190 161528 229246 161537
rect 229190 161463 229246 161472
rect 227904 153332 227956 153338
rect 227904 153274 227956 153280
rect 227812 147688 227864 147694
rect 227812 147630 227864 147636
rect 227824 113257 227852 147630
rect 227916 135250 227944 153274
rect 229098 152416 229154 152425
rect 229098 152351 229154 152360
rect 228364 142248 228416 142254
rect 228364 142190 228416 142196
rect 227904 135244 227956 135250
rect 227904 135186 227956 135192
rect 228376 113830 228404 142190
rect 229112 119882 229140 152351
rect 229204 138689 229232 161463
rect 229282 150648 229338 150657
rect 229282 150583 229338 150592
rect 229190 138680 229246 138689
rect 229190 138615 229246 138624
rect 229296 133890 229324 150583
rect 229744 137080 229796 137086
rect 229744 137022 229796 137028
rect 229284 133884 229336 133890
rect 229284 133826 229336 133832
rect 229100 119876 229152 119882
rect 229100 119818 229152 119824
rect 229100 115252 229152 115258
rect 229100 115194 229152 115200
rect 228364 113824 228416 113830
rect 228364 113766 228416 113772
rect 227810 113248 227866 113257
rect 227810 113183 227866 113192
rect 227810 109712 227866 109721
rect 227810 109647 227866 109656
rect 227720 91180 227772 91186
rect 227720 91122 227772 91128
rect 226524 86964 226576 86970
rect 226524 86906 226576 86912
rect 227824 77178 227852 109647
rect 227902 102368 227958 102377
rect 227902 102303 227958 102312
rect 227812 77172 227864 77178
rect 227812 77114 227864 77120
rect 227916 73166 227944 102303
rect 227996 100020 228048 100026
rect 227996 99962 228048 99968
rect 228008 81394 228036 99962
rect 227996 81388 228048 81394
rect 227996 81330 228048 81336
rect 229112 75818 229140 115194
rect 229192 107772 229244 107778
rect 229192 107714 229244 107720
rect 229204 75857 229232 107714
rect 229756 93129 229784 137022
rect 230388 108384 230440 108390
rect 230388 108326 230440 108332
rect 230400 107778 230428 108326
rect 230388 107772 230440 107778
rect 230388 107714 230440 107720
rect 229742 93120 229798 93129
rect 229742 93055 229798 93064
rect 230492 90409 230520 211103
rect 231860 201408 231912 201414
rect 231860 201350 231912 201356
rect 230572 160200 230624 160206
rect 230572 160142 230624 160148
rect 230584 131102 230612 160142
rect 231872 159361 231900 201350
rect 231950 160168 232006 160177
rect 231950 160103 232006 160112
rect 231858 159352 231914 159361
rect 231858 159287 231914 159296
rect 231858 156088 231914 156097
rect 231858 156023 231914 156032
rect 230572 131096 230624 131102
rect 230572 131038 230624 131044
rect 231872 118658 231900 156023
rect 231964 140049 231992 160103
rect 232516 156097 232544 213415
rect 233160 201414 233188 241604
rect 234710 240136 234766 240145
rect 234710 240071 234766 240080
rect 233238 235240 233294 235249
rect 233238 235175 233294 235184
rect 233148 201408 233200 201414
rect 233148 201350 233200 201356
rect 232596 184204 232648 184210
rect 232596 184146 232648 184152
rect 232608 160177 232636 184146
rect 232594 160168 232650 160177
rect 232594 160103 232650 160112
rect 232502 156088 232558 156097
rect 232502 156023 232558 156032
rect 233252 149161 233280 235175
rect 234618 232656 234674 232665
rect 234618 232591 234620 232600
rect 234672 232591 234674 232600
rect 234620 232562 234672 232568
rect 234632 153241 234660 232562
rect 234724 229809 234752 240071
rect 234816 239494 234844 241604
rect 235998 240136 236054 240145
rect 235998 240071 236054 240080
rect 234804 239488 234856 239494
rect 234804 239430 234856 239436
rect 234710 229800 234766 229809
rect 234710 229735 234766 229744
rect 234618 153232 234674 153241
rect 234618 153167 234674 153176
rect 233238 149152 233294 149161
rect 233238 149087 233294 149096
rect 232596 142180 232648 142186
rect 232596 142122 232648 142128
rect 231950 140040 232006 140049
rect 231950 139975 232006 139984
rect 231964 135969 231992 139975
rect 231950 135960 232006 135969
rect 231950 135895 232006 135904
rect 232504 123480 232556 123486
rect 232504 123422 232556 123428
rect 231860 118652 231912 118658
rect 231860 118594 231912 118600
rect 231952 107704 232004 107710
rect 231952 107646 232004 107652
rect 230572 106344 230624 106350
rect 230572 106286 230624 106292
rect 230478 90400 230534 90409
rect 230478 90335 230534 90344
rect 229190 75848 229246 75857
rect 229100 75812 229152 75818
rect 229190 75783 229246 75792
rect 229100 75754 229152 75760
rect 230584 74458 230612 106286
rect 231860 102196 231912 102202
rect 231860 102138 231912 102144
rect 230572 74452 230624 74458
rect 230572 74394 230624 74400
rect 227904 73160 227956 73166
rect 227904 73102 227956 73108
rect 227916 71806 227944 73102
rect 227904 71800 227956 71806
rect 227904 71742 227956 71748
rect 228364 71800 228416 71806
rect 228364 71742 228416 71748
rect 226340 71732 226392 71738
rect 226340 71674 226392 71680
rect 226352 70446 226380 71674
rect 226340 70440 226392 70446
rect 226340 70382 226392 70388
rect 226984 70440 227036 70446
rect 226984 70382 227036 70388
rect 226996 43450 227024 70382
rect 226984 43444 227036 43450
rect 226984 43386 227036 43392
rect 224868 7676 224920 7682
rect 224868 7618 224920 7624
rect 222844 6248 222896 6254
rect 222844 6190 222896 6196
rect 228376 4826 228404 71742
rect 231872 70378 231900 102138
rect 231964 82657 231992 107646
rect 232516 97986 232544 123422
rect 232608 120766 232636 142122
rect 233252 121446 233280 149087
rect 234632 126886 234660 153167
rect 234620 126880 234672 126886
rect 234620 126822 234672 126828
rect 233240 121440 233292 121446
rect 233240 121382 233292 121388
rect 232596 120760 232648 120766
rect 232596 120702 232648 120708
rect 233240 119400 233292 119406
rect 233240 119342 233292 119348
rect 233148 118652 233200 118658
rect 233148 118594 233200 118600
rect 233160 117978 233188 118594
rect 233148 117972 233200 117978
rect 233148 117914 233200 117920
rect 233252 116686 233280 119342
rect 233240 116680 233292 116686
rect 233240 116622 233292 116628
rect 233148 108316 233200 108322
rect 233148 108258 233200 108264
rect 233160 107710 233188 108258
rect 233148 107704 233200 107710
rect 233148 107646 233200 107652
rect 232504 97980 232556 97986
rect 232504 97922 232556 97928
rect 231950 82648 232006 82657
rect 231950 82583 232006 82592
rect 233252 78577 233280 116622
rect 233238 78568 233294 78577
rect 233238 78503 233294 78512
rect 231860 70372 231912 70378
rect 231860 70314 231912 70320
rect 236012 66881 236040 240071
rect 236472 232558 236500 241604
rect 237392 241590 238050 241618
rect 249064 241606 249116 241612
rect 251822 241632 251878 241641
rect 236460 232552 236512 232558
rect 236460 232494 236512 232500
rect 236092 162988 236144 162994
rect 236092 162930 236144 162936
rect 236104 124166 236132 162930
rect 237392 137086 237420 241590
rect 237472 239488 237524 239494
rect 237472 239430 237524 239436
rect 237484 163538 237512 239430
rect 238850 238776 238906 238785
rect 238850 238711 238906 238720
rect 238760 229764 238812 229770
rect 238760 229706 238812 229712
rect 238772 165753 238800 229706
rect 238864 225622 238892 238711
rect 239692 228410 239720 241604
rect 240784 232552 240836 232558
rect 240784 232494 240836 232500
rect 239680 228404 239732 228410
rect 239680 228346 239732 228352
rect 238852 225616 238904 225622
rect 238852 225558 238904 225564
rect 240796 224942 240824 232494
rect 240784 224936 240836 224942
rect 240784 224878 240836 224884
rect 240796 192506 240824 224878
rect 240784 192500 240836 192506
rect 240784 192442 240836 192448
rect 238758 165744 238814 165753
rect 238758 165679 238814 165688
rect 237472 163532 237524 163538
rect 237472 163474 237524 163480
rect 238022 140992 238078 141001
rect 238022 140927 238078 140936
rect 237380 137080 237432 137086
rect 237380 137022 237432 137028
rect 236092 124160 236144 124166
rect 236092 124102 236144 124108
rect 235998 66872 236054 66881
rect 235998 66807 236054 66816
rect 228364 4820 228416 4826
rect 228364 4762 228416 4768
rect 238036 3534 238064 140927
rect 238772 132462 238800 165679
rect 239404 148368 239456 148374
rect 239404 148310 239456 148316
rect 238760 132456 238812 132462
rect 238760 132398 238812 132404
rect 238114 111888 238170 111897
rect 238114 111823 238116 111832
rect 238168 111823 238170 111832
rect 238116 111794 238168 111800
rect 239416 89622 239444 148310
rect 240690 111888 240746 111897
rect 240690 111823 240746 111832
rect 240704 111110 240732 111823
rect 240692 111104 240744 111110
rect 240692 111046 240744 111052
rect 240796 96558 240824 192442
rect 240784 96552 240836 96558
rect 240784 96494 240836 96500
rect 240784 94580 240836 94586
rect 240784 94522 240836 94528
rect 239404 89616 239456 89622
rect 239404 89558 239456 89564
rect 240796 79422 240824 94522
rect 241348 92313 241376 241604
rect 242912 240106 242940 241604
rect 244568 240106 244596 241604
rect 242164 240100 242216 240106
rect 242164 240042 242216 240048
rect 242900 240100 242952 240106
rect 242900 240042 242952 240048
rect 243544 240100 243596 240106
rect 243544 240042 243596 240048
rect 244556 240100 244608 240106
rect 244556 240042 244608 240048
rect 241518 237960 241574 237969
rect 241518 237895 241574 237904
rect 241532 111790 241560 237895
rect 242176 196654 242204 240042
rect 243556 220726 243584 240042
rect 245014 239592 245070 239601
rect 245014 239527 245070 239536
rect 244924 238808 244976 238814
rect 244924 238750 244976 238756
rect 244278 221640 244334 221649
rect 244278 221575 244334 221584
rect 244292 221474 244320 221575
rect 244280 221468 244332 221474
rect 244280 221410 244332 221416
rect 243544 220720 243596 220726
rect 243544 220662 243596 220668
rect 242900 204944 242952 204950
rect 242900 204886 242952 204892
rect 242164 196648 242216 196654
rect 242164 196590 242216 196596
rect 242164 186992 242216 186998
rect 242164 186934 242216 186940
rect 241520 111784 241572 111790
rect 241520 111726 241572 111732
rect 241334 92304 241390 92313
rect 241334 92239 241390 92248
rect 242176 91050 242204 186934
rect 242912 92546 242940 204886
rect 243544 149184 243596 149190
rect 243544 149126 243596 149132
rect 242900 92540 242952 92546
rect 242900 92482 242952 92488
rect 241612 91044 241664 91050
rect 241612 90986 241664 90992
rect 242164 91044 242216 91050
rect 242164 90986 242216 90992
rect 240140 79416 240192 79422
rect 240140 79358 240192 79364
rect 240784 79416 240836 79422
rect 240784 79358 240836 79364
rect 241520 79416 241572 79422
rect 241520 79358 241572 79364
rect 239312 4820 239364 4826
rect 239312 4762 239364 4768
rect 238024 3528 238076 3534
rect 238024 3470 238076 3476
rect 152462 3360 152518 3369
rect 152462 3295 152518 3304
rect 214562 3360 214618 3369
rect 214562 3295 214618 3304
rect 239324 480 239352 4762
rect 240152 490 240180 79358
rect 241532 16574 241560 79358
rect 241624 64870 241652 90986
rect 241612 64864 241664 64870
rect 241612 64806 241664 64812
rect 241624 63578 241652 64806
rect 241612 63572 241664 63578
rect 241612 63514 241664 63520
rect 242164 63572 242216 63578
rect 242164 63514 242216 63520
rect 241532 16546 241744 16574
rect 240336 598 240548 626
rect 240336 490 240364 598
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240152 462 240364 490
rect 240520 480 240548 598
rect 241716 480 241744 16546
rect 242176 6186 242204 63514
rect 243556 26926 243584 149126
rect 244292 108390 244320 221410
rect 244936 202842 244964 238750
rect 245028 229770 245056 239527
rect 245016 229764 245068 229770
rect 245016 229706 245068 229712
rect 245752 207052 245804 207058
rect 245752 206994 245804 207000
rect 244924 202836 244976 202842
rect 244924 202778 244976 202784
rect 244924 171828 244976 171834
rect 244924 171770 244976 171776
rect 244936 146266 244964 171770
rect 245660 162852 245712 162858
rect 245660 162794 245712 162800
rect 245672 162178 245700 162794
rect 245660 162172 245712 162178
rect 245660 162114 245712 162120
rect 244372 146260 244424 146266
rect 244372 146202 244424 146208
rect 244924 146260 244976 146266
rect 244924 146202 244976 146208
rect 244384 144974 244412 146202
rect 244372 144968 244424 144974
rect 244372 144910 244424 144916
rect 244280 108384 244332 108390
rect 244280 108326 244332 108332
rect 244384 107658 244412 144910
rect 245672 128314 245700 162114
rect 245660 128308 245712 128314
rect 245660 128250 245712 128256
rect 245672 127634 245700 128250
rect 245660 127628 245712 127634
rect 245660 127570 245712 127576
rect 244464 113212 244516 113218
rect 244464 113154 244516 113160
rect 244292 107630 244412 107658
rect 244292 104854 244320 107630
rect 244280 104848 244332 104854
rect 244280 104790 244332 104796
rect 244292 104174 244320 104790
rect 244280 104168 244332 104174
rect 244280 104110 244332 104116
rect 244476 82822 244504 113154
rect 245764 94518 245792 206994
rect 246132 171834 246160 241604
rect 247788 209778 247816 241604
rect 249076 227662 249104 241606
rect 249064 227656 249116 227662
rect 249064 227598 249116 227604
rect 247040 209772 247092 209778
rect 247040 209714 247092 209720
rect 247776 209772 247828 209778
rect 247776 209714 247828 209720
rect 246212 207664 246264 207670
rect 246212 207606 246264 207612
rect 246224 207058 246252 207606
rect 246212 207052 246264 207058
rect 246212 206994 246264 207000
rect 246304 193860 246356 193866
rect 246304 193802 246356 193808
rect 246120 171828 246172 171834
rect 246120 171770 246172 171776
rect 245752 94512 245804 94518
rect 245752 94454 245804 94460
rect 244464 82816 244516 82822
rect 244464 82758 244516 82764
rect 244476 81462 244504 82758
rect 244464 81456 244516 81462
rect 244464 81398 244516 81404
rect 244924 81456 244976 81462
rect 246316 81433 246344 193802
rect 246396 171148 246448 171154
rect 246396 171090 246448 171096
rect 246408 162858 246436 171090
rect 246396 162852 246448 162858
rect 246396 162794 246448 162800
rect 247052 100026 247080 209714
rect 249064 196648 249116 196654
rect 249064 196590 249116 196596
rect 249076 102785 249104 196590
rect 249444 171154 249472 241604
rect 250444 213240 250496 213246
rect 250444 213182 250496 213188
rect 249708 211812 249760 211818
rect 249708 211754 249760 211760
rect 249720 211177 249748 211754
rect 249706 211168 249762 211177
rect 249706 211103 249762 211112
rect 249800 211132 249852 211138
rect 249432 171148 249484 171154
rect 249432 171090 249484 171096
rect 249720 158030 249748 211103
rect 249800 211074 249852 211080
rect 249708 158024 249760 158030
rect 249708 157966 249760 157972
rect 249154 143576 249210 143585
rect 249154 143511 249210 143520
rect 249062 102776 249118 102785
rect 249062 102711 249118 102720
rect 247040 100020 247092 100026
rect 247040 99962 247092 99968
rect 249168 93158 249196 143511
rect 249156 93152 249208 93158
rect 249156 93094 249208 93100
rect 249812 92041 249840 211074
rect 249798 92032 249854 92041
rect 249798 91967 249854 91976
rect 248420 82884 248472 82890
rect 248420 82826 248472 82832
rect 244924 81398 244976 81404
rect 246302 81424 246358 81433
rect 244280 28280 244332 28286
rect 244280 28222 244332 28228
rect 243544 26920 243596 26926
rect 243544 26862 243596 26868
rect 244292 6914 244320 28222
rect 244936 15910 244964 81398
rect 246302 81359 246358 81368
rect 246304 77308 246356 77314
rect 246304 77250 246356 77256
rect 244924 15904 244976 15910
rect 244924 15846 244976 15852
rect 244292 6886 245240 6914
rect 244096 6248 244148 6254
rect 244096 6190 244148 6196
rect 242164 6180 242216 6186
rect 242164 6122 242216 6128
rect 242900 3460 242952 3466
rect 242900 3402 242952 3408
rect 242912 480 242940 3402
rect 244108 480 244136 6190
rect 245212 480 245240 6886
rect 246316 3466 246344 77250
rect 246304 3460 246356 3466
rect 246304 3402 246356 3408
rect 247592 3460 247644 3466
rect 247592 3402 247644 3408
rect 246394 3360 246450 3369
rect 246394 3295 246450 3304
rect 246408 480 246436 3295
rect 247604 480 247632 3402
rect 248432 490 248460 82826
rect 250456 77217 250484 213182
rect 251008 211138 251036 241604
rect 251822 241567 251878 241576
rect 251088 240100 251140 240106
rect 251088 240042 251140 240048
rect 251100 215286 251128 240042
rect 251178 227760 251234 227769
rect 251178 227695 251234 227704
rect 251192 216034 251220 227695
rect 251836 218006 251864 241567
rect 251914 240136 251970 240145
rect 251914 240071 251970 240080
rect 251928 228993 251956 240071
rect 251914 228984 251970 228993
rect 251914 228919 251970 228928
rect 251928 227769 251956 228919
rect 251914 227760 251970 227769
rect 251914 227695 251970 227704
rect 252468 224936 252520 224942
rect 252468 224878 252520 224884
rect 252480 224369 252508 224878
rect 252466 224360 252522 224369
rect 252466 224295 252522 224304
rect 251824 218000 251876 218006
rect 251824 217942 251876 217948
rect 251180 216028 251232 216034
rect 251180 215970 251232 215976
rect 251088 215280 251140 215286
rect 251088 215222 251140 215228
rect 251824 214600 251876 214606
rect 251824 214542 251876 214548
rect 250996 211132 251048 211138
rect 250996 211074 251048 211080
rect 251836 207670 251864 214542
rect 251824 207664 251876 207670
rect 251824 207606 251876 207612
rect 252480 178702 252508 224295
rect 252664 200122 252692 241604
rect 252756 221542 252784 264302
rect 253032 258074 253060 267706
rect 252848 258046 253060 258074
rect 252848 241466 252876 258046
rect 252926 242856 252982 242865
rect 252926 242791 252982 242800
rect 252836 241460 252888 241466
rect 252836 241402 252888 241408
rect 252744 221536 252796 221542
rect 252744 221478 252796 221484
rect 252652 200116 252704 200122
rect 252652 200058 252704 200064
rect 252664 184210 252692 200058
rect 252940 189786 252968 242791
rect 253018 242448 253074 242457
rect 253018 242383 253074 242392
rect 253032 238814 253060 242383
rect 253020 238808 253072 238814
rect 253020 238750 253072 238756
rect 253952 238066 253980 293791
rect 254044 278497 254072 312015
rect 254124 307896 254176 307902
rect 254124 307838 254176 307844
rect 254136 291145 254164 307838
rect 254122 291136 254178 291145
rect 254122 291071 254178 291080
rect 254228 287609 254256 321574
rect 255504 305108 255556 305114
rect 255504 305050 255556 305056
rect 255318 302288 255374 302297
rect 255318 302223 255374 302232
rect 255332 299418 255360 302223
rect 255410 299976 255466 299985
rect 255410 299911 255466 299920
rect 255424 299538 255452 299911
rect 255412 299532 255464 299538
rect 255412 299474 255464 299480
rect 255332 299390 255452 299418
rect 255134 299024 255190 299033
rect 255190 298982 255360 299010
rect 255134 298959 255190 298968
rect 255332 298178 255360 298982
rect 255320 298172 255372 298178
rect 255320 298114 255372 298120
rect 255320 298036 255372 298042
rect 255320 297978 255372 297984
rect 254214 287600 254270 287609
rect 254214 287535 254270 287544
rect 255332 287026 255360 297978
rect 255320 287020 255372 287026
rect 255320 286962 255372 286968
rect 255424 286906 255452 299390
rect 255516 298042 255544 305050
rect 255976 302190 256004 336738
rect 256700 335368 256752 335374
rect 256700 335310 256752 335316
rect 256054 321600 256110 321609
rect 256054 321535 256110 321544
rect 255964 302184 256016 302190
rect 255964 302126 256016 302132
rect 255688 301912 255740 301918
rect 255688 301854 255740 301860
rect 255504 298036 255556 298042
rect 255504 297978 255556 297984
rect 255502 297256 255558 297265
rect 255502 297191 255558 297200
rect 255516 296750 255544 297191
rect 255594 296848 255650 296857
rect 255594 296783 255596 296792
rect 255648 296783 255650 296792
rect 255596 296754 255648 296760
rect 255504 296744 255556 296750
rect 255504 296686 255556 296692
rect 255700 296041 255728 301854
rect 255686 296032 255742 296041
rect 255686 295967 255742 295976
rect 255502 295488 255558 295497
rect 255502 295423 255558 295432
rect 255516 295390 255544 295423
rect 255504 295384 255556 295390
rect 255504 295326 255556 295332
rect 255594 295080 255650 295089
rect 255594 295015 255650 295024
rect 255502 294672 255558 294681
rect 255502 294607 255558 294616
rect 255516 294030 255544 294607
rect 255608 294098 255636 295015
rect 255596 294092 255648 294098
rect 255596 294034 255648 294040
rect 255504 294024 255556 294030
rect 255504 293966 255556 293972
rect 255594 293312 255650 293321
rect 255504 293276 255556 293282
rect 255594 293247 255650 293256
rect 255504 293218 255556 293224
rect 255516 292913 255544 293218
rect 255502 292904 255558 292913
rect 255502 292839 255558 292848
rect 255608 292602 255636 293247
rect 255596 292596 255648 292602
rect 255596 292538 255648 292544
rect 255502 292496 255558 292505
rect 255502 292431 255558 292440
rect 255516 291242 255544 292431
rect 255700 291854 255728 295967
rect 256068 295526 256096 321535
rect 256056 295520 256108 295526
rect 256056 295462 256108 295468
rect 255962 294264 256018 294273
rect 255962 294199 256018 294208
rect 255688 291848 255740 291854
rect 255688 291790 255740 291796
rect 255594 291544 255650 291553
rect 255594 291479 255650 291488
rect 255504 291236 255556 291242
rect 255504 291178 255556 291184
rect 255504 291032 255556 291038
rect 255504 290974 255556 290980
rect 255516 290329 255544 290974
rect 255502 290320 255558 290329
rect 255502 290255 255558 290264
rect 255504 289808 255556 289814
rect 255504 289750 255556 289756
rect 255516 288969 255544 289750
rect 255608 289105 255636 291479
rect 255594 289096 255650 289105
rect 255594 289031 255650 289040
rect 255502 288960 255558 288969
rect 255502 288895 255558 288904
rect 255504 288380 255556 288386
rect 255504 288322 255556 288328
rect 255516 288153 255544 288322
rect 255502 288144 255558 288153
rect 255502 288079 255558 288088
rect 255502 287192 255558 287201
rect 255502 287127 255558 287136
rect 255516 287094 255544 287127
rect 255504 287088 255556 287094
rect 255504 287030 255556 287036
rect 255596 287020 255648 287026
rect 255596 286962 255648 286968
rect 255332 286878 255452 286906
rect 255504 286952 255556 286958
rect 255504 286894 255556 286900
rect 255332 285025 255360 286878
rect 255410 286784 255466 286793
rect 255410 286719 255466 286728
rect 255424 286346 255452 286719
rect 255412 286340 255464 286346
rect 255412 286282 255464 286288
rect 255516 285546 255544 286894
rect 255608 286385 255636 286962
rect 255594 286376 255650 286385
rect 255594 286311 255650 286320
rect 255516 285518 255636 285546
rect 255502 285424 255558 285433
rect 255502 285359 255558 285368
rect 255318 285016 255374 285025
rect 255318 284951 255374 284960
rect 255410 284608 255466 284617
rect 255410 284543 255466 284552
rect 255424 284374 255452 284543
rect 255516 284442 255544 285359
rect 255504 284436 255556 284442
rect 255504 284378 255556 284384
rect 255412 284368 255464 284374
rect 255412 284310 255464 284316
rect 255608 284209 255636 285518
rect 255594 284200 255650 284209
rect 255594 284135 255650 284144
rect 255410 283248 255466 283257
rect 255410 283183 255466 283192
rect 255424 282946 255452 283183
rect 255412 282940 255464 282946
rect 255412 282882 255464 282888
rect 255504 282872 255556 282878
rect 255504 282814 255556 282820
rect 255412 282736 255464 282742
rect 255412 282678 255464 282684
rect 255424 282441 255452 282678
rect 255410 282432 255466 282441
rect 255410 282367 255466 282376
rect 255516 282033 255544 282814
rect 255502 282024 255558 282033
rect 255502 281959 255558 281968
rect 255412 281512 255464 281518
rect 255410 281480 255412 281489
rect 255464 281480 255466 281489
rect 255410 281415 255466 281424
rect 255410 280256 255466 280265
rect 255410 280191 255412 280200
rect 255464 280191 255466 280200
rect 255412 280162 255464 280168
rect 255318 279304 255374 279313
rect 255318 279239 255374 279248
rect 255332 278798 255360 279239
rect 255320 278792 255372 278798
rect 255320 278734 255372 278740
rect 255504 278724 255556 278730
rect 255504 278666 255556 278672
rect 254030 278488 254086 278497
rect 254030 278423 254086 278432
rect 255516 278089 255544 278666
rect 255502 278080 255558 278089
rect 255502 278015 255558 278024
rect 255410 277536 255466 277545
rect 255410 277471 255412 277480
rect 255464 277471 255466 277480
rect 255412 277442 255464 277448
rect 255412 277160 255464 277166
rect 255410 277128 255412 277137
rect 255464 277128 255466 277137
rect 255410 277063 255466 277072
rect 255502 276312 255558 276321
rect 255502 276247 255558 276256
rect 255516 276078 255544 276247
rect 255504 276072 255556 276078
rect 255504 276014 255556 276020
rect 255412 276004 255464 276010
rect 255412 275946 255464 275952
rect 255424 275913 255452 275946
rect 255410 275904 255466 275913
rect 255410 275839 255466 275848
rect 255410 275360 255466 275369
rect 255410 275295 255466 275304
rect 255424 274718 255452 275295
rect 255412 274712 255464 274718
rect 255412 274654 255464 274660
rect 255504 274644 255556 274650
rect 255504 274586 255556 274592
rect 255320 274576 255372 274582
rect 255318 274544 255320 274553
rect 255372 274544 255374 274553
rect 255318 274479 255374 274488
rect 255516 274145 255544 274586
rect 255502 274136 255558 274145
rect 255502 274071 255558 274080
rect 255412 273216 255464 273222
rect 255410 273184 255412 273193
rect 255464 273184 255466 273193
rect 255410 273119 255466 273128
rect 255976 271182 256004 294199
rect 256054 285016 256110 285025
rect 256054 284951 256110 284960
rect 255964 271176 256016 271182
rect 255964 271118 256016 271124
rect 255502 270192 255558 270201
rect 255502 270127 255558 270136
rect 255410 269784 255466 269793
rect 255410 269719 255466 269728
rect 255424 269142 255452 269719
rect 255516 269210 255544 270127
rect 255504 269204 255556 269210
rect 255504 269146 255556 269152
rect 255412 269136 255464 269142
rect 255412 269078 255464 269084
rect 255318 268832 255374 268841
rect 255318 268767 255374 268776
rect 255332 267782 255360 268767
rect 255410 268424 255466 268433
rect 255410 268359 255466 268368
rect 255424 267850 255452 268359
rect 255412 267844 255464 267850
rect 255412 267786 255464 267792
rect 255320 267776 255372 267782
rect 255320 267718 255372 267724
rect 255504 267708 255556 267714
rect 255504 267650 255556 267656
rect 255516 267073 255544 267650
rect 255502 267064 255558 267073
rect 255502 266999 255558 267008
rect 255410 266656 255466 266665
rect 255410 266591 255466 266600
rect 255424 266422 255452 266591
rect 255412 266416 255464 266422
rect 255412 266358 255464 266364
rect 254032 266348 254084 266354
rect 254032 266290 254084 266296
rect 254044 266257 254072 266290
rect 254030 266248 254086 266257
rect 254030 266183 254086 266192
rect 253940 238060 253992 238066
rect 253940 238002 253992 238008
rect 254044 222902 254072 266183
rect 255318 265840 255374 265849
rect 255318 265775 255374 265784
rect 255332 265062 255360 265775
rect 255320 265056 255372 265062
rect 255320 264998 255372 265004
rect 255502 264888 255558 264897
rect 255502 264823 255558 264832
rect 255318 264480 255374 264489
rect 255318 264415 255374 264424
rect 255332 263702 255360 264415
rect 255320 263696 255372 263702
rect 255320 263638 255372 263644
rect 255516 263634 255544 264823
rect 256068 264081 256096 284951
rect 256606 283792 256662 283801
rect 256712 283778 256740 335310
rect 259644 325032 259696 325038
rect 259644 324974 259696 324980
rect 256792 322992 256844 322998
rect 256792 322934 256844 322940
rect 256804 288561 256832 322934
rect 258172 312588 258224 312594
rect 258172 312530 258224 312536
rect 258078 307864 258134 307873
rect 258078 307799 258134 307808
rect 256882 303648 256938 303657
rect 256882 303583 256938 303592
rect 256896 302938 256924 303583
rect 256884 302932 256936 302938
rect 256884 302874 256936 302880
rect 256884 302456 256936 302462
rect 256884 302398 256936 302404
rect 256790 288552 256846 288561
rect 256790 288487 256846 288496
rect 256896 287054 256924 302398
rect 256974 292768 257030 292777
rect 256974 292703 257030 292712
rect 256662 283750 256740 283778
rect 256804 287026 256924 287054
rect 256606 283727 256662 283736
rect 256606 280120 256662 280129
rect 256804 280106 256832 287026
rect 256662 280078 256832 280106
rect 256606 280055 256662 280064
rect 256988 277394 257016 292703
rect 256712 277366 257016 277394
rect 256606 271960 256662 271969
rect 256712 271946 256740 277366
rect 258092 274582 258120 307799
rect 258184 282849 258212 312530
rect 259552 311160 259604 311166
rect 259552 311102 259604 311108
rect 258262 302832 258318 302841
rect 258262 302767 258318 302776
rect 258170 282840 258226 282849
rect 258170 282775 258226 282784
rect 258276 282742 258304 302767
rect 258356 295520 258408 295526
rect 258356 295462 258408 295468
rect 258368 287094 258396 295462
rect 258356 287088 258408 287094
rect 258356 287030 258408 287036
rect 259460 287088 259512 287094
rect 259460 287030 259512 287036
rect 258264 282736 258316 282742
rect 258264 282678 258316 282684
rect 258080 274576 258132 274582
rect 258080 274518 258132 274524
rect 256662 271918 256740 271946
rect 256606 271895 256662 271904
rect 256606 271416 256662 271425
rect 256662 271374 256740 271402
rect 256606 271351 256662 271360
rect 256054 264072 256110 264081
rect 256054 264007 256110 264016
rect 255504 263628 255556 263634
rect 255504 263570 255556 263576
rect 255410 263120 255466 263129
rect 255410 263055 255412 263064
rect 255464 263055 255466 263064
rect 255412 263026 255464 263032
rect 255410 262304 255466 262313
rect 255410 262239 255412 262248
rect 255464 262239 255466 262248
rect 255412 262210 255464 262216
rect 255504 262200 255556 262206
rect 255504 262142 255556 262148
rect 255320 262132 255372 262138
rect 255320 262074 255372 262080
rect 255332 261361 255360 262074
rect 255516 261905 255544 262142
rect 255502 261896 255558 261905
rect 255502 261831 255558 261840
rect 255318 261352 255374 261361
rect 255318 261287 255374 261296
rect 255410 260944 255466 260953
rect 255410 260879 255466 260888
rect 255424 260846 255452 260879
rect 255412 260840 255464 260846
rect 255412 260782 255464 260788
rect 255410 259584 255466 259593
rect 255410 259519 255466 259528
rect 255424 259486 255452 259519
rect 255412 259480 255464 259486
rect 255412 259422 255464 259428
rect 255502 259176 255558 259185
rect 255502 259111 255558 259120
rect 255516 258126 255544 259111
rect 255504 258120 255556 258126
rect 255504 258062 255556 258068
rect 255502 257952 255558 257961
rect 255502 257887 255558 257896
rect 255320 257372 255372 257378
rect 255320 257314 255372 257320
rect 255332 257009 255360 257314
rect 255318 257000 255374 257009
rect 255318 256935 255374 256944
rect 255516 256766 255544 257887
rect 255504 256760 255556 256766
rect 255504 256702 255556 256708
rect 255412 256692 255464 256698
rect 255412 256634 255464 256640
rect 255424 256193 255452 256634
rect 255502 256592 255558 256601
rect 255502 256527 255558 256536
rect 255410 256184 255466 256193
rect 255410 256119 255466 256128
rect 255516 255338 255544 256527
rect 255504 255332 255556 255338
rect 255504 255274 255556 255280
rect 255502 255232 255558 255241
rect 255502 255167 255558 255176
rect 255516 254658 255544 255167
rect 255504 254652 255556 254658
rect 255504 254594 255556 254600
rect 255412 254584 255464 254590
rect 255412 254526 255464 254532
rect 255424 254017 255452 254526
rect 255594 254416 255650 254425
rect 255594 254351 255650 254360
rect 255410 254008 255466 254017
rect 255410 253943 255466 253952
rect 255608 253910 255636 254351
rect 255596 253904 255648 253910
rect 255596 253846 255648 253852
rect 255964 253904 256016 253910
rect 255964 253846 256016 253852
rect 255412 253224 255464 253230
rect 255412 253166 255464 253172
rect 255424 252657 255452 253166
rect 255410 252648 255466 252657
rect 255410 252583 255466 252592
rect 255594 252240 255650 252249
rect 255594 252175 255650 252184
rect 255410 251832 255466 251841
rect 255410 251767 255466 251776
rect 255424 251326 255452 251767
rect 255412 251320 255464 251326
rect 255412 251262 255464 251268
rect 255502 250880 255558 250889
rect 255502 250815 255558 250824
rect 255410 250064 255466 250073
rect 255410 249999 255466 250008
rect 255424 249830 255452 249999
rect 255516 249898 255544 250815
rect 255504 249892 255556 249898
rect 255504 249834 255556 249840
rect 255412 249824 255464 249830
rect 255412 249766 255464 249772
rect 255318 249520 255374 249529
rect 255318 249455 255374 249464
rect 255332 248470 255360 249455
rect 255410 249112 255466 249121
rect 255410 249047 255466 249056
rect 255424 248538 255452 249047
rect 255412 248532 255464 248538
rect 255412 248474 255464 248480
rect 255320 248464 255372 248470
rect 255608 248441 255636 252175
rect 255320 248406 255372 248412
rect 255594 248432 255650 248441
rect 255594 248367 255650 248376
rect 255410 248296 255466 248305
rect 255410 248231 255466 248240
rect 255318 247888 255374 247897
rect 255318 247823 255374 247832
rect 254766 245576 254822 245585
rect 254766 245511 254822 245520
rect 254122 243400 254178 243409
rect 254122 243335 254178 243344
rect 254136 240106 254164 243335
rect 254780 240106 254808 245511
rect 254124 240100 254176 240106
rect 254124 240042 254176 240048
rect 254768 240100 254820 240106
rect 254768 240042 254820 240048
rect 254582 238096 254638 238105
rect 254582 238031 254638 238040
rect 254032 222896 254084 222902
rect 254032 222838 254084 222844
rect 254596 221474 254624 238031
rect 255332 232558 255360 247823
rect 255424 247178 255452 248231
rect 255412 247172 255464 247178
rect 255412 247114 255464 247120
rect 255410 246936 255466 246945
rect 255410 246871 255466 246880
rect 255424 245750 255452 246871
rect 255686 246528 255742 246537
rect 255686 246463 255742 246472
rect 255412 245744 255464 245750
rect 255412 245686 255464 245692
rect 255502 245168 255558 245177
rect 255502 245103 255558 245112
rect 255516 244458 255544 245103
rect 255504 244452 255556 244458
rect 255504 244394 255556 244400
rect 255410 244352 255466 244361
rect 255410 244287 255412 244296
rect 255464 244287 255466 244296
rect 255412 244258 255464 244264
rect 255700 241534 255728 246463
rect 255688 241528 255740 241534
rect 255688 241470 255740 241476
rect 255976 235278 256004 253846
rect 256146 253056 256202 253065
rect 256146 252991 256202 253000
rect 256054 250472 256110 250481
rect 256054 250407 256110 250416
rect 256068 241466 256096 250407
rect 256160 247081 256188 252991
rect 256240 251932 256292 251938
rect 256240 251874 256292 251880
rect 256252 251297 256280 251874
rect 256238 251288 256294 251297
rect 256238 251223 256294 251232
rect 256422 248704 256478 248713
rect 256422 248639 256478 248648
rect 256436 247110 256464 248639
rect 256424 247104 256476 247110
rect 256146 247072 256202 247081
rect 256424 247046 256476 247052
rect 256146 247007 256202 247016
rect 256148 241528 256200 241534
rect 256148 241470 256200 241476
rect 256056 241460 256108 241466
rect 256056 241402 256108 241408
rect 256068 237969 256096 241402
rect 256054 237960 256110 237969
rect 256054 237895 256110 237904
rect 256160 236706 256188 241470
rect 256712 240786 256740 271374
rect 258078 271008 258134 271017
rect 258078 270943 258134 270952
rect 256976 251932 257028 251938
rect 256976 251874 257028 251880
rect 256884 247104 256936 247110
rect 256884 247046 256936 247052
rect 256790 246120 256846 246129
rect 256790 246055 256846 246064
rect 256700 240780 256752 240786
rect 256700 240722 256752 240728
rect 256700 240100 256752 240106
rect 256700 240042 256752 240048
rect 256148 236700 256200 236706
rect 256148 236642 256200 236648
rect 256054 235512 256110 235521
rect 256054 235447 256110 235456
rect 255964 235272 256016 235278
rect 255964 235214 256016 235220
rect 255320 232552 255372 232558
rect 255320 232494 255372 232500
rect 255964 231124 256016 231130
rect 255964 231066 256016 231072
rect 254584 221468 254636 221474
rect 254584 221410 254636 221416
rect 253940 215280 253992 215286
rect 253940 215222 253992 215228
rect 253952 203590 253980 215222
rect 255976 209710 256004 231066
rect 256068 223009 256096 235447
rect 256148 227044 256200 227050
rect 256148 226986 256200 226992
rect 256054 223000 256110 223009
rect 256054 222935 256110 222944
rect 256160 217433 256188 226986
rect 256146 217424 256202 217433
rect 256146 217359 256202 217368
rect 255964 209704 256016 209710
rect 255964 209646 256016 209652
rect 255964 207664 256016 207670
rect 255964 207606 256016 207612
rect 253940 203584 253992 203590
rect 253940 203526 253992 203532
rect 253204 202156 253256 202162
rect 253204 202098 253256 202104
rect 252928 189780 252980 189786
rect 252928 189722 252980 189728
rect 252652 184204 252704 184210
rect 252652 184146 252704 184152
rect 252468 178696 252520 178702
rect 252468 178638 252520 178644
rect 252480 178090 252508 178638
rect 251824 178084 251876 178090
rect 251824 178026 251876 178032
rect 252468 178084 252520 178090
rect 252468 178026 252520 178032
rect 251180 176724 251232 176730
rect 251180 176666 251232 176672
rect 250442 77208 250498 77217
rect 250442 77143 250498 77152
rect 250444 69692 250496 69698
rect 250444 69634 250496 69640
rect 249800 29640 249852 29646
rect 249800 29582 249852 29588
rect 249812 16574 249840 29582
rect 250456 28286 250484 69634
rect 250444 28280 250496 28286
rect 250444 28222 250496 28228
rect 249812 16546 250024 16574
rect 248616 598 248828 626
rect 248616 490 248644 598
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248432 462 248644 490
rect 248800 480 248828 598
rect 249996 480 250024 16546
rect 251192 3602 251220 176666
rect 251836 154562 251864 178026
rect 252468 177336 252520 177342
rect 252468 177278 252520 177284
rect 252480 176730 252508 177278
rect 252468 176724 252520 176730
rect 252468 176666 252520 176672
rect 252558 166288 252614 166297
rect 252558 166223 252614 166232
rect 251272 154556 251324 154562
rect 251272 154498 251324 154504
rect 251824 154556 251876 154562
rect 251824 154498 251876 154504
rect 251284 153270 251312 154498
rect 251272 153264 251324 153270
rect 251272 153206 251324 153212
rect 251284 122806 251312 153206
rect 252572 126954 252600 166223
rect 252560 126948 252612 126954
rect 252560 126890 252612 126896
rect 253020 126948 253072 126954
rect 253020 126890 253072 126896
rect 253032 126274 253060 126890
rect 253020 126268 253072 126274
rect 253020 126210 253072 126216
rect 251272 122800 251324 122806
rect 251272 122742 251324 122748
rect 252560 113824 252612 113830
rect 252560 113766 252612 113772
rect 251272 49020 251324 49026
rect 251272 48962 251324 48968
rect 251180 3596 251232 3602
rect 251180 3538 251232 3544
rect 251284 3482 251312 48962
rect 252572 16574 252600 113766
rect 253216 86902 253244 202098
rect 254584 188352 254636 188358
rect 254584 188294 254636 188300
rect 254596 91089 254624 188294
rect 255320 140820 255372 140826
rect 255320 140762 255372 140768
rect 254582 91080 254638 91089
rect 254582 91015 254638 91024
rect 253204 86896 253256 86902
rect 253204 86838 253256 86844
rect 255332 16574 255360 140762
rect 255976 123486 256004 207606
rect 256056 198008 256108 198014
rect 256056 197950 256108 197956
rect 256068 148374 256096 197950
rect 256056 148368 256108 148374
rect 256056 148310 256108 148316
rect 256712 147626 256740 240042
rect 256804 211177 256832 246055
rect 256896 233889 256924 247046
rect 256988 241670 257016 251874
rect 256976 241664 257028 241670
rect 256976 241606 257028 241612
rect 256974 238776 257030 238785
rect 256974 238711 257030 238720
rect 256882 233880 256938 233889
rect 256882 233815 256938 233824
rect 256988 232626 257016 238711
rect 256976 232620 257028 232626
rect 256976 232562 257028 232568
rect 256884 229764 256936 229770
rect 256884 229706 256936 229712
rect 256896 224262 256924 229706
rect 256884 224256 256936 224262
rect 256884 224198 256936 224204
rect 256790 211168 256846 211177
rect 256790 211103 256846 211112
rect 258092 204338 258120 270943
rect 258356 263084 258408 263090
rect 258356 263026 258408 263032
rect 258262 247344 258318 247353
rect 258262 247279 258318 247288
rect 258172 244452 258224 244458
rect 258172 244394 258224 244400
rect 258184 215966 258212 244394
rect 258276 224942 258304 247279
rect 258368 240961 258396 263026
rect 258354 240952 258410 240961
rect 258354 240887 258410 240896
rect 258724 228404 258776 228410
rect 258724 228346 258776 228352
rect 258264 224936 258316 224942
rect 258264 224878 258316 224884
rect 258172 215960 258224 215966
rect 258172 215902 258224 215908
rect 258080 204332 258132 204338
rect 258080 204274 258132 204280
rect 256700 147620 256752 147626
rect 256700 147562 256752 147568
rect 257436 147620 257488 147626
rect 257436 147562 257488 147568
rect 257448 146946 257476 147562
rect 257436 146940 257488 146946
rect 257436 146882 257488 146888
rect 257342 142216 257398 142225
rect 257342 142151 257398 142160
rect 257356 125594 257384 142151
rect 257344 125588 257396 125594
rect 257344 125530 257396 125536
rect 255964 123480 256016 123486
rect 255964 123422 256016 123428
rect 258092 89690 258120 204274
rect 258736 202881 258764 228346
rect 258722 202872 258778 202881
rect 258722 202807 258778 202816
rect 259472 164898 259500 287030
rect 259564 277166 259592 311102
rect 259656 291038 259684 324974
rect 259736 302184 259788 302190
rect 259736 302126 259788 302132
rect 259644 291032 259696 291038
rect 259644 290974 259696 290980
rect 259642 280664 259698 280673
rect 259642 280599 259698 280608
rect 259552 277160 259604 277166
rect 259552 277102 259604 277108
rect 259656 204270 259684 280599
rect 259748 277506 259776 302126
rect 259840 285025 259868 339458
rect 259826 285016 259882 285025
rect 259826 284951 259882 284960
rect 259736 277500 259788 277506
rect 259736 277442 259788 277448
rect 259748 277394 259776 277442
rect 259748 277366 259868 277394
rect 259734 269240 259790 269249
rect 259734 269175 259790 269184
rect 259748 235385 259776 269175
rect 259734 235376 259790 235385
rect 259734 235311 259790 235320
rect 259644 204264 259696 204270
rect 259644 204206 259696 204212
rect 259460 164892 259512 164898
rect 259460 164834 259512 164840
rect 259656 151814 259684 204206
rect 259840 166326 259868 277366
rect 260852 270881 260880 343606
rect 263600 340944 263652 340950
rect 263600 340886 263652 340892
rect 262220 323604 262272 323610
rect 262220 323546 262272 323552
rect 261024 320204 261076 320210
rect 261024 320146 261076 320152
rect 260932 296812 260984 296818
rect 260932 296754 260984 296760
rect 260838 270872 260894 270881
rect 260838 270807 260894 270816
rect 260840 231804 260892 231810
rect 260840 231746 260892 231752
rect 259828 166320 259880 166326
rect 259828 166262 259880 166268
rect 260104 156052 260156 156058
rect 260104 155994 260156 156000
rect 259472 151786 259684 151814
rect 259472 150521 259500 151786
rect 259458 150512 259514 150521
rect 259458 150447 259514 150456
rect 259472 125526 259500 150447
rect 259460 125520 259512 125526
rect 259460 125462 259512 125468
rect 258172 116612 258224 116618
rect 258172 116554 258224 116560
rect 258080 89684 258132 89690
rect 258080 89626 258132 89632
rect 252572 16546 253520 16574
rect 255332 16546 255912 16574
rect 252376 3596 252428 3602
rect 252376 3538 252428 3544
rect 251192 3454 251312 3482
rect 251192 480 251220 3454
rect 252388 480 252416 3538
rect 253492 480 253520 16546
rect 254676 7676 254728 7682
rect 254676 7618 254728 7624
rect 254688 480 254716 7618
rect 255884 480 255912 16546
rect 258184 3466 258212 116554
rect 259552 26920 259604 26926
rect 259552 26862 259604 26868
rect 258264 7608 258316 7614
rect 258264 7550 258316 7556
rect 257068 3460 257120 3466
rect 257068 3402 257120 3408
rect 258172 3460 258224 3466
rect 258172 3402 258224 3408
rect 257080 480 257108 3402
rect 258276 480 258304 7550
rect 259564 6914 259592 26862
rect 259472 6886 259592 6914
rect 259472 480 259500 6886
rect 260116 3466 260144 155994
rect 260852 119406 260880 231746
rect 260944 186998 260972 296754
rect 261036 287026 261064 320146
rect 261116 310548 261168 310554
rect 261116 310490 261168 310496
rect 261024 287020 261076 287026
rect 261024 286962 261076 286968
rect 261128 278905 261156 310490
rect 262232 289814 262260 323546
rect 262404 307828 262456 307834
rect 262404 307770 262456 307776
rect 262312 291236 262364 291242
rect 262312 291178 262364 291184
rect 262220 289808 262272 289814
rect 262220 289750 262272 289756
rect 262220 280220 262272 280226
rect 262220 280162 262272 280168
rect 261114 278896 261170 278905
rect 261114 278831 261170 278840
rect 261206 272232 261262 272241
rect 261206 272167 261262 272176
rect 261024 269204 261076 269210
rect 261024 269146 261076 269152
rect 261036 237153 261064 269146
rect 261114 262712 261170 262721
rect 261114 262647 261170 262656
rect 261022 237144 261078 237153
rect 261022 237079 261078 237088
rect 261128 234569 261156 262647
rect 261114 234560 261170 234569
rect 261114 234495 261170 234504
rect 261220 231810 261248 272167
rect 261208 231804 261260 231810
rect 261208 231746 261260 231752
rect 262232 213926 262260 280162
rect 262220 213920 262272 213926
rect 262220 213862 262272 213868
rect 260932 186992 260984 186998
rect 260932 186934 260984 186940
rect 260840 119400 260892 119406
rect 260840 119342 260892 119348
rect 262232 96626 262260 213862
rect 262324 177342 262352 291178
rect 262416 288386 262444 307770
rect 262494 306504 262550 306513
rect 262494 306439 262550 306448
rect 262404 288380 262456 288386
rect 262404 288322 262456 288328
rect 262402 285696 262458 285705
rect 262402 285631 262458 285640
rect 262416 211206 262444 285631
rect 262508 282878 262536 306439
rect 262496 282872 262548 282878
rect 262496 282814 262548 282820
rect 263612 262138 263640 340886
rect 264256 321570 264284 703326
rect 267660 699825 267688 703520
rect 282184 703316 282236 703322
rect 282184 703258 282236 703264
rect 273904 703248 273956 703254
rect 273904 703190 273956 703196
rect 267646 699816 267702 699825
rect 267646 699751 267702 699760
rect 269764 364404 269816 364410
rect 269764 364346 269816 364352
rect 267832 342304 267884 342310
rect 267832 342246 267884 342252
rect 266452 332716 266504 332722
rect 266452 332658 266504 332664
rect 266360 331288 266412 331294
rect 266360 331230 266412 331236
rect 264244 321564 264296 321570
rect 264244 321506 264296 321512
rect 264256 321094 264284 321506
rect 263784 321088 263836 321094
rect 263784 321030 263836 321036
rect 264244 321088 264296 321094
rect 264244 321030 264296 321036
rect 263690 313304 263746 313313
rect 263690 313239 263746 313248
rect 263704 273222 263732 313239
rect 263692 273216 263744 273222
rect 263692 273158 263744 273164
rect 263796 266354 263824 321030
rect 265072 313404 265124 313410
rect 265072 313346 265124 313352
rect 263876 311908 263928 311914
rect 263876 311850 263928 311856
rect 263888 278730 263916 311850
rect 264978 291816 265034 291825
rect 264978 291751 265034 291760
rect 263876 278724 263928 278730
rect 263876 278666 263928 278672
rect 264058 273456 264114 273465
rect 264058 273391 264114 273400
rect 263966 268152 264022 268161
rect 263966 268087 264022 268096
rect 263784 266348 263836 266354
rect 263784 266290 263836 266296
rect 263690 265432 263746 265441
rect 263690 265367 263746 265376
rect 263704 265062 263732 265367
rect 263692 265056 263744 265062
rect 263692 264998 263744 265004
rect 263600 262132 263652 262138
rect 263600 262074 263652 262080
rect 263704 258074 263732 264998
rect 263704 258046 263824 258074
rect 262496 250572 262548 250578
rect 262496 250514 262548 250520
rect 262508 249898 262536 250514
rect 262496 249892 262548 249898
rect 262496 249834 262548 249840
rect 262508 230489 262536 249834
rect 262494 230480 262550 230489
rect 262494 230415 262550 230424
rect 262404 211200 262456 211206
rect 262404 211142 262456 211148
rect 262312 177336 262364 177342
rect 262312 177278 262364 177284
rect 262416 109750 262444 211142
rect 263600 211132 263652 211138
rect 263600 211074 263652 211080
rect 262404 109744 262456 109750
rect 262404 109686 262456 109692
rect 262220 96620 262272 96626
rect 262220 96562 262272 96568
rect 262864 93152 262916 93158
rect 262864 93094 262916 93100
rect 262218 58576 262274 58585
rect 262218 58511 262274 58520
rect 262232 16574 262260 58511
rect 262232 16546 262536 16574
rect 261760 15904 261812 15910
rect 261760 15846 261812 15852
rect 260656 3528 260708 3534
rect 260656 3470 260708 3476
rect 260104 3460 260156 3466
rect 260104 3402 260156 3408
rect 260668 480 260696 3470
rect 261772 480 261800 15846
rect 262508 490 262536 16546
rect 262876 3330 262904 93094
rect 263612 88330 263640 211074
rect 263796 207641 263824 258046
rect 263876 251864 263928 251870
rect 263876 251806 263928 251812
rect 263888 251326 263916 251806
rect 263876 251320 263928 251326
rect 263876 251262 263928 251268
rect 263888 226302 263916 251262
rect 263980 231849 264008 268087
rect 263966 231840 264022 231849
rect 263966 231775 264022 231784
rect 263876 226296 263928 226302
rect 263876 226238 263928 226244
rect 264072 211138 264100 273391
rect 264888 224460 264940 224466
rect 264888 224402 264940 224408
rect 264060 211132 264112 211138
rect 264060 211074 264112 211080
rect 263782 207632 263838 207641
rect 263782 207567 263838 207576
rect 264900 140146 264928 224402
rect 264992 169046 265020 291751
rect 265084 281518 265112 313346
rect 265162 304192 265218 304201
rect 265162 304127 265218 304136
rect 265072 281512 265124 281518
rect 265072 281454 265124 281460
rect 265176 273057 265204 304127
rect 266372 298081 266400 331230
rect 266358 298072 266414 298081
rect 266358 298007 266414 298016
rect 266360 284436 266412 284442
rect 266360 284378 266412 284384
rect 265162 273048 265218 273057
rect 265162 272983 265218 272992
rect 265164 266416 265216 266422
rect 265164 266358 265216 266364
rect 265072 262268 265124 262274
rect 265072 262210 265124 262216
rect 265084 219337 265112 262210
rect 265176 227730 265204 266358
rect 265256 250504 265308 250510
rect 265256 250446 265308 250452
rect 265268 249830 265296 250446
rect 265256 249824 265308 249830
rect 265256 249766 265308 249772
rect 265164 227724 265216 227730
rect 265164 227666 265216 227672
rect 265268 219434 265296 249766
rect 266372 223582 266400 284378
rect 266464 277001 266492 332658
rect 266634 316160 266690 316169
rect 266634 316095 266690 316104
rect 267740 316124 267792 316130
rect 266544 278792 266596 278798
rect 266544 278734 266596 278740
rect 266450 276992 266506 277001
rect 266450 276927 266506 276936
rect 266452 271176 266504 271182
rect 266452 271118 266504 271124
rect 266360 223576 266412 223582
rect 266360 223518 266412 223524
rect 265256 219428 265308 219434
rect 265256 219370 265308 219376
rect 265070 219328 265126 219337
rect 265070 219263 265126 219272
rect 264980 169040 265032 169046
rect 264980 168982 265032 168988
rect 264888 140140 264940 140146
rect 264888 140082 264940 140088
rect 264900 139466 264928 140082
rect 264888 139460 264940 139466
rect 264888 139402 264940 139408
rect 266372 102134 266400 223518
rect 266464 158817 266492 271118
rect 266556 214606 266584 278734
rect 266648 256698 266676 316095
rect 267740 316066 267792 316072
rect 266910 298072 266966 298081
rect 266910 298007 266966 298016
rect 266924 297401 266952 298007
rect 266910 297392 266966 297401
rect 266910 297327 266966 297336
rect 267752 286346 267780 316066
rect 267740 286340 267792 286346
rect 267740 286282 267792 286288
rect 266636 256692 266688 256698
rect 266636 256634 266688 256640
rect 266728 255264 266780 255270
rect 266728 255206 266780 255212
rect 266740 254658 266768 255206
rect 266728 254652 266780 254658
rect 266728 254594 266780 254600
rect 266740 254017 266768 254594
rect 266726 254008 266782 254017
rect 266726 253943 266782 253952
rect 266636 248464 266688 248470
rect 266636 248406 266688 248412
rect 266648 217326 266676 248406
rect 266636 217320 266688 217326
rect 266636 217262 266688 217268
rect 266544 214600 266596 214606
rect 266544 214542 266596 214548
rect 266450 158808 266506 158817
rect 266450 158743 266506 158752
rect 266464 129742 266492 158743
rect 267752 135250 267780 286282
rect 267844 276010 267872 342246
rect 269212 305652 269264 305658
rect 269212 305594 269264 305600
rect 267924 294092 267976 294098
rect 267924 294034 267976 294040
rect 267832 276004 267884 276010
rect 267832 275946 267884 275952
rect 267832 267844 267884 267850
rect 267832 267786 267884 267792
rect 267844 234598 267872 267786
rect 267832 234592 267884 234598
rect 267832 234534 267884 234540
rect 267844 145586 267872 234534
rect 267936 224466 267964 294034
rect 269120 291848 269172 291854
rect 269120 291790 269172 291796
rect 268016 269136 268068 269142
rect 268016 269078 268068 269084
rect 268028 238513 268056 269078
rect 268108 258052 268160 258058
rect 268108 257994 268160 258000
rect 268120 257378 268148 257994
rect 268108 257372 268160 257378
rect 268108 257314 268160 257320
rect 268120 257281 268148 257314
rect 268106 257272 268162 257281
rect 268106 257207 268162 257216
rect 268014 238504 268070 238513
rect 268014 238439 268070 238448
rect 267924 224460 267976 224466
rect 267924 224402 267976 224408
rect 268382 148336 268438 148345
rect 268382 148271 268438 148280
rect 267832 145580 267884 145586
rect 267832 145522 267884 145528
rect 267740 135244 267792 135250
rect 267740 135186 267792 135192
rect 266452 129736 266504 129742
rect 266452 129678 266504 129684
rect 267832 129736 267884 129742
rect 267832 129678 267884 129684
rect 266360 102128 266412 102134
rect 266360 102070 266412 102076
rect 264244 95940 264296 95946
rect 264244 95882 264296 95888
rect 263600 88324 263652 88330
rect 263600 88266 263652 88272
rect 264256 74497 264284 95882
rect 266360 84312 266412 84318
rect 266360 84254 266412 84260
rect 264242 74488 264298 74497
rect 264242 74423 264298 74432
rect 264256 73273 264284 74423
rect 263598 73264 263654 73273
rect 263598 73199 263654 73208
rect 264242 73264 264298 73273
rect 264242 73199 264298 73208
rect 263612 16574 263640 73199
rect 264980 60036 265032 60042
rect 264980 59978 265032 59984
rect 263612 16546 264192 16574
rect 262864 3324 262916 3330
rect 262864 3266 262916 3272
rect 262784 598 262996 626
rect 262784 490 262812 598
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262508 462 262812 490
rect 262968 480 262996 598
rect 264164 480 264192 16546
rect 264992 490 265020 59978
rect 266372 16574 266400 84254
rect 266372 16546 266584 16574
rect 265176 598 265388 626
rect 265176 490 265204 598
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 264992 462 265204 490
rect 265360 480 265388 598
rect 266556 480 266584 16546
rect 267844 6914 267872 129678
rect 268396 16574 268424 148271
rect 269132 133890 269160 291790
rect 269224 274650 269252 305594
rect 269304 284368 269356 284374
rect 269304 284310 269356 284316
rect 269212 274644 269264 274650
rect 269212 274586 269264 274592
rect 269210 244352 269266 244361
rect 269210 244287 269266 244296
rect 269224 215937 269252 244287
rect 269210 215928 269266 215937
rect 269210 215863 269266 215872
rect 269120 133884 269172 133890
rect 269120 133826 269172 133832
rect 269224 89729 269252 215863
rect 269316 200054 269344 284310
rect 269776 253230 269804 364346
rect 270592 325712 270644 325718
rect 270592 325654 270644 325660
rect 270500 300892 270552 300898
rect 270500 300834 270552 300840
rect 269396 253224 269448 253230
rect 269396 253166 269448 253172
rect 269764 253224 269816 253230
rect 269764 253166 269816 253172
rect 269408 228410 269436 253166
rect 269396 228404 269448 228410
rect 269396 228346 269448 228352
rect 269304 200048 269356 200054
rect 269304 199990 269356 199996
rect 270512 105602 270540 300834
rect 270604 293282 270632 325654
rect 273916 315518 273944 703190
rect 280804 703180 280856 703186
rect 280804 703122 280856 703128
rect 277308 700324 277360 700330
rect 277308 700266 277360 700272
rect 273352 315512 273404 315518
rect 273352 315454 273404 315460
rect 273904 315512 273956 315518
rect 273904 315454 273956 315460
rect 273364 315314 273392 315454
rect 273352 315308 273404 315314
rect 273352 315250 273404 315256
rect 273260 294024 273312 294030
rect 273260 293966 273312 293972
rect 270592 293276 270644 293282
rect 270592 293218 270644 293224
rect 270604 188358 270632 293218
rect 270684 282940 270736 282946
rect 270684 282882 270736 282888
rect 270696 206990 270724 282882
rect 271878 272504 271934 272513
rect 271878 272439 271934 272448
rect 270776 256760 270828 256766
rect 270776 256702 270828 256708
rect 270788 227730 270816 256702
rect 270776 227724 270828 227730
rect 270776 227666 270828 227672
rect 270788 227050 270816 227666
rect 270776 227044 270828 227050
rect 270776 226986 270828 226992
rect 270684 206984 270736 206990
rect 270684 206926 270736 206932
rect 270696 202162 270724 206926
rect 270684 202156 270736 202162
rect 270684 202098 270736 202104
rect 270592 188352 270644 188358
rect 270592 188294 270644 188300
rect 271892 150385 271920 272439
rect 271972 263696 272024 263702
rect 271972 263638 272024 263644
rect 271984 195294 272012 263638
rect 272064 255332 272116 255338
rect 272064 255274 272116 255280
rect 272076 231810 272104 255274
rect 272156 247172 272208 247178
rect 272156 247114 272208 247120
rect 272064 231804 272116 231810
rect 272064 231746 272116 231752
rect 272168 229770 272196 247114
rect 272340 231804 272392 231810
rect 272340 231746 272392 231752
rect 272352 231130 272380 231746
rect 272340 231124 272392 231130
rect 272340 231066 272392 231072
rect 272156 229764 272208 229770
rect 272156 229706 272208 229712
rect 271972 195288 272024 195294
rect 271972 195230 272024 195236
rect 273272 170474 273300 293966
rect 273364 263702 273392 315250
rect 276018 304056 276074 304065
rect 276018 303991 276074 304000
rect 274732 302932 274784 302938
rect 274732 302874 274784 302880
rect 273444 276072 273496 276078
rect 273444 276014 273496 276020
rect 273352 263696 273404 263702
rect 273352 263638 273404 263644
rect 273352 256012 273404 256018
rect 273352 255954 273404 255960
rect 273364 250578 273392 255954
rect 273352 250572 273404 250578
rect 273352 250514 273404 250520
rect 273456 220794 273484 276014
rect 274640 274644 274692 274650
rect 274640 274586 274692 274592
rect 273536 267776 273588 267782
rect 273536 267718 273588 267724
rect 273548 229090 273576 267718
rect 273628 255196 273680 255202
rect 273628 255138 273680 255144
rect 273640 254590 273668 255138
rect 273628 254584 273680 254590
rect 273628 254526 273680 254532
rect 273640 254017 273668 254526
rect 273626 254008 273682 254017
rect 273626 253943 273682 253952
rect 273536 229084 273588 229090
rect 273536 229026 273588 229032
rect 273444 220788 273496 220794
rect 273444 220730 273496 220736
rect 273548 219434 273576 229026
rect 273364 219406 273576 219434
rect 273260 170468 273312 170474
rect 273260 170410 273312 170416
rect 271878 150376 271934 150385
rect 271878 150311 271934 150320
rect 273364 115258 273392 219406
rect 274652 159390 274680 274586
rect 274744 213246 274772 302874
rect 275282 253192 275338 253201
rect 275282 253127 275338 253136
rect 275296 241505 275324 253127
rect 275282 241496 275338 241505
rect 275282 241431 275338 241440
rect 274732 213240 274784 213246
rect 274732 213182 274784 213188
rect 276032 198014 276060 303991
rect 276110 276720 276166 276729
rect 276110 276655 276166 276664
rect 276020 198008 276072 198014
rect 276020 197950 276072 197956
rect 274640 159384 274692 159390
rect 274640 159326 274692 159332
rect 276020 140140 276072 140146
rect 276020 140082 276072 140088
rect 273904 133884 273956 133890
rect 273904 133826 273956 133832
rect 273352 115252 273404 115258
rect 273352 115194 273404 115200
rect 270500 105596 270552 105602
rect 270500 105538 270552 105544
rect 270512 105194 270540 105538
rect 270500 105188 270552 105194
rect 270500 105130 270552 105136
rect 271144 105188 271196 105194
rect 271144 105130 271196 105136
rect 269764 102196 269816 102202
rect 269764 102138 269816 102144
rect 269210 89720 269266 89729
rect 269210 89655 269266 89664
rect 269120 50380 269172 50386
rect 269120 50322 269172 50328
rect 268396 16546 268516 16574
rect 267844 6886 268424 6914
rect 267740 3324 267792 3330
rect 267740 3266 267792 3272
rect 267752 480 267780 3266
rect 268396 490 268424 6886
rect 268488 3330 268516 16546
rect 269132 6914 269160 50322
rect 269776 7614 269804 102138
rect 270500 33788 270552 33794
rect 270500 33730 270552 33736
rect 270512 16574 270540 33730
rect 270512 16546 270816 16574
rect 269764 7608 269816 7614
rect 269764 7550 269816 7556
rect 269132 6886 270080 6914
rect 268476 3324 268528 3330
rect 268476 3266 268528 3272
rect 268672 598 268884 626
rect 268672 490 268700 598
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268396 462 268700 490
rect 268856 480 268884 598
rect 270052 480 270080 6886
rect 270788 490 270816 16546
rect 271156 16250 271184 105130
rect 271144 16244 271196 16250
rect 271144 16186 271196 16192
rect 273916 3466 273944 133826
rect 274824 13116 274876 13122
rect 274824 13058 274876 13064
rect 272432 3460 272484 3466
rect 272432 3402 272484 3408
rect 273904 3460 273956 3466
rect 273904 3402 273956 3408
rect 271064 598 271276 626
rect 271064 490 271092 598
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 270788 462 271092 490
rect 271248 480 271276 598
rect 272444 480 272472 3402
rect 273628 3324 273680 3330
rect 273628 3266 273680 3272
rect 273640 480 273668 3266
rect 274836 480 274864 13058
rect 276032 3602 276060 140082
rect 276124 131102 276152 276655
rect 277320 267714 277348 700266
rect 278044 311908 278096 311914
rect 278044 311850 278096 311856
rect 277398 301064 277454 301073
rect 277398 300999 277454 301008
rect 277308 267708 277360 267714
rect 277308 267650 277360 267656
rect 277320 266422 277348 267650
rect 277308 266416 277360 266422
rect 277308 266358 277360 266364
rect 276202 262984 276258 262993
rect 276202 262919 276258 262928
rect 276216 230450 276244 262919
rect 276204 230444 276256 230450
rect 276204 230386 276256 230392
rect 276216 207670 276244 230386
rect 276204 207664 276256 207670
rect 276204 207606 276256 207612
rect 276112 131096 276164 131102
rect 276112 131038 276164 131044
rect 277412 63510 277440 300999
rect 277492 266416 277544 266422
rect 277492 266358 277544 266364
rect 277504 201482 277532 266358
rect 277584 258120 277636 258126
rect 277584 258062 277636 258068
rect 277596 227633 277624 258062
rect 278056 251938 278084 311850
rect 280250 299568 280306 299577
rect 280250 299503 280306 299512
rect 278778 294536 278834 294545
rect 278778 294471 278834 294480
rect 278688 258732 278740 258738
rect 278688 258674 278740 258680
rect 278700 258126 278728 258674
rect 278688 258120 278740 258126
rect 278688 258062 278740 258068
rect 278044 251932 278096 251938
rect 278044 251874 278096 251880
rect 278044 248532 278096 248538
rect 278044 248474 278096 248480
rect 278056 233306 278084 248474
rect 278044 233300 278096 233306
rect 278044 233242 278096 233248
rect 277582 227624 277638 227633
rect 277582 227559 277638 227568
rect 277492 201476 277544 201482
rect 277492 201418 277544 201424
rect 278056 191826 278084 233242
rect 278044 191820 278096 191826
rect 278044 191762 278096 191768
rect 278792 139398 278820 294471
rect 280160 292596 280212 292602
rect 280160 292538 280212 292544
rect 278872 263628 278924 263634
rect 278872 263570 278924 263576
rect 278884 209681 278912 263570
rect 278870 209672 278926 209681
rect 278870 209607 278926 209616
rect 278780 139392 278832 139398
rect 278780 139334 278832 139340
rect 280068 139392 280120 139398
rect 280068 139334 280120 139340
rect 280080 138718 280108 139334
rect 280068 138712 280120 138718
rect 280068 138654 280120 138660
rect 278044 134564 278096 134570
rect 278044 134506 278096 134512
rect 277400 63504 277452 63510
rect 277400 63446 277452 63452
rect 277400 43444 277452 43450
rect 277400 43386 277452 43392
rect 276112 16244 276164 16250
rect 276112 16186 276164 16192
rect 276020 3596 276072 3602
rect 276020 3538 276072 3544
rect 276124 3482 276152 16186
rect 277412 6914 277440 43386
rect 278056 9042 278084 134506
rect 280172 95946 280200 292538
rect 280264 125594 280292 299503
rect 280816 262993 280844 703122
rect 281538 298752 281594 298761
rect 281538 298687 281594 298696
rect 280802 262984 280858 262993
rect 280802 262919 280858 262928
rect 281552 193866 281580 298687
rect 281632 274712 281684 274718
rect 281632 274654 281684 274660
rect 281644 204950 281672 274654
rect 282196 263634 282224 703258
rect 283852 700330 283880 703520
rect 300136 703118 300164 703520
rect 332520 703390 332548 703520
rect 332508 703384 332560 703390
rect 332508 703326 332560 703332
rect 300124 703112 300176 703118
rect 300124 703054 300176 703060
rect 287704 703044 287756 703050
rect 287704 702986 287756 702992
rect 286324 702976 286376 702982
rect 286324 702918 286376 702924
rect 283840 700324 283892 700330
rect 283840 700266 283892 700272
rect 286336 310457 286364 702918
rect 285678 310448 285734 310457
rect 285678 310383 285734 310392
rect 286322 310448 286378 310457
rect 286322 310383 286378 310392
rect 285692 309369 285720 310383
rect 285678 309360 285734 309369
rect 285678 309295 285734 309304
rect 282920 296744 282972 296750
rect 282920 296686 282972 296692
rect 282184 263628 282236 263634
rect 282184 263570 282236 263576
rect 281632 204944 281684 204950
rect 281632 204886 281684 204892
rect 281540 193860 281592 193866
rect 281540 193802 281592 193808
rect 282932 145625 282960 296686
rect 284392 295384 284444 295390
rect 284392 295326 284444 295332
rect 284298 241768 284354 241777
rect 284298 241703 284354 241712
rect 282918 145616 282974 145625
rect 282918 145551 282920 145560
rect 282972 145551 282974 145560
rect 282920 145522 282972 145528
rect 280252 125588 280304 125594
rect 280252 125530 280304 125536
rect 281448 125588 281500 125594
rect 281448 125530 281500 125536
rect 281460 124914 281488 125530
rect 281448 124908 281500 124914
rect 281448 124850 281500 124856
rect 280160 95940 280212 95946
rect 280160 95882 280212 95888
rect 284312 82754 284340 241703
rect 284404 196654 284432 295326
rect 285692 262206 285720 309295
rect 287060 299532 287112 299538
rect 287060 299474 287112 299480
rect 285680 262200 285732 262206
rect 285680 262142 285732 262148
rect 285772 244316 285824 244322
rect 285772 244258 285824 244264
rect 284392 196648 284444 196654
rect 284392 196590 284444 196596
rect 285680 167068 285732 167074
rect 285680 167010 285732 167016
rect 284944 104168 284996 104174
rect 284944 104110 284996 104116
rect 284300 82748 284352 82754
rect 284300 82690 284352 82696
rect 284312 82142 284340 82690
rect 284300 82136 284352 82142
rect 284300 82078 284352 82084
rect 280804 80708 280856 80714
rect 280804 80650 280856 80656
rect 280158 73808 280214 73817
rect 280158 73743 280214 73752
rect 278688 63504 278740 63510
rect 278688 63446 278740 63452
rect 278700 62830 278728 63446
rect 278688 62824 278740 62830
rect 278688 62766 278740 62772
rect 280172 16574 280200 73743
rect 280172 16546 280752 16574
rect 278044 9036 278096 9042
rect 278044 8978 278096 8984
rect 279516 8968 279568 8974
rect 279516 8910 279568 8916
rect 277412 6886 278360 6914
rect 277124 3596 277176 3602
rect 277124 3538 277176 3544
rect 276032 3454 276152 3482
rect 276032 480 276060 3454
rect 277136 480 277164 3538
rect 278332 480 278360 6886
rect 279528 480 279556 8910
rect 280724 480 280752 16546
rect 280816 3330 280844 80650
rect 281540 71052 281592 71058
rect 281540 70994 281592 71000
rect 280804 3324 280856 3330
rect 280804 3266 280856 3272
rect 281552 490 281580 70994
rect 284392 18624 284444 18630
rect 284392 18566 284444 18572
rect 284404 6914 284432 18566
rect 284956 13122 284984 104110
rect 285692 16574 285720 167010
rect 285784 86970 285812 244258
rect 287072 99346 287100 299474
rect 287716 260846 287744 702986
rect 348804 702545 348832 703520
rect 364996 702914 365024 703520
rect 397472 703322 397500 703520
rect 397460 703316 397512 703322
rect 397460 703258 397512 703264
rect 413664 703254 413692 703520
rect 413652 703248 413704 703254
rect 413652 703190 413704 703196
rect 364984 702908 365036 702914
rect 364984 702850 365036 702856
rect 429856 702778 429884 703520
rect 462332 703186 462360 703520
rect 462320 703180 462372 703186
rect 462320 703122 462372 703128
rect 478524 702846 478552 703520
rect 478512 702840 478564 702846
rect 478512 702782 478564 702788
rect 429844 702772 429896 702778
rect 429844 702714 429896 702720
rect 494808 702710 494836 703520
rect 494796 702704 494848 702710
rect 494796 702646 494848 702652
rect 527192 702642 527220 703520
rect 543476 702982 543504 703520
rect 543464 702976 543516 702982
rect 543464 702918 543516 702924
rect 527180 702636 527232 702642
rect 527180 702578 527232 702584
rect 348790 702536 348846 702545
rect 559668 702506 559696 703520
rect 580172 703044 580224 703050
rect 580172 702986 580224 702992
rect 348790 702471 348846 702480
rect 559656 702500 559708 702506
rect 559656 702442 559708 702448
rect 580184 697241 580212 702986
rect 582380 702568 582432 702574
rect 582380 702510 582432 702516
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 582392 670721 582420 702510
rect 582746 683904 582802 683913
rect 582746 683839 582802 683848
rect 582378 670712 582434 670721
rect 582378 670647 582434 670656
rect 582378 644056 582434 644065
rect 582378 643991 582434 644000
rect 580170 511320 580226 511329
rect 580170 511255 580172 511264
rect 580224 511255 580226 511264
rect 580172 511226 580224 511232
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 580184 364410 580212 365055
rect 580172 364404 580224 364410
rect 580172 364346 580224 364352
rect 574744 351960 574796 351966
rect 580172 351960 580224 351966
rect 574744 351902 574796 351908
rect 580170 351928 580172 351937
rect 580224 351928 580226 351937
rect 288440 298172 288492 298178
rect 288440 298114 288492 298120
rect 287704 260840 287756 260846
rect 287704 260782 287756 260788
rect 287152 245744 287204 245750
rect 287152 245686 287204 245692
rect 287164 124166 287192 245686
rect 288452 155922 288480 298114
rect 309782 297392 309838 297401
rect 309782 297327 309838 297336
rect 289728 260160 289780 260166
rect 289728 260102 289780 260108
rect 289740 259486 289768 260102
rect 288532 259480 288584 259486
rect 288532 259422 288584 259428
rect 289728 259480 289780 259486
rect 289728 259422 289780 259428
rect 288544 212537 288572 259422
rect 288530 212528 288586 212537
rect 288530 212463 288586 212472
rect 288440 155916 288492 155922
rect 288440 155858 288492 155864
rect 287704 140072 287756 140078
rect 287704 140014 287756 140020
rect 287152 124160 287204 124166
rect 287152 124102 287204 124108
rect 287060 99340 287112 99346
rect 287060 99282 287112 99288
rect 285772 86964 285824 86970
rect 285772 86906 285824 86912
rect 285784 86873 285812 86906
rect 285770 86864 285826 86873
rect 285770 86799 285826 86808
rect 287060 35216 287112 35222
rect 287060 35158 287112 35164
rect 287072 16574 287100 35158
rect 285692 16546 286640 16574
rect 287072 16546 287376 16574
rect 284944 13116 284996 13122
rect 284944 13058 284996 13064
rect 284404 6886 284984 6914
rect 283104 3460 283156 3466
rect 283104 3402 283156 3408
rect 281736 598 281948 626
rect 281736 490 281764 598
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281552 462 281764 490
rect 281920 480 281948 598
rect 283116 480 283144 3402
rect 284300 3324 284352 3330
rect 284300 3266 284352 3272
rect 284312 480 284340 3266
rect 284956 490 284984 6886
rect 285232 598 285444 626
rect 285232 490 285260 598
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 284956 462 285260 490
rect 285416 480 285444 598
rect 286612 480 286640 16546
rect 287348 490 287376 16546
rect 287716 3534 287744 140014
rect 288544 108322 288572 212463
rect 295984 175364 296036 175370
rect 295984 175306 296036 175312
rect 289728 155916 289780 155922
rect 289728 155858 289780 155864
rect 289740 155242 289768 155858
rect 289728 155236 289780 155242
rect 289728 155178 289780 155184
rect 289084 140888 289136 140894
rect 289084 140830 289136 140836
rect 288532 108316 288584 108322
rect 288532 108258 288584 108264
rect 288348 99340 288400 99346
rect 288348 99282 288400 99288
rect 288360 98666 288388 99282
rect 288348 98660 288400 98666
rect 288348 98602 288400 98608
rect 288440 28280 288492 28286
rect 288440 28222 288492 28228
rect 288452 16574 288480 28222
rect 288452 16546 289032 16574
rect 287704 3528 287756 3534
rect 287704 3470 287756 3476
rect 287624 598 287836 626
rect 287624 490 287652 598
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287348 462 287652 490
rect 287808 480 287836 598
rect 289004 480 289032 16546
rect 289096 2990 289124 140830
rect 295340 120760 295392 120766
rect 295340 120702 295392 120708
rect 291844 111104 291896 111110
rect 291844 111046 291896 111052
rect 291200 54528 291252 54534
rect 291200 54470 291252 54476
rect 290464 42084 290516 42090
rect 290464 42026 290516 42032
rect 290476 3534 290504 42026
rect 291212 16574 291240 54470
rect 291212 16546 291424 16574
rect 290188 3528 290240 3534
rect 290188 3470 290240 3476
rect 290464 3528 290516 3534
rect 290464 3470 290516 3476
rect 289084 2984 289136 2990
rect 289084 2926 289136 2932
rect 290200 480 290228 3470
rect 291396 480 291424 16546
rect 291856 4486 291884 111046
rect 292672 53100 292724 53106
rect 292672 53042 292724 53048
rect 292684 16574 292712 53042
rect 295352 16574 295380 120702
rect 292684 16546 293264 16574
rect 295352 16546 295656 16574
rect 291844 4480 291896 4486
rect 291844 4422 291896 4428
rect 292580 2984 292632 2990
rect 292580 2926 292632 2932
rect 292592 480 292620 2926
rect 293236 490 293264 16546
rect 294880 3528 294932 3534
rect 294880 3470 294932 3476
rect 293512 598 293724 626
rect 293512 490 293540 598
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293236 462 293540 490
rect 293696 480 293724 598
rect 294892 480 294920 3470
rect 295628 490 295656 16546
rect 295996 3466 296024 175306
rect 306380 163532 306432 163538
rect 306380 163474 306432 163480
rect 302240 152516 302292 152522
rect 302240 152458 302292 152464
rect 298744 145580 298796 145586
rect 298744 145522 298796 145528
rect 298098 87544 298154 87553
rect 298098 87479 298154 87488
rect 297272 4480 297324 4486
rect 297272 4422 297324 4428
rect 295984 3460 296036 3466
rect 295984 3402 296036 3408
rect 295904 598 296116 626
rect 295904 490 295932 598
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 295628 462 295932 490
rect 296088 480 296116 598
rect 297284 480 297312 4422
rect 298112 490 298140 87479
rect 298756 6254 298784 145522
rect 299480 129056 299532 129062
rect 299480 128998 299532 129004
rect 298744 6248 298796 6254
rect 298744 6190 298796 6196
rect 299492 3534 299520 128998
rect 299480 3528 299532 3534
rect 299480 3470 299532 3476
rect 300768 3528 300820 3534
rect 300768 3470 300820 3476
rect 299664 3120 299716 3126
rect 299664 3062 299716 3068
rect 298296 598 298508 626
rect 298296 490 298324 598
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298112 462 298324 490
rect 298480 480 298508 598
rect 299676 480 299704 3062
rect 300780 480 300808 3470
rect 301964 3460 302016 3466
rect 301964 3402 302016 3408
rect 301976 480 302004 3402
rect 302252 3126 302280 152458
rect 305000 150544 305052 150550
rect 305000 150486 305052 150492
rect 304264 117972 304316 117978
rect 304264 117914 304316 117920
rect 303618 24168 303674 24177
rect 303618 24103 303674 24112
rect 303632 16574 303660 24103
rect 303632 16546 303936 16574
rect 303160 6180 303212 6186
rect 303160 6122 303212 6128
rect 302240 3120 302292 3126
rect 302240 3062 302292 3068
rect 303172 480 303200 6122
rect 303908 490 303936 16546
rect 304276 4826 304304 117914
rect 305012 6914 305040 150486
rect 304920 6886 305040 6914
rect 304264 4820 304316 4826
rect 304264 4762 304316 4768
rect 304920 3534 304948 6886
rect 304908 3528 304960 3534
rect 304908 3470 304960 3476
rect 305552 3528 305604 3534
rect 305552 3470 305604 3476
rect 304184 598 304396 626
rect 304184 490 304212 598
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 303908 462 304212 490
rect 304368 480 304396 598
rect 305564 480 305592 3470
rect 306392 490 306420 163474
rect 307760 21412 307812 21418
rect 307760 21354 307812 21360
rect 307772 3534 307800 21354
rect 309796 5574 309824 297327
rect 565084 271924 565136 271930
rect 565084 271866 565136 271872
rect 565096 241466 565124 271866
rect 574756 244225 574784 351902
rect 580170 351863 580226 351872
rect 580906 325272 580962 325281
rect 580906 325207 580962 325216
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 580184 311914 580212 312015
rect 580172 311908 580224 311914
rect 580172 311850 580224 311856
rect 580920 299470 580948 325207
rect 580908 299464 580960 299470
rect 580908 299406 580960 299412
rect 580262 298752 580318 298761
rect 580262 298687 580318 298696
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 580184 271930 580212 272167
rect 580172 271924 580224 271930
rect 580172 271866 580224 271872
rect 580276 256018 580304 298687
rect 582392 260166 582420 643991
rect 582470 630864 582526 630873
rect 582470 630799 582526 630808
rect 582380 260160 582432 260166
rect 582380 260102 582432 260108
rect 582378 258904 582434 258913
rect 582378 258839 582434 258848
rect 580264 256012 580316 256018
rect 580264 255954 580316 255960
rect 582392 250510 582420 258839
rect 582484 258738 582512 630799
rect 582654 617536 582710 617545
rect 582654 617471 582710 617480
rect 582668 585818 582696 617471
rect 582656 585812 582708 585818
rect 582656 585754 582708 585760
rect 582654 577688 582710 577697
rect 582654 577623 582710 577632
rect 582472 258732 582524 258738
rect 582472 258674 582524 258680
rect 582380 250504 582432 250510
rect 582380 250446 582432 250452
rect 582380 248464 582432 248470
rect 582432 248412 582512 248414
rect 582380 248406 582512 248412
rect 582392 248386 582512 248406
rect 582380 247104 582432 247110
rect 582380 247046 582432 247052
rect 574742 244216 574798 244225
rect 574742 244151 574798 244160
rect 565084 241460 565136 241466
rect 565084 241402 565136 241408
rect 580172 233300 580224 233306
rect 580172 233242 580224 233248
rect 580184 232393 580212 233242
rect 580170 232384 580226 232393
rect 580170 232319 580226 232328
rect 580264 229764 580316 229770
rect 580264 229706 580316 229712
rect 580276 205737 580304 229706
rect 582392 219065 582420 247046
rect 582484 245585 582512 248386
rect 582470 245576 582526 245585
rect 582470 245511 582526 245520
rect 582564 241528 582616 241534
rect 582564 241470 582616 241476
rect 582470 236600 582526 236609
rect 582470 236535 582526 236544
rect 582378 219056 582434 219065
rect 582378 218991 582434 219000
rect 580262 205728 580318 205737
rect 580262 205663 580318 205672
rect 580170 192536 580226 192545
rect 580170 192471 580172 192480
rect 580224 192471 580226 192480
rect 580172 192442 580224 192448
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580184 178702 580212 179143
rect 580172 178696 580224 178702
rect 580172 178638 580224 178644
rect 340142 160712 340198 160721
rect 340142 160647 340198 160656
rect 317420 155236 317472 155242
rect 317420 155178 317472 155184
rect 313280 143608 313332 143614
rect 313280 143550 313332 143556
rect 313292 16574 313320 143550
rect 316040 124908 316092 124914
rect 316040 124850 316092 124856
rect 316052 16574 316080 124850
rect 317432 16574 317460 155178
rect 320180 147756 320232 147762
rect 320180 147698 320232 147704
rect 313292 16546 313872 16574
rect 316052 16546 316264 16574
rect 317432 16546 318104 16574
rect 312176 11756 312228 11762
rect 312176 11698 312228 11704
rect 310244 6248 310296 6254
rect 310244 6190 310296 6196
rect 309784 5568 309836 5574
rect 309784 5510 309836 5516
rect 307944 4820 307996 4826
rect 307944 4762 307996 4768
rect 307760 3528 307812 3534
rect 307760 3470 307812 3476
rect 306576 598 306788 626
rect 306576 490 306604 598
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306392 462 306604 490
rect 306760 480 306788 598
rect 307956 480 307984 4762
rect 309048 3528 309100 3534
rect 309048 3470 309100 3476
rect 309060 480 309088 3470
rect 310256 480 310284 6190
rect 311440 5568 311492 5574
rect 311440 5510 311492 5516
rect 311452 480 311480 5510
rect 312188 490 312216 11698
rect 312464 598 312676 626
rect 312464 490 312492 598
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312188 462 312492 490
rect 312648 480 312676 598
rect 313844 480 313872 16546
rect 315028 9036 315080 9042
rect 315028 8978 315080 8984
rect 315040 480 315068 8978
rect 316236 480 316264 16546
rect 317328 7608 317380 7614
rect 317328 7550 317380 7556
rect 317340 480 317368 7550
rect 318076 490 318104 16546
rect 320192 3534 320220 147698
rect 322204 138712 322256 138718
rect 322204 138654 322256 138660
rect 321560 22772 321612 22778
rect 321560 22714 321612 22720
rect 320272 19984 320324 19990
rect 320272 19926 320324 19932
rect 320284 16574 320312 19926
rect 321572 16574 321600 22714
rect 320284 16546 320496 16574
rect 321572 16546 322152 16574
rect 319720 3528 319772 3534
rect 319720 3470 319772 3476
rect 320180 3528 320232 3534
rect 320180 3470 320232 3476
rect 318352 598 318564 626
rect 318352 490 318380 598
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 462 318380 490
rect 318536 480 318564 598
rect 319732 480 319760 3470
rect 320468 490 320496 16546
rect 320744 598 320956 626
rect 320744 490 320772 598
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320468 462 320772 490
rect 320928 480 320956 598
rect 322124 480 322152 16546
rect 322216 4010 322244 138654
rect 323584 127628 323636 127634
rect 323584 127570 323636 127576
rect 322940 31068 322992 31074
rect 322940 31010 322992 31016
rect 322204 4004 322256 4010
rect 322204 3946 322256 3952
rect 322952 490 322980 31010
rect 323596 4826 323624 127570
rect 324320 111852 324372 111858
rect 324320 111794 324372 111800
rect 323584 4820 323636 4826
rect 323584 4762 323636 4768
rect 324332 3534 324360 111794
rect 327724 100020 327776 100026
rect 327724 99962 327776 99968
rect 327080 68332 327132 68338
rect 327080 68274 327132 68280
rect 324412 36576 324464 36582
rect 324412 36518 324464 36524
rect 324320 3528 324372 3534
rect 324320 3470 324372 3476
rect 323136 598 323348 626
rect 323136 490 323164 598
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 322952 462 323164 490
rect 323320 480 323348 598
rect 324424 480 324452 36518
rect 327092 16574 327120 68274
rect 327092 16546 327672 16574
rect 326804 4004 326856 4010
rect 326804 3946 326856 3952
rect 325608 3528 325660 3534
rect 325608 3470 325660 3476
rect 325620 480 325648 3470
rect 326816 480 326844 3946
rect 327644 2802 327672 16546
rect 327736 2990 327764 99962
rect 331220 98660 331272 98666
rect 331220 98602 331272 98608
rect 328460 51740 328512 51746
rect 328460 51682 328512 51688
rect 328472 16574 328500 51682
rect 328472 16546 328776 16574
rect 327724 2984 327776 2990
rect 327724 2926 327776 2932
rect 327644 2774 328040 2802
rect 328012 480 328040 2774
rect 328748 490 328776 16546
rect 330392 13116 330444 13122
rect 330392 13058 330444 13064
rect 329024 598 329236 626
rect 329024 490 329052 598
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 328748 462 329052 490
rect 329208 480 329236 598
rect 330404 480 330432 13058
rect 331232 490 331260 98602
rect 335358 83464 335414 83473
rect 335358 83399 335414 83408
rect 332692 44872 332744 44878
rect 332692 44814 332744 44820
rect 332704 11762 332732 44814
rect 333980 37936 334032 37942
rect 333980 37878 334032 37884
rect 333992 16574 334020 37878
rect 335372 16574 335400 83399
rect 338120 40724 338172 40730
rect 338120 40666 338172 40672
rect 338132 16574 338160 40666
rect 333992 16546 334664 16574
rect 335372 16546 336320 16574
rect 338132 16546 338712 16574
rect 332692 11756 332744 11762
rect 332692 11698 332744 11704
rect 333888 11756 333940 11762
rect 333888 11698 333940 11704
rect 332692 2984 332744 2990
rect 332692 2926 332744 2932
rect 331416 598 331628 626
rect 331416 490 331444 598
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331232 462 331444 490
rect 331600 480 331628 598
rect 332704 480 332732 2926
rect 333900 480 333928 11698
rect 334636 490 334664 16546
rect 334912 598 335124 626
rect 334912 490 334940 598
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 462 334940 490
rect 335096 480 335124 598
rect 336292 480 336320 16546
rect 337476 4820 337528 4826
rect 337476 4762 337528 4768
rect 337488 480 337516 4762
rect 338684 480 338712 16546
rect 340156 3534 340184 160647
rect 580356 158024 580408 158030
rect 580356 157966 580408 157972
rect 580264 146940 580316 146946
rect 580264 146882 580316 146888
rect 341522 135960 341578 135969
rect 341522 135895 341578 135904
rect 340972 32428 341024 32434
rect 340972 32370 341024 32376
rect 340144 3528 340196 3534
rect 340144 3470 340196 3476
rect 339868 2984 339920 2990
rect 339868 2926 339920 2932
rect 339880 480 339908 2926
rect 340984 480 341012 32370
rect 341536 3466 341564 135895
rect 349160 126268 349212 126274
rect 349160 126210 349212 126216
rect 342352 84244 342404 84250
rect 342352 84186 342404 84192
rect 342260 10328 342312 10334
rect 342260 10270 342312 10276
rect 342168 3528 342220 3534
rect 342168 3470 342220 3476
rect 341524 3460 341576 3466
rect 341524 3402 341576 3408
rect 342180 480 342208 3470
rect 342272 2666 342300 10270
rect 342364 2990 342392 84186
rect 345018 64152 345074 64161
rect 345018 64087 345074 64096
rect 343640 47592 343692 47598
rect 343640 47534 343692 47540
rect 343652 16574 343680 47534
rect 345032 16574 345060 64087
rect 343652 16546 344600 16574
rect 345032 16546 345336 16574
rect 342352 2984 342404 2990
rect 342352 2926 342404 2932
rect 342272 2638 342944 2666
rect 342916 490 342944 2638
rect 343192 598 343404 626
rect 343192 490 343220 598
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 462 343220 490
rect 343376 480 343404 598
rect 344572 480 344600 16546
rect 345308 490 345336 16546
rect 349172 5574 349200 126210
rect 580276 126041 580304 146882
rect 580368 139369 580396 157966
rect 580354 139360 580410 139369
rect 580354 139295 580410 139304
rect 580262 126032 580318 126041
rect 580262 125967 580318 125976
rect 353300 106344 353352 106350
rect 353300 106286 353352 106292
rect 351920 62824 351972 62830
rect 351920 62766 351972 62772
rect 348056 5568 348108 5574
rect 348056 5510 348108 5516
rect 349160 5568 349212 5574
rect 349160 5510 349212 5516
rect 346952 4208 347004 4214
rect 346952 4150 347004 4156
rect 345584 598 345796 626
rect 345584 490 345612 598
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345308 462 345612 490
rect 345768 480 345796 598
rect 346964 480 346992 4150
rect 348068 480 348096 5510
rect 351644 4140 351696 4146
rect 351644 4082 351696 4088
rect 350448 3460 350500 3466
rect 350448 3402 350500 3408
rect 349252 3188 349304 3194
rect 349252 3130 349304 3136
rect 349264 480 349292 3130
rect 350460 480 350488 3402
rect 351656 480 351684 4082
rect 351932 3194 351960 62766
rect 353312 4214 353340 106286
rect 582378 99512 582434 99521
rect 582378 99447 582434 99456
rect 580262 90400 580318 90409
rect 580262 90335 580318 90344
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 580276 73001 580304 90335
rect 582392 89729 582420 99447
rect 582378 89720 582434 89729
rect 582378 89655 582434 89664
rect 580262 72992 580318 73001
rect 580262 72927 580318 72936
rect 356060 72480 356112 72486
rect 356060 72422 356112 72428
rect 353300 4208 353352 4214
rect 353300 4150 353352 4156
rect 356072 4146 356100 72422
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 582484 6914 582512 236535
rect 582576 152697 582604 241470
rect 582668 227730 582696 577623
rect 582760 570654 582788 683839
rect 583666 590744 583722 590753
rect 583666 590679 583722 590688
rect 582840 583772 582892 583778
rect 582840 583714 582892 583720
rect 582748 570648 582800 570654
rect 582748 570590 582800 570596
rect 582852 564369 582880 583714
rect 582838 564360 582894 564369
rect 582838 564295 582894 564304
rect 582838 537840 582894 537849
rect 582838 537775 582894 537784
rect 582746 524512 582802 524521
rect 582746 524447 582802 524456
rect 582760 231810 582788 524447
rect 582852 258058 582880 537775
rect 582930 484664 582986 484673
rect 582930 484599 582986 484608
rect 582840 258052 582892 258058
rect 582840 257994 582892 258000
rect 582944 235929 582972 484599
rect 583022 471472 583078 471481
rect 583022 471407 583078 471416
rect 583036 255270 583064 471407
rect 583114 458144 583170 458153
rect 583114 458079 583170 458088
rect 583128 438190 583156 458079
rect 583116 438184 583168 438190
rect 583116 438126 583168 438132
rect 583206 431624 583262 431633
rect 583206 431559 583262 431568
rect 583114 289096 583170 289105
rect 583114 289031 583170 289040
rect 583024 255264 583076 255270
rect 583024 255206 583076 255212
rect 582930 235920 582986 235929
rect 582930 235855 582986 235864
rect 582930 232520 582986 232529
rect 582930 232455 582986 232464
rect 582748 231804 582800 231810
rect 582748 231746 582800 231752
rect 582656 227724 582708 227730
rect 582656 227666 582708 227672
rect 582746 165880 582802 165889
rect 582746 165815 582802 165824
rect 582656 161492 582708 161498
rect 582656 161434 582708 161440
rect 582562 152688 582618 152697
rect 582562 152623 582618 152632
rect 582562 138680 582618 138689
rect 582562 138615 582618 138624
rect 582576 19825 582604 138615
rect 582668 59673 582696 161434
rect 582760 124166 582788 165815
rect 582838 142760 582894 142769
rect 582838 142695 582894 142704
rect 582748 124160 582800 124166
rect 582748 124102 582800 124108
rect 582852 112849 582880 142695
rect 582838 112840 582894 112849
rect 582838 112775 582894 112784
rect 582748 82136 582800 82142
rect 582748 82078 582800 82084
rect 582654 59664 582710 59673
rect 582654 59599 582710 59608
rect 582562 19816 582618 19825
rect 582562 19751 582618 19760
rect 582392 6886 582512 6914
rect 356060 4140 356112 4146
rect 356060 4082 356112 4088
rect 582392 3482 582420 6886
rect 582760 6633 582788 82078
rect 582840 79348 582892 79354
rect 582840 79290 582892 79296
rect 582852 33153 582880 79290
rect 582838 33144 582894 33153
rect 582838 33079 582894 33088
rect 582944 16574 582972 232455
rect 582944 16546 583064 16574
rect 582746 6624 582802 6633
rect 582746 6559 582802 6568
rect 582208 3454 582420 3482
rect 351920 3188 351972 3194
rect 351920 3130 351972 3136
rect 581000 2984 581052 2990
rect 581000 2926 581052 2932
rect 581012 480 581040 2926
rect 582208 480 582236 3454
rect 583036 2530 583064 16546
rect 583128 2990 583156 289031
rect 583220 253910 583248 431559
rect 583390 418296 583446 418305
rect 583390 418231 583446 418240
rect 583298 404968 583354 404977
rect 583298 404903 583354 404912
rect 583208 253904 583260 253910
rect 583208 253846 583260 253852
rect 583312 240145 583340 404903
rect 583404 255202 583432 418231
rect 583482 378176 583538 378185
rect 583482 378111 583538 378120
rect 583392 255196 583444 255202
rect 583392 255138 583444 255144
rect 583496 253201 583524 378111
rect 583576 299464 583628 299470
rect 583576 299406 583628 299412
rect 583482 253192 583538 253201
rect 583482 253127 583538 253136
rect 583588 251870 583616 299406
rect 583576 251864 583628 251870
rect 583576 251806 583628 251812
rect 583298 240136 583354 240145
rect 583298 240071 583354 240080
rect 583680 238649 583708 590679
rect 583666 238640 583722 238649
rect 583666 238575 583722 238584
rect 583116 2984 583168 2990
rect 583116 2926 583168 2932
rect 583036 2502 583432 2530
rect 583404 480 583432 2502
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 2778 606056 2834 606112
rect 3330 579944 3386 580000
rect 3514 671200 3570 671256
rect 3514 658144 3570 658200
rect 3514 632068 3516 632088
rect 3516 632068 3568 632088
rect 3568 632068 3570 632088
rect 3514 632032 3570 632068
rect 15842 621560 15898 621616
rect 3514 619112 3570 619168
rect 3422 566888 3478 566944
rect 3514 553852 3570 553888
rect 3514 553832 3516 553852
rect 3516 553832 3568 553852
rect 3568 553832 3570 553852
rect 4802 542408 4858 542464
rect 17222 541048 17278 541104
rect 3514 527876 3570 527912
rect 3514 527856 3516 527876
rect 3516 527856 3568 527876
rect 3568 527856 3570 527876
rect 3514 514820 3570 514856
rect 3514 514800 3516 514820
rect 3516 514800 3568 514820
rect 3568 514800 3570 514820
rect 3422 501744 3478 501800
rect 3422 475632 3478 475688
rect 3146 449520 3202 449576
rect 2778 423580 2780 423600
rect 2780 423580 2832 423600
rect 2832 423580 2834 423600
rect 2778 423544 2834 423580
rect 2870 410488 2926 410544
rect 3514 462576 3570 462632
rect 3514 397432 3570 397488
rect 3422 371320 3478 371376
rect 14462 388728 14518 388784
rect 3330 358400 3386 358456
rect 3330 345344 3386 345400
rect 12346 328480 12402 328536
rect 3422 319232 3478 319288
rect 1306 306720 1362 306776
rect 3238 306176 3294 306232
rect 4066 297336 4122 297392
rect 3422 293120 3478 293176
rect 3514 267144 3570 267200
rect 3146 254088 3202 254144
rect 3514 241032 3570 241088
rect 3422 214920 3478 214976
rect 3330 201864 3386 201920
rect 3146 149776 3202 149832
rect 3514 188808 3570 188864
rect 3514 162868 3516 162888
rect 3516 162868 3568 162888
rect 3568 162868 3570 162888
rect 3514 162832 3570 162868
rect 3514 136720 3570 136776
rect 3146 110608 3202 110664
rect 3054 97552 3110 97608
rect 3422 84632 3478 84688
rect 3422 71576 3478 71632
rect 3514 58520 3570 58576
rect 3422 45500 3424 45520
rect 3424 45500 3476 45520
rect 3476 45500 3478 45520
rect 3422 45464 3478 45500
rect 2870 32408 2926 32464
rect 3422 19352 3478 19408
rect 3422 6432 3478 6488
rect 12254 298832 12310 298888
rect 5446 196560 5502 196616
rect 8758 3304 8814 3360
rect 17866 309168 17922 309224
rect 16486 301280 16542 301336
rect 15106 235184 15162 235240
rect 13726 226888 13782 226944
rect 18694 241168 18750 241224
rect 21362 236000 21418 236056
rect 18602 233416 18658 233472
rect 19246 211792 19302 211848
rect 19430 4800 19486 4856
rect 30286 311888 30342 311944
rect 26146 294480 26202 294536
rect 24766 221448 24822 221504
rect 28906 232464 28962 232520
rect 29642 224168 29698 224224
rect 31022 302776 31078 302832
rect 39854 531936 39910 531992
rect 35162 313384 35218 313440
rect 34426 310528 34482 310584
rect 32402 253816 32458 253872
rect 39302 314744 39358 314800
rect 37186 310664 37242 310720
rect 35806 254496 35862 254552
rect 35806 222808 35862 222864
rect 35162 3304 35218 3360
rect 39854 269728 39910 269784
rect 43994 530576 44050 530632
rect 41234 242936 41290 242992
rect 39946 120672 40002 120728
rect 42706 218592 42762 218648
rect 41326 204856 41382 204912
rect 41234 91704 41290 91760
rect 45466 210296 45522 210352
rect 45374 199280 45430 199336
rect 48134 436056 48190 436112
rect 48042 385600 48098 385656
rect 46846 258712 46902 258768
rect 48134 254088 48190 254144
rect 49606 266464 49662 266520
rect 49514 217232 49570 217288
rect 48226 206216 48282 206272
rect 50526 264968 50582 265024
rect 50894 268368 50950 268424
rect 50894 264968 50950 265024
rect 51722 389136 51778 389192
rect 52182 384240 52238 384296
rect 52090 285912 52146 285968
rect 50894 231784 50950 231840
rect 50710 153040 50766 153096
rect 50710 151816 50766 151872
rect 51998 223488 52054 223544
rect 54942 433472 54998 433528
rect 53470 391448 53526 391504
rect 52274 239808 52330 239864
rect 52366 238040 52422 238096
rect 52274 223488 52330 223544
rect 52274 222264 52330 222320
rect 52090 175344 52146 175400
rect 50802 150728 50858 150784
rect 50894 148280 50950 148336
rect 53746 251232 53802 251288
rect 53654 149640 53710 149696
rect 53562 149096 53618 149152
rect 52366 90888 52422 90944
rect 54942 289720 54998 289776
rect 55126 289720 55182 289776
rect 55034 211112 55090 211168
rect 54942 157392 54998 157448
rect 54482 136040 54538 136096
rect 59266 581168 59322 581224
rect 57610 290400 57666 290456
rect 55034 95784 55090 95840
rect 57702 244432 57758 244488
rect 57702 212608 57758 212664
rect 57886 244432 57942 244488
rect 59082 277616 59138 277672
rect 60370 271904 60426 271960
rect 59174 228928 59230 228984
rect 59082 143520 59138 143576
rect 56506 89664 56562 89720
rect 57242 86536 57298 86592
rect 60554 273264 60610 273320
rect 60646 270544 60702 270600
rect 61014 251232 61070 251288
rect 61934 432792 61990 432848
rect 61750 284280 61806 284336
rect 61658 283192 61714 283248
rect 61750 273264 61806 273320
rect 63406 578856 63462 578912
rect 63314 434696 63370 434752
rect 63038 268368 63094 268424
rect 62026 263608 62082 263664
rect 61842 248512 61898 248568
rect 61934 248240 61990 248296
rect 61934 216688 61990 216744
rect 61842 169768 61898 169824
rect 60554 160792 60610 160848
rect 60646 155216 60702 155272
rect 57886 73072 57942 73128
rect 57242 71848 57298 71904
rect 57886 71848 57942 71904
rect 62118 241576 62174 241632
rect 63406 420824 63462 420880
rect 65982 568792 66038 568848
rect 66810 579944 66866 580000
rect 66810 578584 66866 578640
rect 66534 575864 66590 575920
rect 66442 573144 66498 573200
rect 66718 571784 66774 571840
rect 66718 564712 66774 564768
rect 66442 564168 66498 564224
rect 66166 561992 66222 562048
rect 66074 545944 66130 546000
rect 65890 449928 65946 449984
rect 63130 144880 63186 144936
rect 62026 139440 62082 139496
rect 63406 241576 63462 241632
rect 63314 142160 63370 142216
rect 64694 284280 64750 284336
rect 64694 274760 64750 274816
rect 64602 239944 64658 240000
rect 66074 429256 66130 429312
rect 65982 403688 66038 403744
rect 65706 265140 65708 265160
rect 65708 265140 65760 265160
rect 65760 265140 65762 265160
rect 65706 265104 65762 265140
rect 64786 263608 64842 263664
rect 64602 138760 64658 138816
rect 66534 549480 66590 549536
rect 66718 544584 66774 544640
rect 66258 433356 66314 433392
rect 66258 433336 66260 433356
rect 66260 433336 66312 433356
rect 66312 433336 66314 433356
rect 66442 432520 66498 432576
rect 66718 431432 66774 431488
rect 66718 430344 66774 430400
rect 66718 428168 66774 428224
rect 66718 427352 66774 427408
rect 66534 425176 66590 425232
rect 66718 424088 66774 424144
rect 66718 423272 66774 423328
rect 66626 418920 66682 418976
rect 66626 415928 66682 415984
rect 66718 414840 66774 414896
rect 66718 411848 66774 411904
rect 66258 408856 66314 408912
rect 66442 406680 66498 406736
rect 67454 577224 67510 577280
rect 66902 570152 66958 570208
rect 66994 567432 67050 567488
rect 66994 560632 67050 560688
rect 66994 559272 67050 559328
rect 66994 557912 67050 557968
rect 66994 555192 67050 555248
rect 66994 553560 67050 553616
rect 66994 546760 67050 546816
rect 66994 421096 67050 421152
rect 66902 420008 66958 420064
rect 66994 418104 67050 418160
rect 67362 418104 67418 418160
rect 66902 417016 66958 417072
rect 66902 414024 66958 414080
rect 66902 412936 66958 412992
rect 66902 410760 66958 410816
rect 66902 407768 66958 407824
rect 67546 575320 67602 575376
rect 76470 591096 76526 591152
rect 77206 591096 77262 591152
rect 71778 584840 71834 584896
rect 72422 582664 72478 582720
rect 69478 582392 69534 582448
rect 70306 582392 70362 582448
rect 74906 582392 74962 582448
rect 77206 590688 77262 590744
rect 75366 580896 75422 580952
rect 70858 580760 70914 580816
rect 79046 581032 79102 581088
rect 83002 581168 83058 581224
rect 88246 582528 88302 582584
rect 79782 580760 79838 580816
rect 84198 580760 84254 580816
rect 88706 580760 88762 580816
rect 92386 580760 92442 580816
rect 68650 578856 68706 578912
rect 67638 566616 67694 566672
rect 67822 556552 67878 556608
rect 67730 552200 67786 552256
rect 67638 550840 67694 550896
rect 95238 574776 95294 574832
rect 94778 563624 94834 563680
rect 94686 552472 94742 552528
rect 94686 540232 94742 540288
rect 70306 539708 70362 539744
rect 70306 539688 70308 539708
rect 70308 539688 70360 539708
rect 70360 539688 70362 539708
rect 67454 405592 67510 405648
rect 66902 404504 66958 404560
rect 66718 402600 66774 402656
rect 66534 399608 66590 399664
rect 66626 398520 66682 398576
rect 66902 401512 66958 401568
rect 66810 400424 66866 400480
rect 67086 396344 67142 396400
rect 66810 395256 66866 395312
rect 66166 394576 66222 394632
rect 66350 394440 66406 394496
rect 66810 393372 66866 393408
rect 66810 393352 66812 393372
rect 66812 393352 66864 393372
rect 66864 393352 66866 393372
rect 66810 392264 66866 392320
rect 66810 391176 66866 391232
rect 68926 449948 68982 449984
rect 68926 449928 68928 449948
rect 68928 449928 68980 449948
rect 68980 449928 68982 449948
rect 68926 436192 68982 436248
rect 71042 436192 71098 436248
rect 69938 436056 69994 436112
rect 76746 539552 76802 539608
rect 72606 476720 72662 476776
rect 74446 534656 74502 534712
rect 73434 434696 73490 434752
rect 76470 536696 76526 536752
rect 76470 535608 76526 535664
rect 76102 535472 76158 535528
rect 77206 535608 77262 535664
rect 76746 535472 76802 535528
rect 76562 522280 76618 522336
rect 76102 441632 76158 441688
rect 77390 437144 77446 437200
rect 77482 436328 77538 436384
rect 77390 436192 77446 436248
rect 74722 434288 74778 434344
rect 76194 434288 76250 434344
rect 78402 437416 78458 437472
rect 78034 437144 78090 437200
rect 81438 479440 81494 479496
rect 80058 450472 80114 450528
rect 81346 438096 81402 438152
rect 80242 435240 80298 435296
rect 81346 434424 81402 434480
rect 83738 436056 83794 436112
rect 68926 433608 68982 433664
rect 83186 433744 83242 433800
rect 75458 433608 75514 433664
rect 78218 433608 78274 433664
rect 78954 433608 79010 433664
rect 83094 433608 83150 433664
rect 84474 433608 84530 433664
rect 85670 436056 85726 436112
rect 88430 468560 88486 468616
rect 93950 538872 94006 538928
rect 88430 440272 88486 440328
rect 86314 436056 86370 436112
rect 87142 436056 87198 436112
rect 88246 436056 88302 436112
rect 89902 436192 89958 436248
rect 94778 474000 94834 474056
rect 96250 574776 96306 574832
rect 96894 578856 96950 578912
rect 97078 577496 97134 577552
rect 97906 576716 97908 576736
rect 97908 576716 97960 576736
rect 97960 576716 97962 576736
rect 97906 576680 97962 576716
rect 97906 573416 97962 573472
rect 97262 572192 97318 572248
rect 96618 569064 96674 569120
rect 95422 565800 95478 565856
rect 95330 558864 95386 558920
rect 95330 555464 95386 555520
rect 96802 560904 96858 560960
rect 95882 558864 95938 558920
rect 95330 523640 95386 523696
rect 96710 556824 96766 556880
rect 96618 552064 96674 552120
rect 97906 570016 97962 570072
rect 97906 569064 97962 569120
rect 97354 562264 97410 562320
rect 96894 554104 96950 554160
rect 96986 552744 97042 552800
rect 96710 545672 96766 545728
rect 94502 437552 94558 437608
rect 94410 436056 94466 436112
rect 95284 434560 95340 434616
rect 94778 434288 94834 434344
rect 96342 434288 96398 434344
rect 97906 550704 97962 550760
rect 97538 544312 97594 544368
rect 98090 542952 98146 543008
rect 100022 582528 100078 582584
rect 98642 439456 98698 439512
rect 97078 437416 97134 437472
rect 102782 581032 102838 581088
rect 100758 436328 100814 436384
rect 92662 434152 92718 434208
rect 96986 434152 97042 434208
rect 91466 433880 91522 433936
rect 99194 433880 99250 433936
rect 87326 433744 87382 433800
rect 92938 433744 92994 433800
rect 98366 433744 98422 433800
rect 103334 436328 103390 436384
rect 103334 436056 103390 436112
rect 85670 433608 85726 433664
rect 85946 433608 86002 433664
rect 87142 433608 87198 433664
rect 87970 433608 88026 433664
rect 89994 433608 90050 433664
rect 91374 433608 91430 433664
rect 98458 433608 98514 433664
rect 99930 433608 99986 433664
rect 101218 433608 101274 433664
rect 102690 433608 102746 433664
rect 104898 436192 104954 436248
rect 104346 436056 104402 436112
rect 107566 437416 107622 437472
rect 110418 436328 110474 436384
rect 109406 434288 109462 434344
rect 108946 434016 109002 434072
rect 104162 433608 104218 433664
rect 105450 433608 105506 433664
rect 106738 433608 106794 433664
rect 110878 433644 110880 433664
rect 110880 433644 110932 433664
rect 110932 433644 110934 433664
rect 110878 433608 110934 433644
rect 111890 433608 111946 433664
rect 68650 432792 68706 432848
rect 67730 397840 67786 397896
rect 67270 312160 67326 312216
rect 66902 312024 66958 312080
rect 67454 396344 67510 396400
rect 66442 291080 66498 291136
rect 66902 291080 66958 291136
rect 66442 290400 66498 290456
rect 66074 271904 66130 271960
rect 66074 252728 66130 252784
rect 65982 147736 66038 147792
rect 65890 144744 65946 144800
rect 65890 143656 65946 143712
rect 66810 282920 66866 282976
rect 66534 278840 66590 278896
rect 66810 278044 66866 278080
rect 66810 278024 66812 278044
rect 66812 278024 66864 278044
rect 66864 278024 66866 278044
rect 66810 277208 66866 277264
rect 66902 276392 66958 276448
rect 66626 275576 66682 275632
rect 66810 273128 66866 273184
rect 66258 270680 66314 270736
rect 66810 268232 66866 268288
rect 66810 266600 66866 266656
rect 66902 263336 66958 263392
rect 66534 262520 66590 262576
rect 66258 260888 66314 260944
rect 66810 260072 66866 260128
rect 66442 258032 66498 258088
rect 66810 257624 66866 257680
rect 66258 256808 66314 256864
rect 66810 255992 66866 256048
rect 66810 254360 66866 254416
rect 66534 252728 66590 252784
rect 66258 251912 66314 251968
rect 66810 251096 66866 251152
rect 66902 250280 66958 250336
rect 66810 248648 66866 248704
rect 66902 247832 66958 247888
rect 67178 247016 67234 247072
rect 66258 243752 66314 243808
rect 66810 242936 66866 242992
rect 66166 226344 66222 226400
rect 65982 118360 66038 118416
rect 65890 114552 65946 114608
rect 64602 92384 64658 92440
rect 66258 131960 66314 132016
rect 66350 131144 66406 131200
rect 66810 127608 66866 127664
rect 66810 125976 66866 126032
rect 66810 124344 66866 124400
rect 66902 123800 66958 123856
rect 66626 122984 66682 123040
rect 66810 122168 66866 122224
rect 66810 121388 66812 121408
rect 66812 121388 66864 121408
rect 66864 121388 66866 121408
rect 66810 121352 66866 121388
rect 66902 120672 66958 120728
rect 66626 120536 66682 120592
rect 66810 120028 66812 120048
rect 66812 120028 66864 120048
rect 66864 120028 66866 120048
rect 66810 119992 66866 120028
rect 66902 119176 66958 119232
rect 66258 117544 66314 117600
rect 66902 117000 66958 117056
rect 66258 116184 66314 116240
rect 66810 115368 66866 115424
rect 66810 113736 66866 113792
rect 66902 113192 66958 113248
rect 66166 111560 66222 111616
rect 66074 103128 66130 103184
rect 65982 82728 66038 82784
rect 62026 77832 62082 77888
rect 66626 110744 66682 110800
rect 66810 110200 66866 110256
rect 66810 108568 66866 108624
rect 66902 107752 66958 107808
rect 66810 106936 66866 106992
rect 66902 106392 66958 106448
rect 66534 105596 66590 105632
rect 66534 105576 66536 105596
rect 66536 105576 66588 105596
rect 66588 105576 66590 105596
rect 66258 104796 66260 104816
rect 66260 104796 66312 104816
rect 66312 104796 66314 104816
rect 66258 104760 66314 104796
rect 66534 102584 66590 102640
rect 66810 101768 66866 101824
rect 66442 100952 66498 101008
rect 66810 99592 66866 99648
rect 66626 98776 66682 98832
rect 67362 247016 67418 247072
rect 67362 246200 67418 246256
rect 68006 280472 68062 280528
rect 67546 244568 67602 244624
rect 67914 257896 67970 257952
rect 67638 233280 67694 233336
rect 67270 129784 67326 129840
rect 67178 97960 67234 98016
rect 66626 96328 66682 96384
rect 67546 147872 67602 147928
rect 67914 238584 67970 238640
rect 113270 431160 113326 431216
rect 113270 427080 113326 427136
rect 113178 420008 113234 420064
rect 112718 405864 112774 405920
rect 84382 390632 84438 390688
rect 70306 364384 70362 364440
rect 70214 317464 70270 317520
rect 69754 317328 69810 317384
rect 69754 316104 69810 316160
rect 69018 292576 69074 292632
rect 69110 285776 69166 285832
rect 69202 285640 69258 285696
rect 70306 317328 70362 317384
rect 69754 285776 69810 285832
rect 69202 283600 69258 283656
rect 71778 389000 71834 389056
rect 71226 387776 71282 387832
rect 71042 298696 71098 298752
rect 72330 390360 72386 390416
rect 72514 389000 72570 389056
rect 71870 388864 71926 388920
rect 73986 390360 74042 390416
rect 73158 387640 73214 387696
rect 73066 380160 73122 380216
rect 72422 313248 72478 313304
rect 71870 299512 71926 299568
rect 70766 283600 70822 283656
rect 71318 286048 71374 286104
rect 73066 299512 73122 299568
rect 71962 284144 72018 284200
rect 75274 387504 75330 387560
rect 77206 390360 77262 390416
rect 76010 389000 76066 389056
rect 76746 389000 76802 389056
rect 77298 387912 77354 387968
rect 75274 326984 75330 327040
rect 73526 304136 73582 304192
rect 73158 283464 73214 283520
rect 77022 318688 77078 318744
rect 76470 291216 76526 291272
rect 75274 285912 75330 285968
rect 74354 283192 74410 283248
rect 77482 385736 77538 385792
rect 79414 390360 79470 390416
rect 78862 389000 78918 389056
rect 80058 389000 80114 389056
rect 79874 383696 79930 383752
rect 79322 378664 79378 378720
rect 77206 365608 77262 365664
rect 77114 314880 77170 314936
rect 77114 291216 77170 291272
rect 78586 318280 78642 318336
rect 77206 289856 77262 289912
rect 79414 323584 79470 323640
rect 78126 286184 78182 286240
rect 79874 318008 79930 318064
rect 80978 389000 81034 389056
rect 81990 390360 82046 390416
rect 81438 388728 81494 388784
rect 81254 385600 81310 385656
rect 84106 375944 84162 376000
rect 83554 339516 83610 339552
rect 83554 339496 83556 339516
rect 83556 339496 83608 339516
rect 83608 339496 83610 339516
rect 84014 330384 84070 330440
rect 80702 320728 80758 320784
rect 81346 319368 81402 319424
rect 79506 286184 79562 286240
rect 80334 288360 80390 288416
rect 80334 287136 80390 287192
rect 81254 303592 81310 303648
rect 75734 283192 75790 283248
rect 81346 288360 81402 288416
rect 81530 318144 81586 318200
rect 82726 289076 82728 289096
rect 82728 289076 82780 289096
rect 82780 289076 82782 289096
rect 82726 289040 82782 289076
rect 82450 285640 82506 285696
rect 102414 390904 102470 390960
rect 106738 390904 106794 390960
rect 86866 380160 86922 380216
rect 84198 294616 84254 294672
rect 86774 288496 86830 288552
rect 85394 283600 85450 283656
rect 88338 389000 88394 389056
rect 87050 316648 87106 316704
rect 86958 293120 87014 293176
rect 89258 389000 89314 389056
rect 89626 385600 89682 385656
rect 89534 326304 89590 326360
rect 88246 319504 88302 319560
rect 89442 312432 89498 312488
rect 89534 288360 89590 288416
rect 89258 287272 89314 287328
rect 70950 282920 71006 282976
rect 80886 282920 80942 282976
rect 81254 282920 81310 282976
rect 87878 282920 87934 282976
rect 88522 282920 88578 282976
rect 91282 387776 91338 387832
rect 91006 373224 91062 373280
rect 90362 322904 90418 322960
rect 89718 300736 89774 300792
rect 89626 285640 89682 285696
rect 89810 283464 89866 283520
rect 92386 386960 92442 387016
rect 91374 383560 91430 383616
rect 91742 383560 91798 383616
rect 92294 308352 92350 308408
rect 93766 384240 93822 384296
rect 93674 353912 93730 353968
rect 92478 351872 92534 351928
rect 93030 293276 93086 293312
rect 93030 293256 93032 293276
rect 93032 293256 93084 293276
rect 93084 293256 93086 293276
rect 91374 285504 91430 285560
rect 91374 284416 91430 284472
rect 91466 284144 91522 284200
rect 92294 285504 92350 285560
rect 94410 387776 94466 387832
rect 94042 382200 94098 382256
rect 95330 389544 95386 389600
rect 97170 375944 97226 376000
rect 96526 374584 96582 374640
rect 95238 321408 95294 321464
rect 93766 287408 93822 287464
rect 93030 286048 93086 286104
rect 93674 286048 93730 286104
rect 92570 283464 92626 283520
rect 94134 286320 94190 286376
rect 96710 330248 96766 330304
rect 96020 283736 96076 283792
rect 100298 390224 100354 390280
rect 99654 389000 99710 389056
rect 100482 389000 100538 389056
rect 100758 389000 100814 389056
rect 97906 375944 97962 376000
rect 97814 330248 97870 330304
rect 97814 329840 97870 329896
rect 99286 332596 99288 332616
rect 99288 332596 99340 332616
rect 99340 332596 99342 332616
rect 99286 332560 99342 332596
rect 98090 327664 98146 327720
rect 97998 287408 98054 287464
rect 97906 282920 97962 282976
rect 69018 282684 69020 282704
rect 69020 282684 69072 282704
rect 69072 282684 69074 282704
rect 69018 282648 69074 282684
rect 68834 281152 68890 281208
rect 68558 279656 68614 279712
rect 98182 270680 98238 270736
rect 98090 247016 98146 247072
rect 69018 244296 69074 244352
rect 69478 241712 69534 241768
rect 70030 241576 70086 241632
rect 68006 229880 68062 229936
rect 69662 208392 69718 208448
rect 67730 133592 67786 133648
rect 67730 128968 67786 129024
rect 67638 112376 67694 112432
rect 67362 97144 67418 97200
rect 67454 95784 67510 95840
rect 67546 94152 67602 94208
rect 66166 74432 66222 74488
rect 64786 10240 64842 10296
rect 63222 3984 63278 4040
rect 67822 128152 67878 128208
rect 69294 137944 69350 138000
rect 69570 134952 69626 135008
rect 70306 141380 70308 141400
rect 70308 141380 70360 141400
rect 70360 141380 70362 141400
rect 70306 141344 70362 141380
rect 70950 241712 71006 241768
rect 72330 241712 72386 241768
rect 71042 241304 71098 241360
rect 71502 240760 71558 240816
rect 73894 241712 73950 241768
rect 83370 241712 83426 241768
rect 84934 241712 84990 241768
rect 72882 239944 72938 240000
rect 75550 241576 75606 241632
rect 74722 238040 74778 238096
rect 74538 230560 74594 230616
rect 72422 161608 72478 161664
rect 70858 137128 70914 137184
rect 72330 137808 72386 137864
rect 71686 137264 71742 137320
rect 73342 159296 73398 159352
rect 72422 137128 72478 137184
rect 73066 140800 73122 140856
rect 74262 141480 74318 141536
rect 76838 236000 76894 236056
rect 76562 213968 76618 214024
rect 75182 137808 75238 137864
rect 75826 138624 75882 138680
rect 75550 137944 75606 138000
rect 74998 135904 75054 135960
rect 79690 240080 79746 240136
rect 78678 236000 78734 236056
rect 77298 153720 77354 153776
rect 76654 140120 76710 140176
rect 76562 138760 76618 138816
rect 81346 241304 81402 241360
rect 79966 236816 80022 236872
rect 79966 236000 80022 236056
rect 80702 206352 80758 206408
rect 82082 240080 82138 240136
rect 84290 240080 84346 240136
rect 85946 241712 86002 241768
rect 86682 241712 86738 241768
rect 88062 241712 88118 241768
rect 84198 235864 84254 235920
rect 81346 141344 81402 141400
rect 82082 168408 82138 168464
rect 81990 146920 82046 146976
rect 82082 137944 82138 138000
rect 85578 236544 85634 236600
rect 86866 239944 86922 240000
rect 85486 145560 85542 145616
rect 84566 143656 84622 143712
rect 84474 139576 84530 139632
rect 85486 136720 85542 136776
rect 86774 156576 86830 156632
rect 89626 239808 89682 239864
rect 90270 239672 90326 239728
rect 91006 235728 91062 235784
rect 88338 234368 88394 234424
rect 92110 241576 92166 241632
rect 91650 240080 91706 240136
rect 92892 241440 92948 241496
rect 93122 241168 93178 241224
rect 92386 210976 92442 211032
rect 94318 240080 94374 240136
rect 94870 240080 94926 240136
rect 93766 236952 93822 237008
rect 95054 238448 95110 238504
rect 95054 238176 95110 238232
rect 95238 237224 95294 237280
rect 96434 241712 96490 241768
rect 87602 176704 87658 176760
rect 86958 167048 87014 167104
rect 86314 137264 86370 137320
rect 88982 173984 89038 174040
rect 87602 139576 87658 139632
rect 89166 143656 89222 143712
rect 89166 142704 89222 142760
rect 89626 140800 89682 140856
rect 88982 136720 89038 136776
rect 92478 171128 92534 171184
rect 91098 136040 91154 136096
rect 91282 136040 91338 136096
rect 92662 161472 92718 161528
rect 93030 144064 93086 144120
rect 94962 143928 95018 143984
rect 94134 135088 94190 135144
rect 68834 133320 68890 133376
rect 94594 124888 94650 124944
rect 67822 93336 67878 93392
rect 68006 91704 68062 91760
rect 68006 91024 68062 91080
rect 95146 138216 95202 138272
rect 69662 87488 69718 87544
rect 67822 60560 67878 60616
rect 72974 92692 72976 92712
rect 72976 92692 73028 92712
rect 73028 92692 73030 92712
rect 72974 92656 73030 92692
rect 70306 91160 70362 91216
rect 71042 91160 71098 91216
rect 71134 91024 71190 91080
rect 71686 76472 71742 76528
rect 71042 71712 71098 71768
rect 69754 70216 69810 70272
rect 70122 14456 70178 14512
rect 74262 90888 74318 90944
rect 74814 91024 74870 91080
rect 76286 92384 76342 92440
rect 78034 89800 78090 89856
rect 79506 92112 79562 92168
rect 78954 90888 79010 90944
rect 78402 85448 78458 85504
rect 82082 89392 82138 89448
rect 83002 89256 83058 89312
rect 82266 88168 82322 88224
rect 84106 88032 84162 88088
rect 82818 81368 82874 81424
rect 83462 62736 83518 62792
rect 73802 3440 73858 3496
rect 79322 15816 79378 15872
rect 82082 8880 82138 8936
rect 86130 86808 86186 86864
rect 87234 85312 87290 85368
rect 85486 17176 85542 17232
rect 88246 82048 88302 82104
rect 89258 88168 89314 88224
rect 89810 86672 89866 86728
rect 93260 92656 93316 92712
rect 91006 92384 91062 92440
rect 92386 92384 92442 92440
rect 91834 92248 91890 92304
rect 91282 89528 91338 89584
rect 94778 92384 94834 92440
rect 94686 86536 94742 86592
rect 95422 138216 95478 138272
rect 95514 127608 95570 127664
rect 95422 124072 95478 124128
rect 95330 120264 95386 120320
rect 96802 240080 96858 240136
rect 97722 241304 97778 241360
rect 97262 233416 97318 233472
rect 97722 233416 97778 233472
rect 97262 166232 97318 166288
rect 97814 166232 97870 166288
rect 96526 147076 96582 147112
rect 96526 147056 96528 147076
rect 96528 147056 96580 147076
rect 96580 147056 96582 147076
rect 96710 133864 96766 133920
rect 96710 133048 96766 133104
rect 96618 131416 96674 131472
rect 96618 130056 96674 130112
rect 96710 128424 96766 128480
rect 97170 126248 97226 126304
rect 99378 277752 99434 277808
rect 99286 271224 99342 271280
rect 98734 268368 98790 268424
rect 99194 247560 99250 247616
rect 97906 130872 97962 130928
rect 97538 129240 97594 129296
rect 97446 124616 97502 124672
rect 97354 123256 97410 123312
rect 97906 127064 97962 127120
rect 97262 122440 97318 122496
rect 97170 120808 97226 120864
rect 96066 120300 96068 120320
rect 96068 120300 96120 120320
rect 96120 120300 96122 120320
rect 96066 120264 96122 120300
rect 97262 114008 97318 114064
rect 96802 111052 96804 111072
rect 96804 111052 96856 111072
rect 96856 111052 96858 111072
rect 96802 111016 96858 111052
rect 97170 109656 97226 109712
rect 96618 96600 96674 96656
rect 97906 121624 97962 121680
rect 97814 118632 97870 118688
rect 97906 117816 97962 117872
rect 97906 117000 97962 117056
rect 97814 116456 97870 116512
rect 97906 115640 97962 115696
rect 97814 114824 97870 114880
rect 97538 113464 97594 113520
rect 97814 112648 97870 112704
rect 97906 111868 97908 111888
rect 97908 111868 97960 111888
rect 97960 111868 97962 111888
rect 97906 111832 97962 111868
rect 97446 110236 97448 110256
rect 97448 110236 97500 110256
rect 97500 110236 97502 110256
rect 97446 110200 97502 110236
rect 97906 108024 97962 108080
rect 97538 107208 97594 107264
rect 97906 106664 97962 106720
rect 97906 105848 97962 105904
rect 97538 105032 97594 105088
rect 97906 104216 97962 104272
rect 97722 103420 97778 103456
rect 97722 103400 97724 103420
rect 97724 103400 97776 103420
rect 97776 103400 97778 103420
rect 97906 102856 97962 102912
rect 97630 102040 97686 102096
rect 97906 101224 97962 101280
rect 97814 100408 97870 100464
rect 97906 99592 97962 99648
rect 97538 99084 97540 99104
rect 97540 99084 97592 99104
rect 97592 99084 97594 99104
rect 97538 99048 97594 99084
rect 97814 98232 97870 98288
rect 99470 270408 99526 270464
rect 99562 242528 99618 242584
rect 100114 284416 100170 284472
rect 100298 270444 100300 270464
rect 100300 270444 100352 270464
rect 100352 270444 100354 270464
rect 100298 270408 100354 270444
rect 100758 282648 100814 282704
rect 100758 281016 100814 281072
rect 100758 279384 100814 279440
rect 100758 276936 100814 276992
rect 100850 274488 100906 274544
rect 100758 273672 100814 273728
rect 100758 272856 100814 272912
rect 101126 272060 101182 272096
rect 101126 272040 101128 272060
rect 101128 272040 101180 272060
rect 101180 272040 101182 272060
rect 100758 268776 100814 268832
rect 101218 267960 101274 268016
rect 100758 267144 100814 267200
rect 100850 265512 100906 265568
rect 100758 263880 100814 263936
rect 100758 262268 100814 262304
rect 100758 262248 100760 262268
rect 100760 262248 100812 262268
rect 100812 262248 100814 262268
rect 101862 291896 101918 291952
rect 101494 280200 101550 280256
rect 103886 390632 103942 390688
rect 102782 387776 102838 387832
rect 101678 263064 101734 263120
rect 100942 261432 100998 261488
rect 101402 261432 101458 261488
rect 100758 260616 100814 260672
rect 100758 258984 100814 259040
rect 100758 258204 100760 258224
rect 100760 258204 100812 258224
rect 100812 258204 100814 258224
rect 100758 258168 100814 258204
rect 100390 256672 100446 256728
rect 100114 242528 100170 242584
rect 100114 241712 100170 241768
rect 100022 234504 100078 234560
rect 97906 97416 97962 97472
rect 97354 87488 97410 87544
rect 97906 95260 97962 95296
rect 97906 95240 97908 95260
rect 97908 95240 97960 95260
rect 97960 95240 97962 95260
rect 97814 94424 97870 94480
rect 98734 92248 98790 92304
rect 100758 257388 100760 257408
rect 100760 257388 100812 257408
rect 100812 257388 100814 257408
rect 100758 257352 100814 257388
rect 100850 254904 100906 254960
rect 100758 254088 100814 254144
rect 100758 253272 100814 253328
rect 100850 252456 100906 252512
rect 100758 250824 100814 250880
rect 101218 259836 101220 259856
rect 101220 259836 101272 259856
rect 101272 259836 101274 259856
rect 101218 259800 101274 259836
rect 101034 255720 101090 255776
rect 101954 250008 102010 250064
rect 101678 248376 101734 248432
rect 101034 246744 101090 246800
rect 101126 245928 101182 245984
rect 101034 242664 101090 242720
rect 103426 318280 103482 318336
rect 102782 284144 102838 284200
rect 102230 276120 102286 276176
rect 102782 268504 102838 268560
rect 105266 389000 105322 389056
rect 102414 245656 102470 245712
rect 102322 245112 102378 245168
rect 102230 243480 102286 243536
rect 102414 244296 102470 244352
rect 102230 234504 102286 234560
rect 103426 245656 103482 245712
rect 103426 241576 103482 241632
rect 103426 241304 103482 241360
rect 102782 162832 102838 162888
rect 100114 102176 100170 102232
rect 99010 96056 99066 96112
rect 99010 92384 99066 92440
rect 98826 80008 98882 80064
rect 99286 80008 99342 80064
rect 100758 91044 100814 91080
rect 100758 91024 100760 91044
rect 100760 91024 100812 91044
rect 100812 91024 100814 91044
rect 103426 159296 103482 159352
rect 103426 156576 103482 156632
rect 102874 139440 102930 139496
rect 101494 75792 101550 75848
rect 97262 72936 97318 72992
rect 90362 61376 90418 61432
rect 95146 55800 95202 55856
rect 99286 66816 99342 66872
rect 101034 3304 101090 3360
rect 103702 291216 103758 291272
rect 103610 237088 103666 237144
rect 105818 284144 105874 284200
rect 106186 271088 106242 271144
rect 106186 251640 106242 251696
rect 105634 234368 105690 234424
rect 105634 206352 105690 206408
rect 104990 205672 105046 205728
rect 105634 205672 105690 205728
rect 104806 203496 104862 203552
rect 104162 138080 104218 138136
rect 103610 86808 103666 86864
rect 104714 86808 104770 86864
rect 104714 86536 104770 86592
rect 105082 142160 105138 142216
rect 104990 124208 105046 124264
rect 107750 390496 107806 390552
rect 107658 390224 107714 390280
rect 107750 389136 107806 389192
rect 106646 254532 106648 254552
rect 106648 254532 106700 254552
rect 106700 254532 106702 254552
rect 106646 254496 106702 254532
rect 107014 292576 107070 292632
rect 107474 251232 107530 251288
rect 107474 241848 107530 241904
rect 106370 238448 106426 238504
rect 106922 213152 106978 213208
rect 108946 236544 109002 236600
rect 108302 229744 108358 229800
rect 108486 154536 108542 154592
rect 111706 390360 111762 390416
rect 110510 288496 110566 288552
rect 109130 90888 109186 90944
rect 108394 90344 108450 90400
rect 113362 424904 113418 424960
rect 113822 430072 113878 430128
rect 113454 416744 113510 416800
rect 110694 242528 110750 242584
rect 114650 437416 114706 437472
rect 114650 424088 114706 424144
rect 114558 421912 114614 421968
rect 114650 418920 114706 418976
rect 115570 432248 115626 432304
rect 115846 431160 115902 431216
rect 115754 429256 115810 429312
rect 115846 428168 115902 428224
rect 115846 425992 115902 426048
rect 115754 424904 115810 424960
rect 115846 424088 115902 424144
rect 115846 423000 115902 423056
rect 115754 420824 115810 420880
rect 115846 416780 115848 416800
rect 115848 416780 115900 416800
rect 115900 416780 115902 416800
rect 115846 416744 115902 416780
rect 115846 415692 115848 415712
rect 115848 415692 115900 415712
rect 115900 415692 115902 415712
rect 115846 415656 115902 415692
rect 115846 414860 115902 414896
rect 115846 414840 115848 414860
rect 115848 414840 115900 414860
rect 115900 414840 115902 414860
rect 115846 413752 115902 413808
rect 115110 412664 115166 412720
rect 115202 411576 115258 411632
rect 115846 410488 115902 410544
rect 115846 409672 115902 409728
rect 115018 407516 115074 407552
rect 115018 407496 115020 407516
rect 115020 407496 115072 407516
rect 115072 407496 115074 407516
rect 115846 405628 115848 405648
rect 115848 405628 115900 405648
rect 115900 405628 115902 405648
rect 115846 405592 115902 405628
rect 115846 404540 115848 404560
rect 115848 404540 115900 404560
rect 115900 404540 115902 404560
rect 115846 404504 115902 404540
rect 115846 403416 115902 403472
rect 114558 399472 114614 399528
rect 114558 398792 114614 398848
rect 114558 396344 114614 396400
rect 114558 391992 114614 392048
rect 111614 216008 111670 216064
rect 110418 85448 110474 85504
rect 109314 3440 109370 3496
rect 113178 287136 113234 287192
rect 112626 245656 112682 245712
rect 112442 220224 112498 220280
rect 111798 89392 111854 89448
rect 114098 294616 114154 294672
rect 115846 402328 115902 402384
rect 115202 401240 115258 401296
rect 115018 391196 115074 391232
rect 115018 391176 115020 391196
rect 115020 391176 115072 391196
rect 115072 391176 115074 391196
rect 115846 400424 115902 400480
rect 115386 399336 115442 399392
rect 115570 398248 115626 398304
rect 115846 397160 115902 397216
rect 115846 395256 115902 395312
rect 115386 394168 115442 394224
rect 115202 335416 115258 335472
rect 115846 393080 115902 393136
rect 116582 536696 116638 536752
rect 117318 384240 117374 384296
rect 116582 318280 116638 318336
rect 116030 318144 116086 318200
rect 115294 243480 115350 243536
rect 115202 241576 115258 241632
rect 115386 238584 115442 238640
rect 115202 228928 115258 228984
rect 115754 224984 115810 225040
rect 113178 153720 113234 153776
rect 113270 88032 113326 88088
rect 115846 220088 115902 220144
rect 115202 150456 115258 150512
rect 115754 150456 115810 150512
rect 117226 249056 117282 249112
rect 117226 214512 117282 214568
rect 116674 153176 116730 153232
rect 116582 146920 116638 146976
rect 117962 302504 118018 302560
rect 119986 312160 120042 312216
rect 118698 233180 118700 233200
rect 118700 233180 118752 233200
rect 118752 233180 118754 233200
rect 118698 233144 118754 233180
rect 118790 226208 118846 226264
rect 118790 224984 118846 225040
rect 117962 167184 118018 167240
rect 117962 144064 118018 144120
rect 118606 144064 118662 144120
rect 119342 86672 119398 86728
rect 121458 312024 121514 312080
rect 122102 318280 122158 318336
rect 120722 220224 120778 220280
rect 122102 88168 122158 88224
rect 122654 88168 122710 88224
rect 120170 88032 120226 88088
rect 132590 582664 132646 582720
rect 124770 389036 124772 389056
rect 124772 389036 124824 389056
rect 124824 389036 124826 389056
rect 124770 389000 124826 389036
rect 125414 316684 125416 316704
rect 125416 316684 125468 316704
rect 125468 316684 125470 316704
rect 125414 316648 125470 316684
rect 124218 307808 124274 307864
rect 122930 243480 122986 243536
rect 122838 235864 122894 235920
rect 122838 85312 122894 85368
rect 124034 85312 124090 85368
rect 126242 275984 126298 276040
rect 125598 92520 125654 92576
rect 126334 249056 126390 249112
rect 127714 282920 127770 282976
rect 128450 262792 128506 262848
rect 127714 149096 127770 149152
rect 129738 258712 129794 258768
rect 128542 239808 128598 239864
rect 129002 229880 129058 229936
rect 131118 286320 131174 286376
rect 131854 261432 131910 261488
rect 131762 118904 131818 118960
rect 133234 299512 133290 299568
rect 133970 281560 134026 281616
rect 135902 288496 135958 288552
rect 134614 284280 134670 284336
rect 134522 280744 134578 280800
rect 137282 307944 137338 308000
rect 136638 267008 136694 267064
rect 137466 289856 137522 289912
rect 138662 281560 138718 281616
rect 138018 257216 138074 257272
rect 140778 398792 140834 398848
rect 140134 304136 140190 304192
rect 140870 277344 140926 277400
rect 140870 276664 140926 276720
rect 141054 253136 141110 253192
rect 140134 228928 140190 228984
rect 142802 320184 142858 320240
rect 143538 269728 143594 269784
rect 145654 284824 145710 284880
rect 144918 274488 144974 274544
rect 142986 157392 143042 157448
rect 144274 242120 144330 242176
rect 144826 202136 144882 202192
rect 146206 274488 146262 274544
rect 146206 273808 146262 273864
rect 146298 255856 146354 255912
rect 146298 255312 146354 255368
rect 145654 160112 145710 160168
rect 147678 260752 147734 260808
rect 147678 260072 147734 260128
rect 149794 288496 149850 288552
rect 149702 193840 149758 193896
rect 148414 152360 148470 152416
rect 151174 304952 151230 305008
rect 151174 165688 151230 165744
rect 148322 3440 148378 3496
rect 155222 308080 155278 308136
rect 153934 267008 153990 267064
rect 153198 223488 153254 223544
rect 153842 161744 153898 161800
rect 154210 157392 154266 157448
rect 153842 131144 153898 131200
rect 159362 303864 159418 303920
rect 155406 276664 155462 276720
rect 155314 262792 155370 262848
rect 155406 249056 155462 249112
rect 158074 284824 158130 284880
rect 156694 238448 156750 238504
rect 157246 237904 157302 237960
rect 157246 230424 157302 230480
rect 156602 84088 156658 84144
rect 160098 298696 160154 298752
rect 160742 286320 160798 286376
rect 159454 237088 159510 237144
rect 159914 237088 159970 237144
rect 159454 108976 159510 109032
rect 160006 108976 160062 109032
rect 160926 235320 160982 235376
rect 162214 269728 162270 269784
rect 160742 143520 160798 143576
rect 160834 84088 160890 84144
rect 162122 241576 162178 241632
rect 162214 232600 162270 232656
rect 162122 226072 162178 226128
rect 162122 224984 162178 225040
rect 162766 224984 162822 225040
rect 161570 144880 161626 144936
rect 162122 144880 162178 144936
rect 162122 117136 162178 117192
rect 166170 92384 166226 92440
rect 169298 255856 169354 255912
rect 169114 149640 169170 149696
rect 169298 149096 169354 149152
rect 167826 138624 167882 138680
rect 173254 293120 173310 293176
rect 172426 287680 172482 287736
rect 170586 273808 170642 273864
rect 170586 233280 170642 233336
rect 171874 226344 171930 226400
rect 172334 114552 172390 114608
rect 177302 305088 177358 305144
rect 176014 268368 176070 268424
rect 173346 260072 173402 260128
rect 173346 247560 173402 247616
rect 173254 158752 173310 158808
rect 173806 141480 173862 141536
rect 174634 251232 174690 251288
rect 175186 217368 175242 217424
rect 175186 216688 175242 216744
rect 175830 147056 175886 147112
rect 174542 76472 174598 76528
rect 178038 282940 178094 282976
rect 178038 282920 178040 282940
rect 178040 282920 178092 282940
rect 178092 282920 178094 282940
rect 177302 280744 177358 280800
rect 176566 240760 176622 240816
rect 176566 92384 176622 92440
rect 178682 238584 178738 238640
rect 178682 147736 178738 147792
rect 178774 145560 178830 145616
rect 180154 305224 180210 305280
rect 179418 235456 179474 235512
rect 182822 303728 182878 303784
rect 180246 262792 180302 262848
rect 180154 235592 180210 235648
rect 180338 257216 180394 257272
rect 180338 233960 180394 234016
rect 180154 178608 180210 178664
rect 180154 117952 180210 118008
rect 180706 81368 180762 81424
rect 181534 213968 181590 214024
rect 181534 209616 181590 209672
rect 182086 209616 182142 209672
rect 182178 144744 182234 144800
rect 182178 135904 182234 135960
rect 182086 109112 182142 109168
rect 182914 261432 182970 261488
rect 187054 309440 187110 309496
rect 186962 296656 187018 296712
rect 185766 258712 185822 258768
rect 184202 233824 184258 233880
rect 182914 219272 182970 219328
rect 182914 218048 182970 218104
rect 183466 218048 183522 218104
rect 184478 161608 184534 161664
rect 184202 149640 184258 149696
rect 183466 144744 183522 144800
rect 183466 143520 183522 143576
rect 184294 147192 184350 147248
rect 184478 145696 184534 145752
rect 184294 124208 184350 124264
rect 182822 82048 182878 82104
rect 184294 85312 184350 85368
rect 184202 82592 184258 82648
rect 184754 74432 184810 74488
rect 189722 309304 189778 309360
rect 188342 306584 188398 306640
rect 186226 227568 186282 227624
rect 186134 222944 186190 223000
rect 186134 222264 186190 222320
rect 186134 108160 186190 108216
rect 185582 77832 185638 77888
rect 187054 249056 187110 249112
rect 188710 301280 188766 301336
rect 188526 301144 188582 301200
rect 188434 291080 188490 291136
rect 188342 241576 188398 241632
rect 187238 232464 187294 232520
rect 187054 156032 187110 156088
rect 186962 148280 187018 148336
rect 186226 89528 186282 89584
rect 187146 150456 187202 150512
rect 189906 302368 189962 302424
rect 190458 300872 190514 300928
rect 191102 310800 191158 310856
rect 190550 299784 190606 299840
rect 191102 300600 191158 300656
rect 191286 298560 191342 298616
rect 191194 297472 191250 297528
rect 190366 297336 190422 297392
rect 190458 296248 190514 296304
rect 189906 294480 189962 294536
rect 190550 293936 190606 293992
rect 191102 291624 191158 291680
rect 189722 289720 189778 289776
rect 191010 289312 191066 289368
rect 191010 283600 191066 283656
rect 190458 280064 190514 280120
rect 190366 278976 190422 279032
rect 189722 270544 189778 270600
rect 188986 160656 189042 160712
rect 188434 159296 188490 159352
rect 188066 153720 188122 153776
rect 188342 150728 188398 150784
rect 188066 145832 188122 145888
rect 187698 139440 187754 139496
rect 187698 135088 187754 135144
rect 188894 145560 188950 145616
rect 188434 144200 188490 144256
rect 189814 244568 189870 244624
rect 189906 242936 189962 242992
rect 189906 235184 189962 235240
rect 191010 266328 191066 266384
rect 190642 255856 190698 255912
rect 190826 251268 190828 251288
rect 190828 251268 190880 251288
rect 190880 251268 190882 251288
rect 190826 251232 190882 251268
rect 190642 246608 190698 246664
rect 190366 232464 190422 232520
rect 189814 221448 189870 221504
rect 189722 156576 189778 156632
rect 189722 151816 189778 151872
rect 189078 142296 189134 142352
rect 188986 139440 189042 139496
rect 189722 138488 189778 138544
rect 189906 148552 189962 148608
rect 189814 133864 189870 133920
rect 190366 133728 190422 133784
rect 190366 132504 190422 132560
rect 201498 328480 201554 328536
rect 196990 306720 197046 306776
rect 192482 296520 192538 296576
rect 195978 302776 196034 302832
rect 200210 302368 200266 302424
rect 198278 302232 198334 302288
rect 203614 311888 203670 311944
rect 201774 309168 201830 309224
rect 202510 308216 202566 308272
rect 203430 304952 203486 305008
rect 204902 310664 204958 310720
rect 204258 310528 204314 310584
rect 208398 309440 208454 309496
rect 207846 301824 207902 301880
rect 209778 306584 209834 306640
rect 220910 313384 220966 313440
rect 219990 308080 220046 308136
rect 218058 307944 218114 308000
rect 214838 305224 214894 305280
rect 213918 303628 213920 303648
rect 213920 303628 213972 303648
rect 213972 303628 213974 303648
rect 213918 303592 213974 303628
rect 215482 305088 215538 305144
rect 215298 303864 215354 303920
rect 224038 314744 224094 314800
rect 226982 303592 227038 303648
rect 232502 318824 232558 318880
rect 240138 312160 240194 312216
rect 234618 303728 234674 303784
rect 240046 303628 240048 303648
rect 240048 303628 240100 303648
rect 240100 303628 240102 303648
rect 240046 303592 240102 303628
rect 240690 303612 240746 303648
rect 240690 303592 240692 303612
rect 240692 303592 240744 303612
rect 240744 303592 240746 303612
rect 242990 303592 243046 303648
rect 198738 301416 198794 301472
rect 224774 301280 224830 301336
rect 233790 301280 233846 301336
rect 235630 301280 235686 301336
rect 236918 301280 236974 301336
rect 239494 301280 239550 301336
rect 194230 301144 194286 301200
rect 200578 301144 200634 301200
rect 218426 301008 218482 301064
rect 194690 300872 194746 300928
rect 197358 300872 197414 300928
rect 199290 300872 199346 300928
rect 205638 300872 205694 300928
rect 206282 300872 206338 300928
rect 207110 300872 207166 300928
rect 211526 300872 211582 300928
rect 217046 300872 217102 300928
rect 218978 300872 219034 300928
rect 219438 300908 219440 300928
rect 219440 300908 219492 300928
rect 219492 300908 219494 300928
rect 219438 300872 219494 300908
rect 221646 300872 221702 300928
rect 222382 300872 222438 300928
rect 224130 300872 224186 300928
rect 225970 300872 226026 300928
rect 226522 300872 226578 300928
rect 227258 300872 227314 300928
rect 229834 300872 229890 300928
rect 230570 300872 230626 300928
rect 231214 300872 231270 300928
rect 232042 300872 232098 300928
rect 232502 300872 232558 300928
rect 233330 300872 233386 300928
rect 234986 300872 235042 300928
rect 236642 300872 236698 300928
rect 238850 300872 238906 300928
rect 241426 300872 241482 300928
rect 241978 300872 242034 300928
rect 243266 300872 243322 300928
rect 244922 306992 244978 307048
rect 246118 304000 246174 304056
rect 247682 302776 247738 302832
rect 248510 302504 248566 302560
rect 244554 301008 244610 301064
rect 249154 316648 249210 316704
rect 249154 304136 249210 304192
rect 249338 303864 249394 303920
rect 249982 303592 250038 303648
rect 254030 312024 254086 312080
rect 251914 302232 251970 302288
rect 251822 301688 251878 301744
rect 245106 300872 245162 300928
rect 246394 300872 246450 300928
rect 247774 300872 247830 300928
rect 248510 300872 248566 300928
rect 251546 300872 251602 300928
rect 252466 300872 252522 300928
rect 252926 300600 252982 300656
rect 191378 293120 191434 293176
rect 193126 292848 193182 292904
rect 191746 288224 191802 288280
rect 191286 287680 191342 287736
rect 191654 285912 191710 285968
rect 191194 284824 191250 284880
rect 191562 284688 191618 284744
rect 192390 282376 192446 282432
rect 193034 282376 193090 282432
rect 191746 281288 191802 281344
rect 191654 277752 191710 277808
rect 191654 274352 191710 274408
rect 191562 273128 191618 273184
rect 191654 272040 191710 272096
rect 191654 269728 191710 269784
rect 191654 268640 191710 268696
rect 191286 267416 191342 267472
rect 191562 265104 191618 265160
rect 191654 262792 191710 262848
rect 191654 261704 191710 261760
rect 191286 260480 191342 260536
rect 191654 257080 191710 257136
rect 191654 254768 191710 254824
rect 191654 253544 191710 253600
rect 191654 252456 191710 252512
rect 191654 250144 191710 250200
rect 191654 248920 191710 248976
rect 191654 247832 191710 247888
rect 191562 148416 191618 148472
rect 191654 148280 191710 148336
rect 191562 138216 191618 138272
rect 191562 136312 191618 136368
rect 191562 135496 191618 135552
rect 190366 129784 190422 129840
rect 190642 122984 190698 123040
rect 191102 120264 191158 120320
rect 190366 120128 190422 120184
rect 188986 117408 189042 117464
rect 191102 118632 191158 118688
rect 190366 117136 190422 117192
rect 190642 116728 190698 116784
rect 187146 78512 187202 78568
rect 190366 113464 190422 113520
rect 191010 113212 191066 113248
rect 191010 113192 191012 113212
rect 191012 113192 191064 113212
rect 191064 113192 191066 113212
rect 190366 110744 190422 110800
rect 190366 108976 190422 109032
rect 188342 73072 188398 73128
rect 190458 105032 190514 105088
rect 189078 82728 189134 82784
rect 189078 81504 189134 81560
rect 189722 81504 189778 81560
rect 191010 103400 191066 103456
rect 190642 101496 190698 101552
rect 190642 99864 190698 99920
rect 190826 98776 190882 98832
rect 191654 131960 191710 132016
rect 191654 129240 191710 129296
rect 191654 126520 191710 126576
rect 191654 123800 191710 123856
rect 191654 122168 191710 122224
rect 191562 121352 191618 121408
rect 191562 120128 191618 120184
rect 191654 119448 191710 119504
rect 191194 117408 191250 117464
rect 191654 115912 191710 115968
rect 192482 228792 192538 228848
rect 191838 211112 191894 211168
rect 193218 290536 193274 290592
rect 253478 301008 253534 301064
rect 253938 296384 253994 296440
rect 253938 293800 253994 293856
rect 253018 290128 253074 290184
rect 252926 289720 252982 289776
rect 252834 281288 252890 281344
rect 252834 274760 252890 274816
rect 252926 267280 252982 267336
rect 193402 258848 193458 258904
rect 193586 242800 193642 242856
rect 195978 241440 196034 241496
rect 195242 237904 195298 237960
rect 195242 235456 195298 235512
rect 193770 224304 193826 224360
rect 193862 181328 193918 181384
rect 192850 137400 192906 137456
rect 192482 127608 192538 127664
rect 191562 109656 191618 109712
rect 191562 106936 191618 106992
rect 191746 112412 191748 112432
rect 191748 112412 191800 112432
rect 191800 112412 191802 112432
rect 191746 112376 191802 112412
rect 191746 110492 191802 110528
rect 191746 110472 191748 110492
rect 191748 110472 191800 110492
rect 191800 110472 191802 110492
rect 191746 107788 191748 107808
rect 191748 107788 191800 107808
rect 191800 107788 191802 107808
rect 191746 107752 191802 107788
rect 191746 106120 191802 106176
rect 191654 104216 191710 104272
rect 191654 100680 191710 100736
rect 191746 97960 191802 98016
rect 191562 96328 191618 96384
rect 191654 94424 191710 94480
rect 191838 92112 191894 92168
rect 193402 160792 193458 160848
rect 193126 144064 193182 144120
rect 193034 134680 193090 134736
rect 193402 139576 193458 139632
rect 193126 128424 193182 128480
rect 192942 127608 192998 127664
rect 192850 83408 192906 83464
rect 193034 92248 193090 92304
rect 193034 91160 193090 91216
rect 194690 143384 194746 143440
rect 194690 142160 194746 142216
rect 198646 240216 198702 240272
rect 196622 235184 196678 235240
rect 196622 221448 196678 221504
rect 198002 175344 198058 175400
rect 196622 164872 196678 164928
rect 196070 159296 196126 159352
rect 196898 159296 196954 159352
rect 196714 147192 196770 147248
rect 196530 145696 196586 145752
rect 195242 143384 195298 143440
rect 195978 142160 196034 142216
rect 197082 142296 197138 142352
rect 196898 142160 196954 142216
rect 197910 148552 197966 148608
rect 198094 154672 198150 154728
rect 198646 154672 198702 154728
rect 198094 149640 198150 149696
rect 203982 236544 204038 236600
rect 202786 223488 202842 223544
rect 200762 208392 200818 208448
rect 201498 168408 201554 168464
rect 202142 168408 202198 168464
rect 201406 145696 201462 145752
rect 200210 144200 200266 144256
rect 198830 143656 198886 143712
rect 198002 143384 198058 143440
rect 198922 143384 198978 143440
rect 198646 141072 198702 141128
rect 201314 143520 201370 143576
rect 201406 142160 201462 142216
rect 205546 235864 205602 235920
rect 205454 171672 205510 171728
rect 203522 140392 203578 140448
rect 204442 145832 204498 145888
rect 205086 156168 205142 156224
rect 204902 143520 204958 143576
rect 205638 169768 205694 169824
rect 205546 156168 205602 156224
rect 207110 233824 207166 233880
rect 206374 173848 206430 173904
rect 205638 144064 205694 144120
rect 205546 143520 205602 143576
rect 204994 141344 205050 141400
rect 205454 141344 205510 141400
rect 205086 140936 205142 140992
rect 208490 228792 208546 228848
rect 208490 227704 208546 227760
rect 211066 233144 211122 233200
rect 212078 227024 212134 227080
rect 213182 206216 213238 206272
rect 213182 177248 213238 177304
rect 208398 150320 208454 150376
rect 210238 148416 210294 148472
rect 210054 146920 210110 146976
rect 215942 240896 215998 240952
rect 215390 240080 215446 240136
rect 213458 142704 213514 142760
rect 213458 142160 213514 142216
rect 214562 173984 214618 174040
rect 215482 167048 215538 167104
rect 214746 141072 214802 141128
rect 216034 167048 216090 167104
rect 215942 152360 215998 152416
rect 216678 157392 216734 157448
rect 222382 240080 222438 240136
rect 223486 240080 223542 240136
rect 221002 233960 221058 234016
rect 217414 157392 217470 157448
rect 218794 141344 218850 141400
rect 218886 140800 218942 140856
rect 219530 142704 219586 142760
rect 222106 238584 222162 238640
rect 222198 172352 222254 172408
rect 222198 171128 222254 171184
rect 221002 142704 221058 142760
rect 222290 162696 222346 162752
rect 222290 161472 222346 161528
rect 222842 238040 222898 238096
rect 223578 226480 223634 226536
rect 223578 224168 223634 224224
rect 222934 172352 222990 172408
rect 224958 207032 225014 207088
rect 224866 173168 224922 173224
rect 223578 167184 223634 167240
rect 224222 167184 224278 167240
rect 222842 162696 222898 162752
rect 222934 156168 222990 156224
rect 222382 148416 222438 148472
rect 222934 142024 222990 142080
rect 225326 141344 225382 141400
rect 226338 137128 226394 137184
rect 225326 135496 225382 135552
rect 226338 126520 226394 126576
rect 225142 123800 225198 123856
rect 226338 122168 226394 122224
rect 225050 118088 225106 118144
rect 226338 117544 226394 117600
rect 225142 116728 225198 116784
rect 193402 100680 193458 100736
rect 225326 111288 225382 111344
rect 226338 105848 226394 105904
rect 226246 102720 226302 102776
rect 225234 102312 225290 102368
rect 226246 100680 226302 100736
rect 216126 93336 216182 93392
rect 201406 92928 201462 92984
rect 193862 92792 193918 92848
rect 195518 92792 195574 92848
rect 194690 71712 194746 71768
rect 194690 70352 194746 70408
rect 195242 70352 195298 70408
rect 194598 70216 194654 70272
rect 194598 69808 194654 69864
rect 195334 69808 195390 69864
rect 195334 64096 195390 64152
rect 196530 92384 196586 92440
rect 198002 91976 198058 92032
rect 198370 89664 198426 89720
rect 200486 92792 200542 92848
rect 200762 91840 200818 91896
rect 201590 92792 201646 92848
rect 203522 92248 203578 92304
rect 204166 92420 204168 92440
rect 204168 92420 204220 92440
rect 204220 92420 204222 92440
rect 204166 92384 204222 92420
rect 203614 90344 203670 90400
rect 204626 92656 204682 92712
rect 204442 89800 204498 89856
rect 205086 92656 205142 92712
rect 205086 90888 205142 90944
rect 204994 85448 205050 85504
rect 207110 92792 207166 92848
rect 207386 90208 207442 90264
rect 208306 90208 208362 90264
rect 204626 60560 204682 60616
rect 204626 60152 204682 60208
rect 204994 60152 205050 60208
rect 208398 86808 208454 86864
rect 208766 92792 208822 92848
rect 209870 81368 209926 81424
rect 210054 92792 210110 92848
rect 210330 89256 210386 89312
rect 211066 81368 211122 81424
rect 209962 77152 210018 77208
rect 213642 92792 213698 92848
rect 214010 86536 214066 86592
rect 212538 81368 212594 81424
rect 212538 80144 212594 80200
rect 213182 80144 213238 80200
rect 224498 93336 224554 93392
rect 217690 88032 217746 88088
rect 218242 86672 218298 86728
rect 219898 90344 219954 90400
rect 220082 89528 220138 89584
rect 221922 88168 221978 88224
rect 223578 92384 223634 92440
rect 223762 91024 223818 91080
rect 224866 91024 224922 91080
rect 224222 72936 224278 72992
rect 225142 97960 225198 98016
rect 226154 97960 226210 98016
rect 225050 84088 225106 84144
rect 226522 134680 226578 134736
rect 227718 239672 227774 239728
rect 228362 239672 228418 239728
rect 226706 134680 226762 134736
rect 226706 133592 226762 133648
rect 227074 132776 227130 132832
rect 226706 131960 226762 132016
rect 226706 130872 226762 130928
rect 226706 129240 226762 129296
rect 226706 128424 226762 128480
rect 226614 127336 226670 127392
rect 226706 125704 226762 125760
rect 226706 124616 226762 124672
rect 226706 122984 226762 123040
rect 226706 120264 226762 120320
rect 226522 119448 226578 119504
rect 226614 118360 226670 118416
rect 226706 115912 226762 115968
rect 226522 114824 226578 114880
rect 227350 114008 227406 114064
rect 226522 110472 226578 110528
rect 226614 108568 226670 108624
rect 226706 107752 226762 107808
rect 226706 106936 226762 106992
rect 226614 105032 226670 105088
rect 226522 104216 226578 104272
rect 226430 96056 226486 96112
rect 226614 103400 226670 103456
rect 226706 101496 226762 101552
rect 226614 97144 226670 97200
rect 226614 95240 226670 95296
rect 226706 94424 226762 94480
rect 227534 99592 227590 99648
rect 226982 93608 227038 93664
rect 227810 234368 227866 234424
rect 231122 239400 231178 239456
rect 227810 164192 227866 164248
rect 232502 213424 232558 213480
rect 230478 211112 230534 211168
rect 231122 211112 231178 211168
rect 229190 162696 229246 162752
rect 229742 162696 229798 162752
rect 229190 161472 229246 161528
rect 229098 152360 229154 152416
rect 229282 150592 229338 150648
rect 229190 138624 229246 138680
rect 227810 113192 227866 113248
rect 227810 109656 227866 109712
rect 227902 102312 227958 102368
rect 229742 93064 229798 93120
rect 231950 160112 232006 160168
rect 231858 159296 231914 159352
rect 231858 156032 231914 156088
rect 234710 240080 234766 240136
rect 233238 235184 233294 235240
rect 232594 160112 232650 160168
rect 232502 156032 232558 156088
rect 234618 232620 234674 232656
rect 234618 232600 234620 232620
rect 234620 232600 234672 232620
rect 234672 232600 234674 232620
rect 235998 240080 236054 240136
rect 234710 229744 234766 229800
rect 234618 153176 234674 153232
rect 233238 149096 233294 149152
rect 231950 139984 232006 140040
rect 231950 135904 232006 135960
rect 230478 90344 230534 90400
rect 229190 75792 229246 75848
rect 231950 82592 232006 82648
rect 233238 78512 233294 78568
rect 238850 238720 238906 238776
rect 238758 165688 238814 165744
rect 238022 140936 238078 140992
rect 235998 66816 236054 66872
rect 238114 111852 238170 111888
rect 238114 111832 238116 111852
rect 238116 111832 238168 111852
rect 238168 111832 238170 111852
rect 240690 111832 240746 111888
rect 241518 237904 241574 237960
rect 245014 239536 245070 239592
rect 244278 221584 244334 221640
rect 241334 92248 241390 92304
rect 152462 3304 152518 3360
rect 214562 3304 214618 3360
rect 249706 211112 249762 211168
rect 249154 143520 249210 143576
rect 249062 102720 249118 102776
rect 249798 91976 249854 92032
rect 246302 81368 246358 81424
rect 246394 3304 246450 3360
rect 251822 241576 251878 241632
rect 251178 227704 251234 227760
rect 251914 240080 251970 240136
rect 251914 228928 251970 228984
rect 251914 227704 251970 227760
rect 252466 224304 252522 224360
rect 252926 242800 252982 242856
rect 253018 242392 253074 242448
rect 254122 291080 254178 291136
rect 255318 302232 255374 302288
rect 255410 299920 255466 299976
rect 255134 298968 255190 299024
rect 254214 287544 254270 287600
rect 256054 321544 256110 321600
rect 255502 297200 255558 297256
rect 255594 296812 255650 296848
rect 255594 296792 255596 296812
rect 255596 296792 255648 296812
rect 255648 296792 255650 296812
rect 255686 295976 255742 296032
rect 255502 295432 255558 295488
rect 255594 295024 255650 295080
rect 255502 294616 255558 294672
rect 255594 293256 255650 293312
rect 255502 292848 255558 292904
rect 255502 292440 255558 292496
rect 255962 294208 256018 294264
rect 255594 291488 255650 291544
rect 255502 290264 255558 290320
rect 255594 289040 255650 289096
rect 255502 288904 255558 288960
rect 255502 288088 255558 288144
rect 255502 287136 255558 287192
rect 255410 286728 255466 286784
rect 255594 286320 255650 286376
rect 255502 285368 255558 285424
rect 255318 284960 255374 285016
rect 255410 284552 255466 284608
rect 255594 284144 255650 284200
rect 255410 283192 255466 283248
rect 255410 282376 255466 282432
rect 255502 281968 255558 282024
rect 255410 281460 255412 281480
rect 255412 281460 255464 281480
rect 255464 281460 255466 281480
rect 255410 281424 255466 281460
rect 255410 280220 255466 280256
rect 255410 280200 255412 280220
rect 255412 280200 255464 280220
rect 255464 280200 255466 280220
rect 255318 279248 255374 279304
rect 254030 278432 254086 278488
rect 255502 278024 255558 278080
rect 255410 277500 255466 277536
rect 255410 277480 255412 277500
rect 255412 277480 255464 277500
rect 255464 277480 255466 277500
rect 255410 277108 255412 277128
rect 255412 277108 255464 277128
rect 255464 277108 255466 277128
rect 255410 277072 255466 277108
rect 255502 276256 255558 276312
rect 255410 275848 255466 275904
rect 255410 275304 255466 275360
rect 255318 274524 255320 274544
rect 255320 274524 255372 274544
rect 255372 274524 255374 274544
rect 255318 274488 255374 274524
rect 255502 274080 255558 274136
rect 255410 273164 255412 273184
rect 255412 273164 255464 273184
rect 255464 273164 255466 273184
rect 255410 273128 255466 273164
rect 256054 284960 256110 285016
rect 255502 270136 255558 270192
rect 255410 269728 255466 269784
rect 255318 268776 255374 268832
rect 255410 268368 255466 268424
rect 255502 267008 255558 267064
rect 255410 266600 255466 266656
rect 254030 266192 254086 266248
rect 255318 265784 255374 265840
rect 255502 264832 255558 264888
rect 255318 264424 255374 264480
rect 256606 283736 256662 283792
rect 258078 307808 258134 307864
rect 256882 303592 256938 303648
rect 256790 288496 256846 288552
rect 256974 292712 257030 292768
rect 256606 280064 256662 280120
rect 256606 271904 256662 271960
rect 258262 302776 258318 302832
rect 258170 282784 258226 282840
rect 256606 271360 256662 271416
rect 256054 264016 256110 264072
rect 255410 263084 255466 263120
rect 255410 263064 255412 263084
rect 255412 263064 255464 263084
rect 255464 263064 255466 263084
rect 255410 262268 255466 262304
rect 255410 262248 255412 262268
rect 255412 262248 255464 262268
rect 255464 262248 255466 262268
rect 255502 261840 255558 261896
rect 255318 261296 255374 261352
rect 255410 260888 255466 260944
rect 255410 259528 255466 259584
rect 255502 259120 255558 259176
rect 255502 257896 255558 257952
rect 255318 256944 255374 257000
rect 255502 256536 255558 256592
rect 255410 256128 255466 256184
rect 255502 255176 255558 255232
rect 255594 254360 255650 254416
rect 255410 253952 255466 254008
rect 255410 252592 255466 252648
rect 255594 252184 255650 252240
rect 255410 251776 255466 251832
rect 255502 250824 255558 250880
rect 255410 250008 255466 250064
rect 255318 249464 255374 249520
rect 255410 249056 255466 249112
rect 255594 248376 255650 248432
rect 255410 248240 255466 248296
rect 255318 247832 255374 247888
rect 254766 245520 254822 245576
rect 254122 243344 254178 243400
rect 254582 238040 254638 238096
rect 255410 246880 255466 246936
rect 255686 246472 255742 246528
rect 255502 245112 255558 245168
rect 255410 244316 255466 244352
rect 255410 244296 255412 244316
rect 255412 244296 255464 244316
rect 255464 244296 255466 244316
rect 256146 253000 256202 253056
rect 256054 250416 256110 250472
rect 256238 251232 256294 251288
rect 256422 248648 256478 248704
rect 256146 247016 256202 247072
rect 256054 237904 256110 237960
rect 258078 270952 258134 271008
rect 256790 246064 256846 246120
rect 256054 235456 256110 235512
rect 256054 222944 256110 223000
rect 256146 217368 256202 217424
rect 250442 77152 250498 77208
rect 252558 166232 252614 166288
rect 254582 91024 254638 91080
rect 256974 238720 257030 238776
rect 256882 233824 256938 233880
rect 256790 211112 256846 211168
rect 258262 247288 258318 247344
rect 258354 240896 258410 240952
rect 257342 142160 257398 142216
rect 258722 202816 258778 202872
rect 259642 280608 259698 280664
rect 259826 284960 259882 285016
rect 259734 269184 259790 269240
rect 259734 235320 259790 235376
rect 260838 270816 260894 270872
rect 259458 150456 259514 150512
rect 261114 278840 261170 278896
rect 261206 272176 261262 272232
rect 261114 262656 261170 262712
rect 261022 237088 261078 237144
rect 261114 234504 261170 234560
rect 262494 306448 262550 306504
rect 262402 285640 262458 285696
rect 267646 699760 267702 699816
rect 263690 313248 263746 313304
rect 264978 291760 265034 291816
rect 264058 273400 264114 273456
rect 263966 268096 264022 268152
rect 263690 265376 263746 265432
rect 262494 230424 262550 230480
rect 262218 58520 262274 58576
rect 263966 231784 264022 231840
rect 263782 207576 263838 207632
rect 265162 304136 265218 304192
rect 266358 298016 266414 298072
rect 265162 272992 265218 273048
rect 266634 316104 266690 316160
rect 266450 276936 266506 276992
rect 265070 219272 265126 219328
rect 266910 298016 266966 298072
rect 266910 297336 266966 297392
rect 266726 253952 266782 254008
rect 266450 158752 266506 158808
rect 268106 257216 268162 257272
rect 268014 238448 268070 238504
rect 268382 148280 268438 148336
rect 264242 74432 264298 74488
rect 263598 73208 263654 73264
rect 264242 73208 264298 73264
rect 269210 244296 269266 244352
rect 269210 215872 269266 215928
rect 271878 272448 271934 272504
rect 276018 304000 276074 304056
rect 273626 253952 273682 254008
rect 271878 150320 271934 150376
rect 275282 253136 275338 253192
rect 275282 241440 275338 241496
rect 276110 276664 276166 276720
rect 269210 89664 269266 89720
rect 277398 301008 277454 301064
rect 276202 262928 276258 262984
rect 280250 299512 280306 299568
rect 278778 294480 278834 294536
rect 277582 227568 277638 227624
rect 278870 209616 278926 209672
rect 281538 298696 281594 298752
rect 280802 262928 280858 262984
rect 285678 310392 285734 310448
rect 286322 310392 286378 310448
rect 285678 309304 285734 309360
rect 284298 241712 284354 241768
rect 282918 145580 282974 145616
rect 282918 145560 282920 145580
rect 282920 145560 282972 145580
rect 282972 145560 282974 145580
rect 280158 73752 280214 73808
rect 348790 702480 348846 702536
rect 580170 697176 580226 697232
rect 582746 683848 582802 683904
rect 582378 670656 582434 670712
rect 582378 644000 582434 644056
rect 580170 511284 580226 511320
rect 580170 511264 580172 511284
rect 580172 511264 580224 511284
rect 580224 511264 580226 511284
rect 580170 365064 580226 365120
rect 580170 351908 580172 351928
rect 580172 351908 580224 351928
rect 580224 351908 580226 351928
rect 309782 297336 309838 297392
rect 288530 212472 288586 212528
rect 285770 86808 285826 86864
rect 298098 87488 298154 87544
rect 303618 24112 303674 24168
rect 580170 351872 580226 351908
rect 580906 325216 580962 325272
rect 580170 312024 580226 312080
rect 580262 298696 580318 298752
rect 580170 272176 580226 272232
rect 582470 630808 582526 630864
rect 582378 258848 582434 258904
rect 582654 617480 582710 617536
rect 582654 577632 582710 577688
rect 574742 244160 574798 244216
rect 580170 232328 580226 232384
rect 582470 245520 582526 245576
rect 582470 236544 582526 236600
rect 582378 219000 582434 219056
rect 580262 205672 580318 205728
rect 580170 192500 580226 192536
rect 580170 192480 580172 192500
rect 580172 192480 580224 192500
rect 580224 192480 580226 192500
rect 580170 179152 580226 179208
rect 340142 160656 340198 160712
rect 335358 83408 335414 83464
rect 341522 135904 341578 135960
rect 345018 64096 345074 64152
rect 580354 139304 580410 139360
rect 580262 125976 580318 126032
rect 582378 99456 582434 99512
rect 580262 90344 580318 90400
rect 580170 86128 580226 86184
rect 582378 89664 582434 89720
rect 580262 72936 580318 72992
rect 580170 46280 580226 46336
rect 583666 590688 583722 590744
rect 582838 564304 582894 564360
rect 582838 537784 582894 537840
rect 582746 524456 582802 524512
rect 582930 484608 582986 484664
rect 583022 471416 583078 471472
rect 583114 458088 583170 458144
rect 583206 431568 583262 431624
rect 583114 289040 583170 289096
rect 582930 235864 582986 235920
rect 582930 232464 582986 232520
rect 582746 165824 582802 165880
rect 582562 152632 582618 152688
rect 582562 138624 582618 138680
rect 582838 142704 582894 142760
rect 582838 112784 582894 112840
rect 582654 59608 582710 59664
rect 582562 19760 582618 19816
rect 582838 33088 582894 33144
rect 582746 6568 582802 6624
rect 583390 418240 583446 418296
rect 583298 404912 583354 404968
rect 583482 378120 583538 378176
rect 583482 253136 583538 253192
rect 583298 240080 583354 240136
rect 583666 238584 583722 238640
<< metal3 >>
rect 268326 702476 268332 702540
rect 268396 702538 268402 702540
rect 348785 702538 348851 702541
rect 268396 702536 348851 702538
rect 268396 702480 348790 702536
rect 348846 702480 348851 702536
rect 268396 702478 348851 702480
rect 268396 702476 268402 702478
rect 348785 702475 348851 702478
rect 260046 699756 260052 699820
rect 260116 699818 260122 699820
rect 267641 699818 267707 699821
rect 260116 699816 267707 699818
rect 260116 699760 267646 699816
rect 267702 699760 267707 699816
rect 260116 699758 267707 699760
rect 260116 699756 260122 699758
rect 267641 699755 267707 699758
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 582741 683906 582807 683909
rect 583520 683906 584960 683996
rect 582741 683904 584960 683906
rect 582741 683848 582746 683904
rect 582802 683848 584960 683904
rect 582741 683846 584960 683848
rect 582741 683843 582807 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 582373 670714 582439 670717
rect 583520 670714 584960 670804
rect 582373 670712 584960 670714
rect 582373 670656 582378 670712
rect 582434 670656 584960 670712
rect 582373 670654 584960 670656
rect 582373 670651 582439 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3509 658202 3575 658205
rect -960 658200 3575 658202
rect -960 658144 3514 658200
rect 3570 658144 3575 658200
rect -960 658142 3575 658144
rect -960 658052 480 658142
rect 3509 658139 3575 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 582373 644058 582439 644061
rect 583520 644058 584960 644148
rect 582373 644056 584960 644058
rect 582373 644000 582378 644056
rect 582434 644000 584960 644056
rect 582373 643998 584960 644000
rect 582373 643995 582439 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3509 632090 3575 632093
rect -960 632088 3575 632090
rect -960 632032 3514 632088
rect 3570 632032 3575 632088
rect -960 632030 3575 632032
rect -960 631940 480 632030
rect 3509 632027 3575 632030
rect 582465 630866 582531 630869
rect 583520 630866 584960 630956
rect 582465 630864 584960 630866
rect 582465 630808 582470 630864
rect 582526 630808 584960 630864
rect 582465 630806 584960 630808
rect 582465 630803 582531 630806
rect 583520 630716 584960 630806
rect 15837 621618 15903 621621
rect 74574 621618 74580 621620
rect 15837 621616 74580 621618
rect 15837 621560 15842 621616
rect 15898 621560 74580 621616
rect 15837 621558 74580 621560
rect 15837 621555 15903 621558
rect 74574 621556 74580 621558
rect 74644 621556 74650 621620
rect -960 619170 480 619260
rect 3509 619170 3575 619173
rect -960 619168 3575 619170
rect -960 619112 3514 619168
rect 3570 619112 3575 619168
rect -960 619110 3575 619112
rect -960 619020 480 619110
rect 3509 619107 3575 619110
rect 582649 617538 582715 617541
rect 583520 617538 584960 617628
rect 582649 617536 584960 617538
rect 582649 617480 582654 617536
rect 582710 617480 584960 617536
rect 582649 617478 584960 617480
rect 582649 617475 582715 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 2773 606114 2839 606117
rect -960 606112 2839 606114
rect -960 606056 2778 606112
rect 2834 606056 2839 606112
rect -960 606054 2839 606056
rect -960 605964 480 606054
rect 2773 606051 2839 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 76465 591154 76531 591157
rect 77201 591154 77267 591157
rect 76465 591152 77267 591154
rect 76465 591096 76470 591152
rect 76526 591096 77206 591152
rect 77262 591096 77267 591152
rect 76465 591094 77267 591096
rect 76465 591091 76531 591094
rect 77201 591091 77267 591094
rect 583520 591018 584960 591108
rect 583342 590958 584960 591018
rect 583342 590882 583402 590958
rect 583520 590882 584960 590958
rect 583342 590868 584960 590882
rect 583342 590822 583586 590868
rect 77201 590746 77267 590749
rect 125726 590746 125732 590748
rect 77201 590744 125732 590746
rect 77201 590688 77206 590744
rect 77262 590688 125732 590744
rect 77201 590686 125732 590688
rect 77201 590683 77267 590686
rect 125726 590684 125732 590686
rect 125796 590684 125802 590748
rect 583526 590746 583586 590822
rect 583661 590746 583727 590749
rect 583526 590744 583727 590746
rect 583526 590688 583666 590744
rect 583722 590688 583727 590744
rect 583526 590686 583727 590688
rect 583661 590683 583727 590686
rect 71773 584898 71839 584901
rect 76046 584898 76052 584900
rect 71773 584896 76052 584898
rect 71773 584840 71778 584896
rect 71834 584840 76052 584896
rect 71773 584838 76052 584840
rect 71773 584835 71839 584838
rect 76046 584836 76052 584838
rect 76116 584836 76122 584900
rect 72417 582722 72483 582725
rect 132585 582722 132651 582725
rect 72417 582720 132651 582722
rect 72417 582664 72422 582720
rect 72478 582664 132590 582720
rect 132646 582664 132651 582720
rect 72417 582662 132651 582664
rect 72417 582659 72483 582662
rect 132585 582659 132651 582662
rect 88241 582586 88307 582589
rect 100017 582586 100083 582589
rect 88241 582584 100083 582586
rect 88241 582528 88246 582584
rect 88302 582528 100022 582584
rect 100078 582528 100083 582584
rect 88241 582526 100083 582528
rect 88241 582523 88307 582526
rect 100017 582523 100083 582526
rect 69473 582450 69539 582453
rect 70301 582450 70367 582453
rect 69473 582448 70367 582450
rect 69473 582392 69478 582448
rect 69534 582392 70306 582448
rect 70362 582392 70367 582448
rect 69473 582390 70367 582392
rect 69473 582387 69539 582390
rect 70301 582387 70367 582390
rect 74574 582388 74580 582452
rect 74644 582450 74650 582452
rect 74901 582450 74967 582453
rect 74644 582448 74967 582450
rect 74644 582392 74906 582448
rect 74962 582392 74967 582448
rect 74644 582390 74967 582392
rect 74644 582388 74650 582390
rect 74901 582387 74967 582390
rect 59261 581226 59327 581229
rect 82997 581226 83063 581229
rect 59261 581224 83063 581226
rect 59261 581168 59266 581224
rect 59322 581168 83002 581224
rect 83058 581168 83063 581224
rect 59261 581166 83063 581168
rect 59261 581163 59327 581166
rect 82997 581163 83063 581166
rect 79041 581090 79107 581093
rect 102777 581090 102843 581093
rect 79041 581088 102843 581090
rect 79041 581032 79046 581088
rect 79102 581032 102782 581088
rect 102838 581032 102843 581088
rect 79041 581030 102843 581032
rect 79041 581027 79107 581030
rect 102777 581027 102843 581030
rect 75361 580954 75427 580957
rect 75678 580954 75684 580956
rect 75361 580952 75684 580954
rect 75361 580896 75366 580952
rect 75422 580896 75684 580952
rect 75361 580894 75684 580896
rect 75361 580891 75427 580894
rect 75678 580892 75684 580894
rect 75748 580892 75754 580956
rect 70526 580756 70532 580820
rect 70596 580818 70602 580820
rect 70853 580818 70919 580821
rect 79777 580820 79843 580821
rect 79726 580818 79732 580820
rect 70596 580816 70919 580818
rect 70596 580760 70858 580816
rect 70914 580760 70919 580816
rect 70596 580758 70919 580760
rect 79686 580758 79732 580818
rect 79796 580816 79843 580820
rect 79838 580760 79843 580816
rect 70596 580756 70602 580758
rect 70853 580755 70919 580758
rect 79726 580756 79732 580758
rect 79796 580756 79843 580760
rect 83958 580756 83964 580820
rect 84028 580818 84034 580820
rect 84193 580818 84259 580821
rect 84028 580816 84259 580818
rect 84028 580760 84198 580816
rect 84254 580760 84259 580816
rect 84028 580758 84259 580760
rect 84028 580756 84034 580758
rect 79777 580755 79843 580756
rect 84193 580755 84259 580758
rect 88374 580756 88380 580820
rect 88444 580818 88450 580820
rect 88701 580818 88767 580821
rect 88444 580816 88767 580818
rect 88444 580760 88706 580816
rect 88762 580760 88767 580816
rect 88444 580758 88767 580760
rect 88444 580756 88450 580758
rect 88701 580755 88767 580758
rect 91502 580756 91508 580820
rect 91572 580818 91578 580820
rect 92381 580818 92447 580821
rect 91572 580816 92447 580818
rect 91572 580760 92386 580816
rect 92442 580760 92447 580816
rect 91572 580758 92447 580760
rect 91572 580756 91578 580758
rect 92381 580755 92447 580758
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 66805 580002 66871 580005
rect 68878 580002 68938 580584
rect 66805 580000 68938 580002
rect 66805 579944 66810 580000
rect 66866 579944 68938 580000
rect 66805 579942 68938 579944
rect 66805 579939 66871 579942
rect 63401 578914 63467 578917
rect 68645 578914 68711 578917
rect 63401 578912 68711 578914
rect 63401 578856 63406 578912
rect 63462 578856 68650 578912
rect 68706 578856 68711 578912
rect 63401 578854 68711 578856
rect 63401 578851 63467 578854
rect 68645 578851 68711 578854
rect 66805 578642 66871 578645
rect 68878 578642 68938 579224
rect 94638 578914 94698 579496
rect 96889 578914 96955 578917
rect 94638 578912 96955 578914
rect 94638 578856 96894 578912
rect 96950 578856 96955 578912
rect 94638 578854 96955 578856
rect 96889 578851 96955 578854
rect 66805 578640 68938 578642
rect 66805 578584 66810 578640
rect 66866 578584 68938 578640
rect 66805 578582 68938 578584
rect 66805 578579 66871 578582
rect 67449 577282 67515 577285
rect 68878 577282 68938 577864
rect 94638 577554 94698 578136
rect 582649 577690 582715 577693
rect 583520 577690 584960 577780
rect 582649 577688 584960 577690
rect 582649 577632 582654 577688
rect 582710 577632 584960 577688
rect 582649 577630 584960 577632
rect 582649 577627 582715 577630
rect 97073 577554 97139 577557
rect 94638 577552 97139 577554
rect 94638 577496 97078 577552
rect 97134 577496 97139 577552
rect 583520 577540 584960 577630
rect 94638 577494 97139 577496
rect 97073 577491 97139 577494
rect 67449 577280 68938 577282
rect 67449 577224 67454 577280
rect 67510 577224 68938 577280
rect 67449 577222 68938 577224
rect 67449 577219 67515 577222
rect 94638 576738 94698 576776
rect 97901 576738 97967 576741
rect 94638 576736 97967 576738
rect 94638 576680 97906 576736
rect 97962 576680 97967 576736
rect 94638 576678 97967 576680
rect 97901 576675 97967 576678
rect 66529 575922 66595 575925
rect 68878 575922 68938 576504
rect 66529 575920 68938 575922
rect 66529 575864 66534 575920
rect 66590 575864 68938 575920
rect 66529 575862 68938 575864
rect 66529 575859 66595 575862
rect 67541 575378 67607 575381
rect 67541 575376 68938 575378
rect 67541 575320 67546 575376
rect 67602 575320 68938 575376
rect 67541 575318 68938 575320
rect 67541 575315 67607 575318
rect 68878 575144 68938 575318
rect 94638 574834 94698 575416
rect 95233 574834 95299 574837
rect 96245 574834 96311 574837
rect 94638 574832 96311 574834
rect 94638 574776 95238 574832
rect 95294 574776 96250 574832
rect 96306 574776 96311 574832
rect 94638 574774 96311 574776
rect 95233 574771 95299 574774
rect 96245 574771 96311 574774
rect 66437 573202 66503 573205
rect 68878 573202 68938 573784
rect 94638 573474 94698 574056
rect 97901 573474 97967 573477
rect 94638 573472 97967 573474
rect 94638 573416 97906 573472
rect 97962 573416 97967 573472
rect 94638 573414 97967 573416
rect 97901 573411 97967 573414
rect 66437 573200 68938 573202
rect 66437 573144 66442 573200
rect 66498 573144 68938 573200
rect 66437 573142 68938 573144
rect 66437 573139 66503 573142
rect 66713 571842 66779 571845
rect 68878 571842 68938 572424
rect 94638 572250 94698 572696
rect 97257 572250 97323 572253
rect 94638 572248 97323 572250
rect 94638 572192 97262 572248
rect 97318 572192 97323 572248
rect 94638 572190 97323 572192
rect 97257 572187 97323 572190
rect 66713 571840 68938 571842
rect 66713 571784 66718 571840
rect 66774 571784 68938 571840
rect 66713 571782 68938 571784
rect 66713 571779 66779 571782
rect 104934 571434 104940 571436
rect 94638 571374 104940 571434
rect 94638 571336 94698 571374
rect 104934 571372 104940 571374
rect 105004 571372 105010 571436
rect 66897 570210 66963 570213
rect 68878 570210 68938 570792
rect 66897 570208 68938 570210
rect 66897 570152 66902 570208
rect 66958 570152 68938 570208
rect 66897 570150 68938 570152
rect 66897 570147 66963 570150
rect 97901 570074 97967 570077
rect 94638 570072 97967 570074
rect 94638 570016 97906 570072
rect 97962 570016 97967 570072
rect 94638 570014 97967 570016
rect 94638 569976 94698 570014
rect 97901 570011 97967 570014
rect 65977 568850 66043 568853
rect 68878 568850 68938 569432
rect 96613 569122 96679 569125
rect 97901 569122 97967 569125
rect 65977 568848 68938 568850
rect 65977 568792 65982 568848
rect 66038 568792 68938 568848
rect 65977 568790 68938 568792
rect 94638 569120 97967 569122
rect 94638 569064 96618 569120
rect 96674 569064 97906 569120
rect 97962 569064 97967 569120
rect 94638 569062 97967 569064
rect 65977 568787 66043 568790
rect 94638 568616 94698 569062
rect 96613 569059 96679 569062
rect 97901 569059 97967 569062
rect 66989 567490 67055 567493
rect 68878 567490 68938 568072
rect 66989 567488 68938 567490
rect 66989 567432 66994 567488
rect 67050 567432 68938 567488
rect 66989 567430 68938 567432
rect 66989 567427 67055 567430
rect 94086 567084 94146 567256
rect -960 566946 480 567036
rect 94078 567020 94084 567084
rect 94148 567020 94154 567084
rect 3417 566946 3483 566949
rect -960 566944 3483 566946
rect -960 566888 3422 566944
rect 3478 566888 3483 566944
rect -960 566886 3483 566888
rect -960 566796 480 566886
rect 3417 566883 3483 566886
rect 67633 566674 67699 566677
rect 68878 566674 68938 566712
rect 67633 566672 68938 566674
rect 67633 566616 67638 566672
rect 67694 566616 68938 566672
rect 67633 566614 68938 566616
rect 67633 566611 67699 566614
rect 94638 565858 94698 565896
rect 95417 565858 95483 565861
rect 94638 565856 95483 565858
rect 94638 565800 95422 565856
rect 95478 565800 95483 565856
rect 94638 565798 95483 565800
rect 95417 565795 95483 565798
rect 66713 564770 66779 564773
rect 68878 564770 68938 565352
rect 66713 564768 68938 564770
rect 66713 564712 66718 564768
rect 66774 564712 68938 564768
rect 66713 564710 68938 564712
rect 66713 564707 66779 564710
rect 582833 564362 582899 564365
rect 583520 564362 584960 564452
rect 582833 564360 584960 564362
rect 582833 564304 582838 564360
rect 582894 564304 584960 564360
rect 582833 564302 584960 564304
rect 582833 564299 582899 564302
rect 66437 564226 66503 564229
rect 66437 564224 68938 564226
rect 66437 564168 66442 564224
rect 66498 564168 68938 564224
rect 66437 564166 68938 564168
rect 66437 564163 66503 564166
rect 68878 563992 68938 564166
rect 94638 563682 94698 564264
rect 583520 564212 584960 564302
rect 94773 563682 94839 563685
rect 94638 563680 94839 563682
rect 94638 563624 94778 563680
rect 94834 563624 94839 563680
rect 94638 563622 94839 563624
rect 94773 563619 94839 563622
rect 66161 562050 66227 562053
rect 68878 562050 68938 562632
rect 94638 562322 94698 562904
rect 97349 562322 97415 562325
rect 94638 562320 97415 562322
rect 94638 562264 97354 562320
rect 97410 562264 97415 562320
rect 94638 562262 97415 562264
rect 97349 562259 97415 562262
rect 66161 562048 68938 562050
rect 66161 561992 66166 562048
rect 66222 561992 68938 562048
rect 66161 561990 68938 561992
rect 66161 561987 66227 561990
rect 66989 560690 67055 560693
rect 68878 560690 68938 561272
rect 94638 560962 94698 561544
rect 96797 560962 96863 560965
rect 94638 560960 96863 560962
rect 94638 560904 96802 560960
rect 96858 560904 96863 560960
rect 94638 560902 96863 560904
rect 96797 560899 96863 560902
rect 66989 560688 68938 560690
rect 66989 560632 66994 560688
rect 67050 560632 68938 560688
rect 66989 560630 68938 560632
rect 66989 560627 67055 560630
rect 66989 559330 67055 559333
rect 68878 559330 68938 559912
rect 94638 559466 94698 560184
rect 110638 559466 110644 559468
rect 94638 559406 110644 559466
rect 110638 559404 110644 559406
rect 110708 559404 110714 559468
rect 66989 559328 68938 559330
rect 66989 559272 66994 559328
rect 67050 559272 68938 559328
rect 66989 559270 68938 559272
rect 66989 559267 67055 559270
rect 95325 558922 95391 558925
rect 95877 558922 95943 558925
rect 94638 558920 95943 558922
rect 94638 558864 95330 558920
rect 95386 558864 95882 558920
rect 95938 558864 95943 558920
rect 94638 558862 95943 558864
rect 94638 558824 94698 558862
rect 95325 558859 95391 558862
rect 95877 558859 95943 558862
rect 66989 557970 67055 557973
rect 68878 557970 68938 558552
rect 66989 557968 68938 557970
rect 66989 557912 66994 557968
rect 67050 557912 68938 557968
rect 66989 557910 68938 557912
rect 66989 557907 67055 557910
rect 67817 556610 67883 556613
rect 68878 556610 68938 557192
rect 94638 556882 94698 557464
rect 96705 556882 96771 556885
rect 94638 556880 96771 556882
rect 94638 556824 96710 556880
rect 96766 556824 96771 556880
rect 94638 556822 96771 556824
rect 96705 556819 96771 556822
rect 67817 556608 68938 556610
rect 67817 556552 67822 556608
rect 67878 556552 68938 556608
rect 67817 556550 68938 556552
rect 67817 556547 67883 556550
rect 66989 555250 67055 555253
rect 68878 555250 68938 555832
rect 94638 555522 94698 556104
rect 95325 555522 95391 555525
rect 94638 555520 95391 555522
rect 94638 555464 95330 555520
rect 95386 555464 95391 555520
rect 94638 555462 95391 555464
rect 95325 555459 95391 555462
rect 66989 555248 68938 555250
rect 66989 555192 66994 555248
rect 67050 555192 68938 555248
rect 66989 555190 68938 555192
rect 66989 555187 67055 555190
rect -960 553890 480 553980
rect 3509 553890 3575 553893
rect -960 553888 3575 553890
rect -960 553832 3514 553888
rect 3570 553832 3575 553888
rect -960 553830 3575 553832
rect -960 553740 480 553830
rect 3509 553827 3575 553830
rect 66989 553618 67055 553621
rect 68878 553618 68938 554200
rect 94638 554162 94698 554744
rect 96889 554162 96955 554165
rect 94638 554160 96955 554162
rect 94638 554104 96894 554160
rect 96950 554104 96955 554160
rect 94638 554102 96955 554104
rect 96889 554099 96955 554102
rect 66989 553616 68938 553618
rect 66989 553560 66994 553616
rect 67050 553560 68938 553616
rect 66989 553558 68938 553560
rect 66989 553555 67055 553558
rect 67725 552258 67791 552261
rect 68878 552258 68938 552840
rect 94638 552802 94698 553384
rect 96981 552802 97047 552805
rect 94638 552800 97047 552802
rect 94638 552744 96986 552800
rect 97042 552744 97047 552800
rect 94638 552742 97047 552744
rect 96981 552739 97047 552742
rect 94681 552530 94747 552533
rect 67725 552256 68938 552258
rect 67725 552200 67730 552256
rect 67786 552200 68938 552256
rect 67725 552198 68938 552200
rect 94638 552528 94747 552530
rect 94638 552472 94686 552528
rect 94742 552472 94747 552528
rect 94638 552467 94747 552472
rect 67725 552195 67791 552198
rect 94638 552122 94698 552467
rect 96613 552122 96679 552125
rect 94638 552120 96679 552122
rect 94638 552064 96618 552120
rect 96674 552064 96679 552120
rect 94638 552062 96679 552064
rect 94638 552024 94698 552062
rect 96613 552059 96679 552062
rect 67633 550898 67699 550901
rect 68878 550898 68938 551480
rect 583520 551020 584960 551260
rect 67633 550896 68938 550898
rect 67633 550840 67638 550896
rect 67694 550840 68938 550896
rect 67633 550838 68938 550840
rect 67633 550835 67699 550838
rect 97901 550762 97967 550765
rect 94638 550760 97967 550762
rect 94638 550704 97906 550760
rect 97962 550704 97967 550760
rect 94638 550702 97967 550704
rect 94638 550664 94698 550702
rect 97901 550699 97967 550702
rect 66529 549538 66595 549541
rect 68878 549538 68938 550120
rect 66529 549536 68938 549538
rect 66529 549480 66534 549536
rect 66590 549480 68938 549536
rect 66529 549478 68938 549480
rect 66529 549475 66595 549478
rect 100702 549402 100708 549404
rect 94638 549342 100708 549402
rect 94638 549304 94698 549342
rect 100702 549340 100708 549342
rect 100772 549340 100778 549404
rect 69062 548316 69122 548760
rect 69054 548252 69060 548316
rect 69124 548252 69130 548316
rect 66989 546818 67055 546821
rect 68878 546818 68938 547400
rect 94638 547090 94698 547672
rect 96654 547090 96660 547092
rect 94638 547030 96660 547090
rect 96654 547028 96660 547030
rect 96724 547028 96730 547092
rect 66989 546816 68938 546818
rect 66989 546760 66994 546816
rect 67050 546760 68938 546816
rect 66989 546758 68938 546760
rect 66989 546755 67055 546758
rect 66069 546002 66135 546005
rect 68878 546002 68938 546040
rect 66069 546000 68938 546002
rect 66069 545944 66074 546000
rect 66130 545944 68938 546000
rect 66069 545942 68938 545944
rect 66069 545939 66135 545942
rect 94638 545730 94698 546312
rect 96705 545730 96771 545733
rect 94638 545728 96771 545730
rect 94638 545672 96710 545728
rect 96766 545672 96771 545728
rect 94638 545670 96771 545672
rect 96705 545667 96771 545670
rect 66713 544642 66779 544645
rect 68878 544642 68938 544680
rect 66713 544640 68938 544642
rect 66713 544584 66718 544640
rect 66774 544584 68938 544640
rect 66713 544582 68938 544584
rect 66713 544579 66779 544582
rect 94638 544370 94698 544952
rect 97533 544370 97599 544373
rect 94638 544368 97599 544370
rect 94638 544312 97538 544368
rect 97594 544312 97599 544368
rect 94638 544310 97599 544312
rect 97533 544307 97599 544310
rect 4797 542466 4863 542469
rect 67766 542466 67772 542468
rect 4797 542464 67772 542466
rect 4797 542408 4802 542464
rect 4858 542408 67772 542464
rect 4797 542406 67772 542408
rect 4797 542403 4863 542406
rect 67766 542404 67772 542406
rect 67836 542466 67842 542468
rect 68878 542466 68938 543320
rect 94638 543010 94698 543592
rect 98085 543010 98151 543013
rect 94638 543008 98151 543010
rect 94638 542952 98090 543008
rect 98146 542952 98151 543008
rect 94638 542950 98151 542952
rect 98085 542947 98151 542950
rect 67836 542406 68938 542466
rect 67836 542404 67842 542406
rect 69422 542132 69428 542196
rect 69492 542132 69498 542196
rect 17217 541106 17283 541109
rect 69430 541106 69490 542132
rect 94638 541650 94698 542232
rect 96838 541650 96844 541652
rect 94638 541590 96844 541650
rect 96838 541588 96844 541590
rect 96908 541588 96914 541652
rect 17217 541104 69490 541106
rect 17217 541048 17222 541104
rect 17278 541048 69490 541104
rect 17217 541046 69490 541048
rect 17217 541043 17283 541046
rect -960 540684 480 540924
rect 69430 539882 69490 540600
rect 94638 540293 94698 540872
rect 94638 540288 94747 540293
rect 94638 540232 94686 540288
rect 94742 540232 94747 540288
rect 94638 540230 94747 540232
rect 94681 540227 94747 540230
rect 69430 539822 69674 539882
rect 69614 539746 69674 539822
rect 70301 539746 70367 539749
rect 69614 539744 70367 539746
rect 69614 539688 70306 539744
rect 70362 539688 70367 539744
rect 69614 539686 70367 539688
rect 70301 539683 70367 539686
rect 76046 539548 76052 539612
rect 76116 539610 76122 539612
rect 76741 539610 76807 539613
rect 76116 539608 76807 539610
rect 76116 539552 76746 539608
rect 76802 539552 76807 539608
rect 76116 539550 76807 539552
rect 76116 539548 76122 539550
rect 76741 539547 76807 539550
rect 93945 538930 94011 538933
rect 94086 538930 94146 539512
rect 93945 538928 94146 538930
rect 93945 538872 93950 538928
rect 94006 538872 94146 538928
rect 93945 538870 94146 538872
rect 93945 538867 94011 538870
rect 582833 537842 582899 537845
rect 583520 537842 584960 537932
rect 582833 537840 584960 537842
rect 582833 537784 582838 537840
rect 582894 537784 584960 537840
rect 582833 537782 584960 537784
rect 582833 537779 582899 537782
rect 583520 537692 584960 537782
rect 76465 536754 76531 536757
rect 116577 536754 116643 536757
rect 76465 536752 116643 536754
rect 76465 536696 76470 536752
rect 76526 536696 116582 536752
rect 116638 536696 116643 536752
rect 76465 536694 116643 536696
rect 76465 536691 76531 536694
rect 116577 536691 116643 536694
rect 76465 535666 76531 535669
rect 77201 535666 77267 535669
rect 76465 535664 77267 535666
rect 76465 535608 76470 535664
rect 76526 535608 77206 535664
rect 77262 535608 77267 535664
rect 76465 535606 77267 535608
rect 76465 535603 76531 535606
rect 77201 535603 77267 535606
rect 76097 535530 76163 535533
rect 76741 535530 76807 535533
rect 76097 535528 76807 535530
rect 76097 535472 76102 535528
rect 76158 535472 76746 535528
rect 76802 535472 76807 535528
rect 76097 535470 76807 535472
rect 76097 535467 76163 535470
rect 76741 535467 76807 535470
rect 74441 534714 74507 534717
rect 111742 534714 111748 534716
rect 74441 534712 111748 534714
rect 74441 534656 74446 534712
rect 74502 534656 111748 534712
rect 74441 534654 111748 534656
rect 74441 534651 74507 534654
rect 111742 534652 111748 534654
rect 111812 534652 111818 534716
rect 39849 531994 39915 531997
rect 96838 531994 96844 531996
rect 39849 531992 96844 531994
rect 39849 531936 39854 531992
rect 39910 531936 96844 531992
rect 39849 531934 96844 531936
rect 39849 531931 39915 531934
rect 96838 531932 96844 531934
rect 96908 531932 96914 531996
rect 79910 530708 79916 530772
rect 79980 530770 79986 530772
rect 93894 530770 93900 530772
rect 79980 530710 93900 530770
rect 79980 530708 79986 530710
rect 93894 530708 93900 530710
rect 93964 530708 93970 530772
rect 43989 530634 44055 530637
rect 96654 530634 96660 530636
rect 43989 530632 96660 530634
rect 43989 530576 43994 530632
rect 44050 530576 96660 530632
rect 43989 530574 96660 530576
rect 43989 530571 44055 530574
rect 96654 530572 96660 530574
rect 96724 530572 96730 530636
rect -960 527914 480 528004
rect 3509 527914 3575 527917
rect -960 527912 3575 527914
rect -960 527856 3514 527912
rect 3570 527856 3575 527912
rect -960 527854 3575 527856
rect -960 527764 480 527854
rect 3509 527851 3575 527854
rect 73470 524996 73476 525060
rect 73540 525058 73546 525060
rect 91502 525058 91508 525060
rect 73540 524998 91508 525058
rect 73540 524996 73546 524998
rect 91502 524996 91508 524998
rect 91572 524996 91578 525060
rect 582741 524514 582807 524517
rect 583520 524514 584960 524604
rect 582741 524512 584960 524514
rect 582741 524456 582746 524512
rect 582802 524456 584960 524512
rect 582741 524454 584960 524456
rect 582741 524451 582807 524454
rect 583520 524364 584960 524454
rect 77150 523636 77156 523700
rect 77220 523698 77226 523700
rect 95325 523698 95391 523701
rect 77220 523696 95391 523698
rect 77220 523640 95330 523696
rect 95386 523640 95391 523696
rect 77220 523638 95391 523640
rect 77220 523636 77226 523638
rect 95325 523635 95391 523638
rect 76557 522338 76623 522341
rect 102174 522338 102180 522340
rect 76557 522336 102180 522338
rect 76557 522280 76562 522336
rect 76618 522280 102180 522336
rect 76557 522278 102180 522280
rect 76557 522275 76623 522278
rect 102174 522276 102180 522278
rect 102244 522276 102250 522340
rect -960 514858 480 514948
rect 3509 514858 3575 514861
rect -960 514856 3575 514858
rect -960 514800 3514 514856
rect 3570 514800 3575 514856
rect -960 514798 3575 514800
rect -960 514708 480 514798
rect 3509 514795 3575 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3417 501802 3483 501805
rect -960 501800 3483 501802
rect -960 501744 3422 501800
rect 3478 501744 3483 501800
rect -960 501742 3483 501744
rect -960 501652 480 501742
rect 3417 501739 3483 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 582925 484666 582991 484669
rect 583520 484666 584960 484756
rect 582925 484664 584960 484666
rect 582925 484608 582930 484664
rect 582986 484608 584960 484664
rect 582925 484606 584960 484608
rect 582925 484603 582991 484606
rect 583520 484516 584960 484606
rect 81433 479498 81499 479501
rect 107694 479498 107700 479500
rect 81433 479496 107700 479498
rect 81433 479440 81438 479496
rect 81494 479440 107700 479496
rect 81433 479438 107700 479440
rect 81433 479435 81499 479438
rect 107694 479436 107700 479438
rect 107764 479436 107770 479500
rect 72601 476778 72667 476781
rect 100150 476778 100156 476780
rect 72601 476776 100156 476778
rect 72601 476720 72606 476776
rect 72662 476720 100156 476776
rect 72601 476718 100156 476720
rect 72601 476715 72667 476718
rect 100150 476716 100156 476718
rect 100220 476716 100226 476780
rect -960 475690 480 475780
rect 3417 475690 3483 475693
rect -960 475688 3483 475690
rect -960 475632 3422 475688
rect 3478 475632 3483 475688
rect -960 475630 3483 475632
rect -960 475540 480 475630
rect 3417 475627 3483 475630
rect 72366 473996 72372 474060
rect 72436 474058 72442 474060
rect 94773 474058 94839 474061
rect 72436 474056 94839 474058
rect 72436 474000 94778 474056
rect 94834 474000 94839 474056
rect 72436 473998 94839 474000
rect 72436 473996 72442 473998
rect 94773 473995 94839 473998
rect 81934 471820 81940 471884
rect 82004 471882 82010 471884
rect 83958 471882 83964 471884
rect 82004 471822 83964 471882
rect 82004 471820 82010 471822
rect 83958 471820 83964 471822
rect 84028 471820 84034 471884
rect 583017 471474 583083 471477
rect 583520 471474 584960 471564
rect 583017 471472 584960 471474
rect 583017 471416 583022 471472
rect 583078 471416 584960 471472
rect 583017 471414 584960 471416
rect 583017 471411 583083 471414
rect 583520 471324 584960 471414
rect 88425 468618 88491 468621
rect 106406 468618 106412 468620
rect 88425 468616 106412 468618
rect 88425 468560 88430 468616
rect 88486 468560 106412 468616
rect 88425 468558 106412 468560
rect 88425 468555 88491 468558
rect 106406 468556 106412 468558
rect 106476 468556 106482 468620
rect 69606 468420 69612 468484
rect 69676 468482 69682 468484
rect 88742 468482 88748 468484
rect 69676 468422 88748 468482
rect 69676 468420 69682 468422
rect 88742 468420 88748 468422
rect 88812 468420 88818 468484
rect 75678 462844 75684 462908
rect 75748 462906 75754 462908
rect 93894 462906 93900 462908
rect 75748 462846 93900 462906
rect 75748 462844 75754 462846
rect 93894 462844 93900 462846
rect 93964 462844 93970 462908
rect -960 462634 480 462724
rect 3509 462634 3575 462637
rect -960 462632 3575 462634
rect -960 462576 3514 462632
rect 3570 462576 3575 462632
rect -960 462574 3575 462576
rect -960 462484 480 462574
rect 3509 462571 3575 462574
rect 583109 458146 583175 458149
rect 583520 458146 584960 458236
rect 583109 458144 584960 458146
rect 583109 458088 583114 458144
rect 583170 458088 584960 458144
rect 583109 458086 584960 458088
rect 583109 458083 583175 458086
rect 583520 457996 584960 458086
rect 79726 456044 79732 456108
rect 79796 456106 79802 456108
rect 80094 456106 80100 456108
rect 79796 456046 80100 456106
rect 79796 456044 79802 456046
rect 80094 456044 80100 456046
rect 80164 456044 80170 456108
rect 80053 450530 80119 450533
rect 114318 450530 114324 450532
rect 80053 450528 114324 450530
rect 80053 450472 80058 450528
rect 80114 450472 114324 450528
rect 80053 450470 114324 450472
rect 80053 450467 80119 450470
rect 114318 450468 114324 450470
rect 114388 450468 114394 450532
rect 65885 449986 65951 449989
rect 67766 449986 67772 449988
rect 65885 449984 67772 449986
rect 65885 449928 65890 449984
rect 65946 449928 67772 449984
rect 65885 449926 67772 449928
rect 65885 449923 65951 449926
rect 67766 449924 67772 449926
rect 67836 449986 67842 449988
rect 68921 449986 68987 449989
rect 67836 449984 68987 449986
rect 67836 449928 68926 449984
rect 68982 449928 68987 449984
rect 67836 449926 68987 449928
rect 67836 449924 67842 449926
rect 68921 449923 68987 449926
rect -960 449578 480 449668
rect 3141 449578 3207 449581
rect -960 449576 3207 449578
rect -960 449520 3146 449576
rect 3202 449520 3207 449576
rect -960 449518 3207 449520
rect -960 449428 480 449518
rect 3141 449515 3207 449518
rect 583520 444668 584960 444908
rect 67766 442852 67772 442916
rect 67836 442914 67842 442916
rect 70526 442914 70532 442916
rect 67836 442854 70532 442914
rect 67836 442852 67842 442854
rect 70526 442852 70532 442854
rect 70596 442852 70602 442916
rect 71446 441628 71452 441692
rect 71516 441690 71522 441692
rect 76097 441690 76163 441693
rect 71516 441688 76163 441690
rect 71516 441632 76102 441688
rect 76158 441632 76163 441688
rect 71516 441630 76163 441632
rect 71516 441628 71522 441630
rect 76097 441627 76163 441630
rect 88425 440330 88491 440333
rect 115974 440330 115980 440332
rect 88425 440328 115980 440330
rect 88425 440272 88430 440328
rect 88486 440272 115980 440328
rect 88425 440270 115980 440272
rect 88425 440267 88491 440270
rect 115974 440268 115980 440270
rect 116044 440268 116050 440332
rect 98637 439514 98703 439517
rect 109534 439514 109540 439516
rect 98637 439512 109540 439514
rect 98637 439456 98642 439512
rect 98698 439456 109540 439512
rect 98637 439454 109540 439456
rect 98637 439451 98703 439454
rect 109534 439452 109540 439454
rect 109604 439452 109610 439516
rect 81341 438154 81407 438157
rect 88374 438154 88380 438156
rect 81341 438152 88380 438154
rect 81341 438096 81346 438152
rect 81402 438096 88380 438152
rect 81341 438094 88380 438096
rect 81341 438091 81407 438094
rect 88374 438092 88380 438094
rect 88444 438092 88450 438156
rect 94497 437610 94563 437613
rect 94497 437608 97090 437610
rect 94497 437552 94502 437608
rect 94558 437552 97090 437608
rect 94497 437550 97090 437552
rect 94497 437547 94563 437550
rect 97030 437477 97090 437550
rect 78397 437476 78463 437477
rect 78397 437472 78444 437476
rect 78508 437474 78514 437476
rect 78397 437416 78402 437472
rect 78397 437412 78444 437416
rect 78508 437414 78554 437474
rect 97030 437472 97139 437477
rect 97030 437416 97078 437472
rect 97134 437416 97139 437472
rect 97030 437414 97139 437416
rect 78508 437412 78514 437414
rect 78397 437411 78463 437412
rect 97073 437411 97139 437414
rect 107561 437474 107627 437477
rect 114645 437474 114711 437477
rect 107561 437472 114711 437474
rect 107561 437416 107566 437472
rect 107622 437416 114650 437472
rect 114706 437416 114711 437472
rect 107561 437414 114711 437416
rect 107561 437411 107627 437414
rect 114645 437411 114711 437414
rect 77385 437202 77451 437205
rect 78029 437202 78095 437205
rect 77385 437200 78095 437202
rect 77385 437144 77390 437200
rect 77446 437144 78034 437200
rect 78090 437144 78095 437200
rect 77385 437142 78095 437144
rect 77385 437139 77451 437142
rect 78029 437139 78095 437142
rect -960 436508 480 436748
rect 71630 436324 71636 436388
rect 71700 436386 71706 436388
rect 77477 436386 77543 436389
rect 71700 436384 77543 436386
rect 71700 436328 77482 436384
rect 77538 436328 77543 436384
rect 71700 436326 77543 436328
rect 71700 436324 71706 436326
rect 77477 436323 77543 436326
rect 90214 436324 90220 436388
rect 90284 436386 90290 436388
rect 100753 436386 100819 436389
rect 90284 436384 100819 436386
rect 90284 436328 100758 436384
rect 100814 436328 100819 436384
rect 90284 436326 100819 436328
rect 90284 436324 90290 436326
rect 100753 436323 100819 436326
rect 103329 436386 103395 436389
rect 110413 436386 110479 436389
rect 103329 436384 110479 436386
rect 103329 436328 103334 436384
rect 103390 436328 110418 436384
rect 110474 436328 110479 436384
rect 103329 436326 110479 436328
rect 103329 436323 103395 436326
rect 110413 436323 110479 436326
rect 68921 436250 68987 436253
rect 71037 436250 71103 436253
rect 68921 436248 71103 436250
rect 68921 436192 68926 436248
rect 68982 436192 71042 436248
rect 71098 436192 71103 436248
rect 68921 436190 71103 436192
rect 68921 436187 68987 436190
rect 71037 436187 71103 436190
rect 72734 436188 72740 436252
rect 72804 436250 72810 436252
rect 77385 436250 77451 436253
rect 72804 436248 77451 436250
rect 72804 436192 77390 436248
rect 77446 436192 77451 436248
rect 72804 436190 77451 436192
rect 72804 436188 72810 436190
rect 77385 436187 77451 436190
rect 83406 436188 83412 436252
rect 83476 436250 83482 436252
rect 89897 436250 89963 436253
rect 83476 436248 89963 436250
rect 83476 436192 89902 436248
rect 89958 436192 89963 436248
rect 83476 436190 89963 436192
rect 83476 436188 83482 436190
rect 89897 436187 89963 436190
rect 94998 436188 95004 436252
rect 95068 436250 95074 436252
rect 104893 436250 104959 436253
rect 95068 436248 104959 436250
rect 95068 436192 104898 436248
rect 104954 436192 104959 436248
rect 95068 436190 104959 436192
rect 95068 436188 95074 436190
rect 104893 436187 104959 436190
rect 48129 436114 48195 436117
rect 69054 436114 69060 436116
rect 48129 436112 69060 436114
rect 48129 436056 48134 436112
rect 48190 436056 69060 436112
rect 48129 436054 69060 436056
rect 48129 436051 48195 436054
rect 69054 436052 69060 436054
rect 69124 436114 69130 436116
rect 69933 436114 69999 436117
rect 69124 436112 69999 436114
rect 69124 436056 69938 436112
rect 69994 436056 69999 436112
rect 69124 436054 69999 436056
rect 69124 436052 69130 436054
rect 69933 436051 69999 436054
rect 78438 436052 78444 436116
rect 78508 436114 78514 436116
rect 83733 436114 83799 436117
rect 78508 436112 83799 436114
rect 78508 436056 83738 436112
rect 83794 436056 83799 436112
rect 78508 436054 83799 436056
rect 78508 436052 78514 436054
rect 83733 436051 83799 436054
rect 85665 436114 85731 436117
rect 86309 436114 86375 436117
rect 85665 436112 86375 436114
rect 85665 436056 85670 436112
rect 85726 436056 86314 436112
rect 86370 436056 86375 436112
rect 85665 436054 86375 436056
rect 85665 436051 85731 436054
rect 86309 436051 86375 436054
rect 87137 436114 87203 436117
rect 88241 436114 88307 436117
rect 87137 436112 88307 436114
rect 87137 436056 87142 436112
rect 87198 436056 88246 436112
rect 88302 436056 88307 436112
rect 87137 436054 88307 436056
rect 87137 436051 87203 436054
rect 88241 436051 88307 436054
rect 93894 436052 93900 436116
rect 93964 436114 93970 436116
rect 94405 436114 94471 436117
rect 103329 436116 103395 436117
rect 103278 436114 103284 436116
rect 93964 436112 94471 436114
rect 93964 436056 94410 436112
rect 94466 436056 94471 436112
rect 93964 436054 94471 436056
rect 103238 436054 103284 436114
rect 103348 436112 103395 436116
rect 103390 436056 103395 436112
rect 93964 436052 93970 436054
rect 94405 436051 94471 436054
rect 103278 436052 103284 436054
rect 103348 436052 103395 436056
rect 103329 436051 103395 436052
rect 104341 436114 104407 436117
rect 105118 436114 105124 436116
rect 104341 436112 105124 436114
rect 104341 436056 104346 436112
rect 104402 436056 105124 436112
rect 104341 436054 105124 436056
rect 104341 436051 104407 436054
rect 105118 436052 105124 436054
rect 105188 436052 105194 436116
rect 73654 435236 73660 435300
rect 73724 435298 73730 435300
rect 80237 435298 80303 435301
rect 73724 435296 80303 435298
rect 73724 435240 80242 435296
rect 80298 435240 80303 435296
rect 73724 435238 80303 435240
rect 73724 435236 73730 435238
rect 80237 435235 80303 435238
rect 63309 434754 63375 434757
rect 73429 434754 73495 434757
rect 63309 434752 73495 434754
rect 63309 434696 63314 434752
rect 63370 434696 73434 434752
rect 73490 434696 73495 434752
rect 63309 434694 73495 434696
rect 63309 434691 63375 434694
rect 73429 434691 73495 434694
rect 92974 434556 92980 434620
rect 93044 434618 93050 434620
rect 95279 434618 95345 434621
rect 93044 434616 95345 434618
rect 93044 434560 95284 434616
rect 95340 434560 95345 434616
rect 93044 434558 95345 434560
rect 93044 434556 93050 434558
rect 95279 434555 95345 434558
rect 80646 434420 80652 434484
rect 80716 434482 80722 434484
rect 81341 434482 81407 434485
rect 80716 434480 81407 434482
rect 80716 434424 81346 434480
rect 81402 434424 81407 434480
rect 80716 434422 81407 434424
rect 80716 434420 80722 434422
rect 81341 434419 81407 434422
rect 74574 434284 74580 434348
rect 74644 434346 74650 434348
rect 74717 434346 74783 434349
rect 74644 434344 74783 434346
rect 74644 434288 74722 434344
rect 74778 434288 74783 434344
rect 74644 434286 74783 434288
rect 74644 434284 74650 434286
rect 74717 434283 74783 434286
rect 75862 434284 75868 434348
rect 75932 434346 75938 434348
rect 76189 434346 76255 434349
rect 75932 434344 76255 434346
rect 75932 434288 76194 434344
rect 76250 434288 76255 434344
rect 75932 434286 76255 434288
rect 75932 434284 75938 434286
rect 76189 434283 76255 434286
rect 94773 434348 94839 434349
rect 96337 434348 96403 434349
rect 94773 434344 94820 434348
rect 94884 434346 94890 434348
rect 96286 434346 96292 434348
rect 94773 434288 94778 434344
rect 94773 434284 94820 434288
rect 94884 434286 94930 434346
rect 96246 434286 96292 434346
rect 96356 434344 96403 434348
rect 96398 434288 96403 434344
rect 94884 434284 94890 434286
rect 96286 434284 96292 434286
rect 96356 434284 96403 434288
rect 108982 434284 108988 434348
rect 109052 434346 109058 434348
rect 109401 434346 109467 434349
rect 109052 434344 109467 434346
rect 109052 434288 109406 434344
rect 109462 434288 109467 434344
rect 109052 434286 109467 434288
rect 109052 434284 109058 434286
rect 94773 434283 94839 434284
rect 96337 434283 96403 434284
rect 109401 434283 109467 434286
rect 92657 434212 92723 434213
rect 92606 434210 92612 434212
rect 92566 434150 92612 434210
rect 92676 434208 92723 434212
rect 92718 434152 92723 434208
rect 92606 434148 92612 434150
rect 92676 434148 92723 434152
rect 96838 434148 96844 434212
rect 96908 434210 96914 434212
rect 96981 434210 97047 434213
rect 96908 434208 97047 434210
rect 96908 434152 96986 434208
rect 97042 434152 97047 434208
rect 96908 434150 97047 434152
rect 96908 434148 96914 434150
rect 92657 434147 92723 434148
rect 96981 434147 97047 434150
rect 96470 434012 96476 434076
rect 96540 434074 96546 434076
rect 108941 434074 109007 434077
rect 96540 434072 109007 434074
rect 96540 434016 108946 434072
rect 109002 434016 109007 434072
rect 96540 434014 109007 434016
rect 96540 434012 96546 434014
rect 108941 434011 109007 434014
rect 109534 434012 109540 434076
rect 109604 434074 109610 434076
rect 112110 434074 112116 434076
rect 109604 434014 112116 434074
rect 109604 434012 109610 434014
rect 112110 434012 112116 434014
rect 112180 434012 112186 434076
rect 82670 433876 82676 433940
rect 82740 433938 82746 433940
rect 91461 433938 91527 433941
rect 82740 433936 91527 433938
rect 82740 433880 91466 433936
rect 91522 433880 91527 433936
rect 82740 433878 91527 433880
rect 82740 433876 82746 433878
rect 91461 433875 91527 433878
rect 97206 433876 97212 433940
rect 97276 433938 97282 433940
rect 99189 433938 99255 433941
rect 97276 433936 99255 433938
rect 97276 433880 99194 433936
rect 99250 433880 99255 433936
rect 97276 433878 99255 433880
rect 97276 433876 97282 433878
rect 99189 433875 99255 433878
rect 75678 433740 75684 433804
rect 75748 433802 75754 433804
rect 83181 433802 83247 433805
rect 75748 433800 83247 433802
rect 75748 433744 83186 433800
rect 83242 433744 83247 433800
rect 75748 433742 83247 433744
rect 75748 433740 75754 433742
rect 83181 433739 83247 433742
rect 86166 433740 86172 433804
rect 86236 433802 86242 433804
rect 87321 433802 87387 433805
rect 86236 433800 87387 433802
rect 86236 433744 87326 433800
rect 87382 433744 87387 433800
rect 86236 433742 87387 433744
rect 86236 433740 86242 433742
rect 87321 433739 87387 433742
rect 91318 433740 91324 433804
rect 91388 433802 91394 433804
rect 92933 433802 92999 433805
rect 91388 433800 92999 433802
rect 91388 433744 92938 433800
rect 92994 433744 92999 433800
rect 91388 433742 92999 433744
rect 91388 433740 91394 433742
rect 92933 433739 92999 433742
rect 98361 433802 98427 433805
rect 98494 433802 98500 433804
rect 98361 433800 98500 433802
rect 98361 433744 98366 433800
rect 98422 433744 98500 433800
rect 98361 433742 98500 433744
rect 98361 433739 98427 433742
rect 98494 433740 98500 433742
rect 98564 433740 98570 433804
rect 108430 433740 108436 433804
rect 108500 433802 108506 433804
rect 108500 433742 112178 433802
rect 108500 433740 108506 433742
rect 68921 433666 68987 433669
rect 64830 433664 68987 433666
rect 64830 433608 68926 433664
rect 68982 433608 68987 433664
rect 64830 433606 68987 433608
rect 54937 433530 55003 433533
rect 64830 433530 64890 433606
rect 68921 433603 68987 433606
rect 69606 433604 69612 433668
rect 69676 433666 69682 433668
rect 75453 433666 75519 433669
rect 69676 433664 75519 433666
rect 69676 433608 75458 433664
rect 75514 433608 75519 433664
rect 69676 433606 75519 433608
rect 69676 433604 69682 433606
rect 75453 433603 75519 433606
rect 77334 433604 77340 433668
rect 77404 433666 77410 433668
rect 78213 433666 78279 433669
rect 77404 433664 78279 433666
rect 77404 433608 78218 433664
rect 78274 433608 78279 433664
rect 77404 433606 78279 433608
rect 77404 433604 77410 433606
rect 78213 433603 78279 433606
rect 78622 433604 78628 433668
rect 78692 433666 78698 433668
rect 78949 433666 79015 433669
rect 78692 433664 79015 433666
rect 78692 433608 78954 433664
rect 79010 433608 79015 433664
rect 78692 433606 79015 433608
rect 78692 433604 78698 433606
rect 78949 433603 79015 433606
rect 83089 433666 83155 433669
rect 83590 433666 83596 433668
rect 83089 433664 83596 433666
rect 83089 433608 83094 433664
rect 83150 433608 83596 433664
rect 83089 433606 83596 433608
rect 83089 433603 83155 433606
rect 83590 433604 83596 433606
rect 83660 433604 83666 433668
rect 84142 433604 84148 433668
rect 84212 433666 84218 433668
rect 84469 433666 84535 433669
rect 84212 433664 84535 433666
rect 84212 433608 84474 433664
rect 84530 433608 84535 433664
rect 84212 433606 84535 433608
rect 84212 433604 84218 433606
rect 84469 433603 84535 433606
rect 85246 433604 85252 433668
rect 85316 433666 85322 433668
rect 85665 433666 85731 433669
rect 85316 433664 85731 433666
rect 85316 433608 85670 433664
rect 85726 433608 85731 433664
rect 85316 433606 85731 433608
rect 85316 433604 85322 433606
rect 85665 433603 85731 433606
rect 85798 433604 85804 433668
rect 85868 433666 85874 433668
rect 85941 433666 86007 433669
rect 87137 433668 87203 433669
rect 85868 433664 86007 433666
rect 85868 433608 85946 433664
rect 86002 433608 86007 433664
rect 85868 433606 86007 433608
rect 85868 433604 85874 433606
rect 85941 433603 86007 433606
rect 87086 433604 87092 433668
rect 87156 433666 87203 433668
rect 87156 433664 87248 433666
rect 87198 433608 87248 433664
rect 87156 433606 87248 433608
rect 87156 433604 87203 433606
rect 87454 433604 87460 433668
rect 87524 433666 87530 433668
rect 87965 433666 88031 433669
rect 87524 433664 88031 433666
rect 87524 433608 87970 433664
rect 88026 433608 88031 433664
rect 87524 433606 88031 433608
rect 87524 433604 87530 433606
rect 87137 433603 87203 433604
rect 87965 433603 88031 433606
rect 89846 433604 89852 433668
rect 89916 433666 89922 433668
rect 89989 433666 90055 433669
rect 89916 433664 90055 433666
rect 89916 433608 89994 433664
rect 90050 433608 90055 433664
rect 89916 433606 90055 433608
rect 89916 433604 89922 433606
rect 89989 433603 90055 433606
rect 91369 433666 91435 433669
rect 91502 433666 91508 433668
rect 91369 433664 91508 433666
rect 91369 433608 91374 433664
rect 91430 433608 91508 433664
rect 91369 433606 91508 433608
rect 91369 433603 91435 433606
rect 91502 433604 91508 433606
rect 91572 433604 91578 433668
rect 98310 433604 98316 433668
rect 98380 433666 98386 433668
rect 98453 433666 98519 433669
rect 99925 433668 99991 433669
rect 99925 433666 99972 433668
rect 98380 433664 98519 433666
rect 98380 433608 98458 433664
rect 98514 433608 98519 433664
rect 98380 433606 98519 433608
rect 99880 433664 99972 433666
rect 99880 433608 99930 433664
rect 99880 433606 99972 433608
rect 98380 433604 98386 433606
rect 98453 433603 98519 433606
rect 99925 433604 99972 433606
rect 100036 433604 100042 433668
rect 100886 433604 100892 433668
rect 100956 433666 100962 433668
rect 101213 433666 101279 433669
rect 100956 433664 101279 433666
rect 100956 433608 101218 433664
rect 101274 433608 101279 433664
rect 100956 433606 101279 433608
rect 100956 433604 100962 433606
rect 99925 433603 99991 433604
rect 101213 433603 101279 433606
rect 102174 433604 102180 433668
rect 102244 433666 102250 433668
rect 102685 433666 102751 433669
rect 104157 433668 104223 433669
rect 104157 433666 104204 433668
rect 102244 433664 102751 433666
rect 102244 433608 102690 433664
rect 102746 433608 102751 433664
rect 102244 433606 102751 433608
rect 104112 433664 104204 433666
rect 104112 433608 104162 433664
rect 104112 433606 104204 433608
rect 102244 433604 102250 433606
rect 102685 433603 102751 433606
rect 104157 433604 104204 433606
rect 104268 433604 104274 433668
rect 105118 433604 105124 433668
rect 105188 433666 105194 433668
rect 105445 433666 105511 433669
rect 105188 433664 105511 433666
rect 105188 433608 105450 433664
rect 105506 433608 105511 433664
rect 105188 433606 105511 433608
rect 105188 433604 105194 433606
rect 104157 433603 104223 433604
rect 105445 433603 105511 433606
rect 106406 433604 106412 433668
rect 106476 433666 106482 433668
rect 106733 433666 106799 433669
rect 106476 433664 106799 433666
rect 106476 433608 106738 433664
rect 106794 433608 106799 433664
rect 106476 433606 106799 433608
rect 106476 433604 106482 433606
rect 106733 433603 106799 433606
rect 110638 433604 110644 433668
rect 110708 433666 110714 433668
rect 110873 433666 110939 433669
rect 110708 433664 110939 433666
rect 110708 433608 110878 433664
rect 110934 433608 110939 433664
rect 110708 433606 110939 433608
rect 110708 433604 110714 433606
rect 110873 433603 110939 433606
rect 111885 433668 111951 433669
rect 111885 433664 111932 433668
rect 111996 433666 112002 433668
rect 111885 433608 111890 433664
rect 111885 433604 111932 433608
rect 111996 433606 112042 433666
rect 111996 433604 112002 433606
rect 111885 433603 111951 433604
rect 54937 433528 64890 433530
rect 54937 433472 54942 433528
rect 54998 433472 64890 433528
rect 54937 433470 64890 433472
rect 54937 433467 55003 433470
rect 66253 433394 66319 433397
rect 66253 433392 68908 433394
rect 66253 433336 66258 433392
rect 66314 433336 68908 433392
rect 112118 433364 112178 433742
rect 66253 433334 68908 433336
rect 66253 433331 66319 433334
rect 61929 432850 61995 432853
rect 68645 432850 68711 432853
rect 61929 432848 68711 432850
rect 61929 432792 61934 432848
rect 61990 432792 68650 432848
rect 68706 432792 68711 432848
rect 61929 432790 68711 432792
rect 61929 432787 61995 432790
rect 68645 432787 68711 432790
rect 112110 432788 112116 432852
rect 112180 432788 112186 432852
rect 66437 432578 66503 432581
rect 66437 432576 68908 432578
rect 66437 432520 66442 432576
rect 66498 432520 68908 432576
rect 66437 432518 68908 432520
rect 66437 432515 66503 432518
rect 112118 432306 112178 432788
rect 115565 432306 115631 432309
rect 112118 432304 115631 432306
rect 112118 432276 115570 432304
rect 112148 432248 115570 432276
rect 115626 432248 115631 432304
rect 112148 432246 115631 432248
rect 115565 432243 115631 432246
rect 583201 431626 583267 431629
rect 583520 431626 584960 431716
rect 583201 431624 584960 431626
rect 583201 431568 583206 431624
rect 583262 431568 584960 431624
rect 583201 431566 584960 431568
rect 583201 431563 583267 431566
rect 66713 431490 66779 431493
rect 66713 431488 68908 431490
rect 66713 431432 66718 431488
rect 66774 431432 68908 431488
rect 583520 431476 584960 431566
rect 66713 431430 68908 431432
rect 66713 431427 66779 431430
rect 113265 431218 113331 431221
rect 115841 431218 115907 431221
rect 112700 431216 115907 431218
rect 112700 431160 113270 431216
rect 113326 431160 115846 431216
rect 115902 431160 115907 431216
rect 112700 431158 115907 431160
rect 113265 431155 113331 431158
rect 115841 431155 115907 431158
rect 66713 430402 66779 430405
rect 66713 430400 68908 430402
rect 66713 430344 66718 430400
rect 66774 430344 68908 430400
rect 66713 430342 68908 430344
rect 66713 430339 66779 430342
rect 113817 430130 113883 430133
rect 112700 430128 113883 430130
rect 112700 430072 113822 430128
rect 113878 430072 113883 430128
rect 112700 430070 113883 430072
rect 113817 430067 113883 430070
rect 66069 429314 66135 429317
rect 115749 429314 115815 429317
rect 66069 429312 68908 429314
rect 66069 429256 66074 429312
rect 66130 429256 68908 429312
rect 66069 429254 68908 429256
rect 112700 429312 115815 429314
rect 112700 429256 115754 429312
rect 115810 429256 115815 429312
rect 112700 429254 115815 429256
rect 66069 429251 66135 429254
rect 115749 429251 115815 429254
rect 66713 428226 66779 428229
rect 115841 428226 115907 428229
rect 66713 428224 68908 428226
rect 66713 428168 66718 428224
rect 66774 428168 68908 428224
rect 66713 428166 68908 428168
rect 112700 428224 115907 428226
rect 112700 428168 115846 428224
rect 115902 428168 115907 428224
rect 112700 428166 115907 428168
rect 66713 428163 66779 428166
rect 115841 428163 115907 428166
rect 66713 427410 66779 427413
rect 66713 427408 68908 427410
rect 66713 427352 66718 427408
rect 66774 427352 68908 427408
rect 66713 427350 68908 427352
rect 66713 427347 66779 427350
rect 113265 427138 113331 427141
rect 112700 427136 113331 427138
rect 112700 427080 113270 427136
rect 113326 427080 113331 427136
rect 112700 427078 113331 427080
rect 113265 427075 113331 427078
rect 68878 425642 68938 426292
rect 115841 426050 115907 426053
rect 112700 426048 115907 426050
rect 112700 425992 115846 426048
rect 115902 425992 115907 426048
rect 112700 425990 115907 425992
rect 115841 425987 115907 425990
rect 64830 425582 68938 425642
rect 64638 425172 64644 425236
rect 64708 425234 64714 425236
rect 64830 425234 64890 425582
rect 64708 425174 64890 425234
rect 66529 425234 66595 425237
rect 66529 425232 68908 425234
rect 66529 425176 66534 425232
rect 66590 425176 68908 425232
rect 66529 425174 68908 425176
rect 64708 425172 64714 425174
rect 66529 425171 66595 425174
rect 113357 424962 113423 424965
rect 115749 424962 115815 424965
rect 112700 424960 115815 424962
rect 112700 424904 113362 424960
rect 113418 424904 115754 424960
rect 115810 424904 115815 424960
rect 112700 424902 115815 424904
rect 113357 424899 113423 424902
rect 115749 424899 115815 424902
rect 66713 424146 66779 424149
rect 114645 424146 114711 424149
rect 115841 424146 115907 424149
rect 66713 424144 68908 424146
rect 66713 424088 66718 424144
rect 66774 424088 68908 424144
rect 66713 424086 68908 424088
rect 112700 424144 115907 424146
rect 112700 424088 114650 424144
rect 114706 424088 115846 424144
rect 115902 424088 115907 424144
rect 112700 424086 115907 424088
rect 66713 424083 66779 424086
rect 114645 424083 114711 424086
rect 115841 424083 115907 424086
rect -960 423602 480 423692
rect 2773 423602 2839 423605
rect -960 423600 2839 423602
rect -960 423544 2778 423600
rect 2834 423544 2839 423600
rect -960 423542 2839 423544
rect -960 423452 480 423542
rect 2773 423539 2839 423542
rect 66713 423330 66779 423333
rect 66713 423328 68908 423330
rect 66713 423272 66718 423328
rect 66774 423272 68908 423328
rect 66713 423270 68908 423272
rect 66713 423267 66779 423270
rect 115841 423058 115907 423061
rect 112700 423056 115907 423058
rect 112700 423000 115846 423056
rect 115902 423000 115907 423056
rect 112700 422998 115907 423000
rect 115841 422995 115907 422998
rect 66846 422180 66852 422244
rect 66916 422242 66922 422244
rect 66916 422182 68908 422242
rect 66916 422180 66922 422182
rect 114553 421970 114619 421973
rect 112700 421968 114619 421970
rect 112700 421912 114558 421968
rect 114614 421912 114619 421968
rect 112700 421910 114619 421912
rect 114553 421907 114619 421910
rect 66989 421154 67055 421157
rect 66989 421152 68908 421154
rect 66989 421096 66994 421152
rect 67050 421096 68908 421152
rect 66989 421094 68908 421096
rect 66989 421091 67055 421094
rect 63401 420882 63467 420885
rect 66846 420882 66852 420884
rect 63401 420880 66852 420882
rect 63401 420824 63406 420880
rect 63462 420824 66852 420880
rect 63401 420822 66852 420824
rect 63401 420819 63467 420822
rect 66846 420820 66852 420822
rect 66916 420820 66922 420884
rect 115749 420882 115815 420885
rect 112700 420880 115815 420882
rect 112700 420824 115754 420880
rect 115810 420824 115815 420880
rect 112700 420822 115815 420824
rect 115749 420819 115815 420822
rect 66897 420066 66963 420069
rect 113173 420066 113239 420069
rect 66897 420064 68908 420066
rect 66897 420008 66902 420064
rect 66958 420008 68908 420064
rect 66897 420006 68908 420008
rect 112700 420064 113239 420066
rect 112700 420008 113178 420064
rect 113234 420008 113239 420064
rect 112700 420006 113239 420008
rect 66897 420003 66963 420006
rect 113173 420003 113239 420006
rect 66621 418978 66687 418981
rect 114645 418978 114711 418981
rect 66621 418976 68908 418978
rect 66621 418920 66626 418976
rect 66682 418920 68908 418976
rect 66621 418918 68908 418920
rect 112700 418976 114711 418978
rect 112700 418920 114650 418976
rect 114706 418920 114711 418976
rect 112700 418918 114711 418920
rect 66621 418915 66687 418918
rect 114645 418915 114711 418918
rect 583385 418298 583451 418301
rect 583520 418298 584960 418388
rect 583385 418296 584960 418298
rect 583385 418240 583390 418296
rect 583446 418240 584960 418296
rect 583385 418238 584960 418240
rect 583385 418235 583451 418238
rect 66989 418162 67055 418165
rect 67357 418162 67423 418165
rect 66989 418160 68908 418162
rect 66989 418104 66994 418160
rect 67050 418104 67362 418160
rect 67418 418104 68908 418160
rect 583520 418148 584960 418238
rect 66989 418102 68908 418104
rect 66989 418099 67055 418102
rect 67357 418099 67423 418102
rect 114502 417890 114508 417892
rect 112700 417830 114508 417890
rect 114502 417828 114508 417830
rect 114572 417828 114578 417892
rect 66897 417074 66963 417077
rect 66897 417072 68908 417074
rect 66897 417016 66902 417072
rect 66958 417016 68908 417072
rect 66897 417014 68908 417016
rect 66897 417011 66963 417014
rect 113449 416802 113515 416805
rect 115841 416802 115907 416805
rect 112700 416800 115907 416802
rect 112700 416744 113454 416800
rect 113510 416744 115846 416800
rect 115902 416744 115907 416800
rect 112700 416742 115907 416744
rect 113449 416739 113515 416742
rect 115841 416739 115907 416742
rect 66110 415924 66116 415988
rect 66180 415986 66186 415988
rect 66621 415986 66687 415989
rect 66180 415984 68908 415986
rect 66180 415928 66626 415984
rect 66682 415928 68908 415984
rect 66180 415926 68908 415928
rect 66180 415924 66186 415926
rect 66621 415923 66687 415926
rect 115841 415714 115907 415717
rect 112700 415712 115907 415714
rect 112700 415656 115846 415712
rect 115902 415656 115907 415712
rect 112700 415654 115907 415656
rect 115841 415651 115907 415654
rect 66713 414898 66779 414901
rect 115841 414898 115907 414901
rect 66713 414896 68908 414898
rect 66713 414840 66718 414896
rect 66774 414840 68908 414896
rect 66713 414838 68908 414840
rect 112700 414896 115907 414898
rect 112700 414840 115846 414896
rect 115902 414840 115907 414896
rect 112700 414838 115907 414840
rect 66713 414835 66779 414838
rect 115841 414835 115907 414838
rect 66897 414082 66963 414085
rect 66897 414080 68908 414082
rect 66897 414024 66902 414080
rect 66958 414024 68908 414080
rect 66897 414022 68908 414024
rect 66897 414019 66963 414022
rect 115841 413810 115907 413813
rect 112700 413808 115907 413810
rect 112700 413752 115846 413808
rect 115902 413752 115907 413808
rect 112700 413750 115907 413752
rect 115841 413747 115907 413750
rect 66897 412994 66963 412997
rect 66897 412992 68908 412994
rect 66897 412936 66902 412992
rect 66958 412936 68908 412992
rect 66897 412934 68908 412936
rect 66897 412931 66963 412934
rect 115105 412722 115171 412725
rect 112700 412720 115171 412722
rect 112700 412664 115110 412720
rect 115166 412664 115171 412720
rect 112700 412662 115171 412664
rect 115105 412659 115171 412662
rect 66713 411906 66779 411909
rect 66713 411904 68908 411906
rect 66713 411848 66718 411904
rect 66774 411848 68908 411904
rect 66713 411846 68908 411848
rect 66713 411843 66779 411846
rect 115197 411634 115263 411637
rect 112700 411632 115263 411634
rect 112700 411576 115202 411632
rect 115258 411576 115263 411632
rect 112700 411574 115263 411576
rect 115197 411571 115263 411574
rect 66897 410818 66963 410821
rect 66897 410816 68908 410818
rect 66897 410760 66902 410816
rect 66958 410760 68908 410816
rect 66897 410758 68908 410760
rect 66897 410755 66963 410758
rect -960 410546 480 410636
rect 2865 410546 2931 410549
rect 115841 410546 115907 410549
rect -960 410544 2931 410546
rect -960 410488 2870 410544
rect 2926 410488 2931 410544
rect -960 410486 2931 410488
rect 112700 410544 115907 410546
rect 112700 410488 115846 410544
rect 115902 410488 115907 410544
rect 112700 410486 115907 410488
rect -960 410396 480 410486
rect 2865 410483 2931 410486
rect 115841 410483 115907 410486
rect 66662 409668 66668 409732
rect 66732 409730 66738 409732
rect 67766 409730 67772 409732
rect 66732 409670 67772 409730
rect 66732 409668 66738 409670
rect 67766 409668 67772 409670
rect 67836 409730 67842 409732
rect 115841 409730 115907 409733
rect 67836 409670 68908 409730
rect 112700 409728 115907 409730
rect 112700 409672 115846 409728
rect 115902 409672 115907 409728
rect 112700 409670 115907 409672
rect 67836 409668 67842 409670
rect 115841 409667 115907 409670
rect 66253 408914 66319 408917
rect 66253 408912 68908 408914
rect 66253 408856 66258 408912
rect 66314 408856 68908 408912
rect 66253 408854 68908 408856
rect 66253 408851 66319 408854
rect 114686 408642 114692 408644
rect 112700 408582 114692 408642
rect 114686 408580 114692 408582
rect 114756 408580 114762 408644
rect 66897 407826 66963 407829
rect 66897 407824 68908 407826
rect 66897 407768 66902 407824
rect 66958 407768 68908 407824
rect 66897 407766 68908 407768
rect 66897 407763 66963 407766
rect 115013 407554 115079 407557
rect 112700 407552 115079 407554
rect 112700 407496 115018 407552
rect 115074 407496 115079 407552
rect 112700 407494 115079 407496
rect 115013 407491 115079 407494
rect 66437 406738 66503 406741
rect 66437 406736 68908 406738
rect 66437 406680 66442 406736
rect 66498 406680 68908 406736
rect 66437 406678 68908 406680
rect 66437 406675 66503 406678
rect 112670 405925 112730 406436
rect 112670 405920 112779 405925
rect 112670 405864 112718 405920
rect 112774 405864 112779 405920
rect 112670 405862 112779 405864
rect 112713 405859 112779 405862
rect 67449 405650 67515 405653
rect 115841 405650 115907 405653
rect 67449 405648 68908 405650
rect 67449 405592 67454 405648
rect 67510 405592 68908 405648
rect 67449 405590 68908 405592
rect 112700 405648 115907 405650
rect 112700 405592 115846 405648
rect 115902 405592 115907 405648
rect 112700 405590 115907 405592
rect 67449 405587 67515 405590
rect 115841 405587 115907 405590
rect 583293 404970 583359 404973
rect 583520 404970 584960 405060
rect 583293 404968 584960 404970
rect 583293 404912 583298 404968
rect 583354 404912 584960 404968
rect 583293 404910 584960 404912
rect 583293 404907 583359 404910
rect 583520 404820 584960 404910
rect 66897 404562 66963 404565
rect 115841 404562 115907 404565
rect 66897 404560 68908 404562
rect 66897 404504 66902 404560
rect 66958 404504 68908 404560
rect 66897 404502 68908 404504
rect 112700 404560 115907 404562
rect 112700 404504 115846 404560
rect 115902 404504 115907 404560
rect 112700 404502 115907 404504
rect 66897 404499 66963 404502
rect 115841 404499 115907 404502
rect 65977 403746 66043 403749
rect 65977 403744 68908 403746
rect 65977 403688 65982 403744
rect 66038 403688 68908 403744
rect 65977 403686 68908 403688
rect 65977 403683 66043 403686
rect 115841 403474 115907 403477
rect 112700 403472 115907 403474
rect 112700 403416 115846 403472
rect 115902 403416 115907 403472
rect 112700 403414 115907 403416
rect 115841 403411 115907 403414
rect 66713 402658 66779 402661
rect 66713 402656 68908 402658
rect 66713 402600 66718 402656
rect 66774 402600 68908 402656
rect 66713 402598 68908 402600
rect 66713 402595 66779 402598
rect 115841 402386 115907 402389
rect 112700 402384 115907 402386
rect 112700 402328 115846 402384
rect 115902 402328 115907 402384
rect 112700 402326 115907 402328
rect 115841 402323 115907 402326
rect 66897 401570 66963 401573
rect 66897 401568 68908 401570
rect 66897 401512 66902 401568
rect 66958 401512 68908 401568
rect 66897 401510 68908 401512
rect 66897 401507 66963 401510
rect 115197 401298 115263 401301
rect 112700 401296 115263 401298
rect 112700 401240 115202 401296
rect 115258 401240 115263 401296
rect 112700 401238 115263 401240
rect 115197 401235 115263 401238
rect 66805 400482 66871 400485
rect 115841 400482 115907 400485
rect 66805 400480 68908 400482
rect 66805 400424 66810 400480
rect 66866 400424 68908 400480
rect 66805 400422 68908 400424
rect 112700 400480 115907 400482
rect 112700 400424 115846 400480
rect 115902 400424 115907 400480
rect 112700 400422 115907 400424
rect 66805 400419 66871 400422
rect 115841 400419 115907 400422
rect 66529 399666 66595 399669
rect 66529 399664 68908 399666
rect 66529 399608 66534 399664
rect 66590 399608 68908 399664
rect 66529 399606 68908 399608
rect 66529 399603 66595 399606
rect 114318 399468 114324 399532
rect 114388 399530 114394 399532
rect 114553 399530 114619 399533
rect 114388 399528 114619 399530
rect 114388 399472 114558 399528
rect 114614 399472 114619 399528
rect 114388 399470 114619 399472
rect 114388 399468 114394 399470
rect 114553 399467 114619 399470
rect 115381 399394 115447 399397
rect 112700 399392 115447 399394
rect 112700 399336 115386 399392
rect 115442 399336 115447 399392
rect 112700 399334 115447 399336
rect 115381 399331 115447 399334
rect 114553 398850 114619 398853
rect 140773 398850 140839 398853
rect 114553 398848 140839 398850
rect 114553 398792 114558 398848
rect 114614 398792 140778 398848
rect 140834 398792 140839 398848
rect 114553 398790 140839 398792
rect 114553 398787 114619 398790
rect 140773 398787 140839 398790
rect 66621 398578 66687 398581
rect 66621 398576 68908 398578
rect 66621 398520 66626 398576
rect 66682 398520 68908 398576
rect 66621 398518 68908 398520
rect 66621 398515 66687 398518
rect 115565 398306 115631 398309
rect 112700 398304 115631 398306
rect 112700 398248 115570 398304
rect 115626 398248 115631 398304
rect 112700 398246 115631 398248
rect 115565 398243 115631 398246
rect 67725 397898 67791 397901
rect 67725 397896 68938 397898
rect 67725 397840 67730 397896
rect 67786 397840 68938 397896
rect 67725 397838 68938 397840
rect 67725 397835 67791 397838
rect -960 397490 480 397580
rect 3509 397490 3575 397493
rect -960 397488 3575 397490
rect -960 397432 3514 397488
rect 3570 397432 3575 397488
rect 68878 397460 68938 397838
rect -960 397430 3575 397432
rect -960 397340 480 397430
rect 3509 397427 3575 397430
rect 115841 397218 115907 397221
rect 112700 397216 115907 397218
rect 112700 397160 115846 397216
rect 115902 397160 115907 397216
rect 112700 397158 115907 397160
rect 115841 397155 115907 397158
rect 67081 396402 67147 396405
rect 67449 396402 67515 396405
rect 114553 396402 114619 396405
rect 67081 396400 68908 396402
rect 67081 396344 67086 396400
rect 67142 396344 67454 396400
rect 67510 396344 68908 396400
rect 67081 396342 68908 396344
rect 112700 396400 114619 396402
rect 112700 396344 114558 396400
rect 114614 396344 114619 396400
rect 112700 396342 114619 396344
rect 67081 396339 67147 396342
rect 67449 396339 67515 396342
rect 114553 396339 114619 396342
rect 66805 395314 66871 395317
rect 115841 395314 115907 395317
rect 66805 395312 68908 395314
rect 66805 395256 66810 395312
rect 66866 395256 68908 395312
rect 66805 395254 68908 395256
rect 112700 395312 115907 395314
rect 112700 395256 115846 395312
rect 115902 395256 115907 395312
rect 112700 395254 115907 395256
rect 66805 395251 66871 395254
rect 115841 395251 115907 395254
rect 66161 394634 66227 394637
rect 68134 394634 68140 394636
rect 66161 394632 68140 394634
rect 66161 394576 66166 394632
rect 66222 394576 68140 394632
rect 66161 394574 68140 394576
rect 66161 394571 66227 394574
rect 68134 394572 68140 394574
rect 68204 394572 68210 394636
rect 66345 394498 66411 394501
rect 66345 394496 68908 394498
rect 66345 394440 66350 394496
rect 66406 394440 68908 394496
rect 66345 394438 68908 394440
rect 66345 394435 66411 394438
rect 115381 394226 115447 394229
rect 112700 394224 115447 394226
rect 112700 394168 115386 394224
rect 115442 394168 115447 394224
rect 112700 394166 115447 394168
rect 115381 394163 115447 394166
rect 66805 393410 66871 393413
rect 66805 393408 68908 393410
rect 66805 393352 66810 393408
rect 66866 393352 68908 393408
rect 66805 393350 68908 393352
rect 66805 393347 66871 393350
rect 115841 393138 115907 393141
rect 112700 393136 115907 393138
rect 112700 393080 115846 393136
rect 115902 393080 115907 393136
rect 112700 393078 115907 393080
rect 115841 393075 115907 393078
rect 66805 392322 66871 392325
rect 66805 392320 68908 392322
rect 66805 392264 66810 392320
rect 66866 392264 68908 392320
rect 66805 392262 68908 392264
rect 66805 392259 66871 392262
rect 114553 392050 114619 392053
rect 112700 392048 114619 392050
rect 112700 391992 114558 392048
rect 114614 391992 114619 392048
rect 112700 391990 114619 391992
rect 114553 391987 114619 391990
rect 583520 391628 584960 391868
rect 53465 391506 53531 391509
rect 53465 391504 99390 391506
rect 53465 391448 53470 391504
rect 53526 391448 99390 391504
rect 53465 391446 99390 391448
rect 53465 391443 53531 391446
rect 66805 391234 66871 391237
rect 66805 391232 68908 391234
rect 66805 391176 66810 391232
rect 66866 391176 68908 391232
rect 66805 391174 68908 391176
rect 66805 391171 66871 391174
rect 84377 390690 84443 390693
rect 85246 390690 85252 390692
rect 84377 390688 85252 390690
rect 84377 390632 84382 390688
rect 84438 390632 85252 390688
rect 84377 390630 85252 390632
rect 84377 390627 84443 390630
rect 85246 390628 85252 390630
rect 85316 390628 85322 390692
rect 99330 390690 99390 391446
rect 115013 391234 115079 391237
rect 112700 391232 115079 391234
rect 112700 391176 115018 391232
rect 115074 391176 115079 391232
rect 112700 391174 115079 391176
rect 115013 391171 115079 391174
rect 102409 390962 102475 390965
rect 103278 390962 103284 390964
rect 102409 390960 103284 390962
rect 102409 390904 102414 390960
rect 102470 390904 103284 390960
rect 102409 390902 103284 390904
rect 102409 390899 102475 390902
rect 103278 390900 103284 390902
rect 103348 390900 103354 390964
rect 106222 390900 106228 390964
rect 106292 390962 106298 390964
rect 106733 390962 106799 390965
rect 106292 390960 106799 390962
rect 106292 390904 106738 390960
rect 106794 390904 106799 390960
rect 106292 390902 106799 390904
rect 106292 390900 106298 390902
rect 106733 390899 106799 390902
rect 103881 390690 103947 390693
rect 99330 390688 103947 390690
rect 99330 390632 103886 390688
rect 103942 390632 103947 390688
rect 99330 390630 103947 390632
rect 72325 390420 72391 390421
rect 72325 390416 72372 390420
rect 72436 390418 72442 390420
rect 72325 390360 72330 390416
rect 72325 390356 72372 390360
rect 72436 390358 72482 390418
rect 72436 390356 72442 390358
rect 73470 390356 73476 390420
rect 73540 390418 73546 390420
rect 73981 390418 74047 390421
rect 77201 390420 77267 390421
rect 77150 390418 77156 390420
rect 73540 390416 74047 390418
rect 73540 390360 73986 390416
rect 74042 390360 74047 390416
rect 73540 390358 74047 390360
rect 77110 390358 77156 390418
rect 77220 390416 77267 390420
rect 77262 390360 77267 390416
rect 73540 390356 73546 390358
rect 72325 390355 72391 390356
rect 73981 390355 74047 390358
rect 77150 390356 77156 390358
rect 77220 390356 77267 390360
rect 77201 390355 77267 390356
rect 79409 390418 79475 390421
rect 81985 390420 82051 390421
rect 79910 390418 79916 390420
rect 79409 390416 79916 390418
rect 79409 390360 79414 390416
rect 79470 390360 79916 390416
rect 79409 390358 79916 390360
rect 79409 390355 79475 390358
rect 79910 390356 79916 390358
rect 79980 390356 79986 390420
rect 81934 390418 81940 390420
rect 81894 390358 81940 390418
rect 82004 390416 82051 390420
rect 82046 390360 82051 390416
rect 81934 390356 81940 390358
rect 82004 390356 82051 390360
rect 81985 390355 82051 390356
rect 100342 390285 100402 390630
rect 103881 390627 103947 390630
rect 107745 390556 107811 390557
rect 107694 390492 107700 390556
rect 107764 390554 107811 390556
rect 107764 390552 107856 390554
rect 107806 390496 107856 390552
rect 107764 390494 107856 390496
rect 107764 390492 107811 390494
rect 107745 390491 107811 390492
rect 111701 390420 111767 390421
rect 111701 390416 111748 390420
rect 111812 390418 111818 390420
rect 111701 390360 111706 390416
rect 111701 390356 111748 390360
rect 111812 390358 111858 390418
rect 111812 390356 111818 390358
rect 111701 390355 111767 390356
rect 100293 390280 100402 390285
rect 100293 390224 100298 390280
rect 100354 390224 100402 390280
rect 100293 390222 100402 390224
rect 107653 390282 107719 390285
rect 108614 390282 108620 390284
rect 107653 390280 108620 390282
rect 107653 390224 107658 390280
rect 107714 390224 108620 390280
rect 107653 390222 108620 390224
rect 100293 390219 100359 390222
rect 107653 390219 107719 390222
rect 108614 390220 108620 390222
rect 108684 390220 108690 390284
rect 95325 389602 95391 389605
rect 96286 389602 96292 389604
rect 95325 389600 96292 389602
rect 95325 389544 95330 389600
rect 95386 389544 96292 389600
rect 95325 389542 96292 389544
rect 95325 389539 95391 389542
rect 96286 389540 96292 389542
rect 96356 389540 96362 389604
rect 51717 389194 51783 389197
rect 107745 389194 107811 389197
rect 51717 389192 107811 389194
rect 51717 389136 51722 389192
rect 51778 389136 107750 389192
rect 107806 389136 107811 389192
rect 51717 389134 107811 389136
rect 51717 389131 51783 389134
rect 107745 389131 107811 389134
rect 71446 388996 71452 389060
rect 71516 389058 71522 389060
rect 71773 389058 71839 389061
rect 72509 389058 72575 389061
rect 71516 389056 72575 389058
rect 71516 389000 71778 389056
rect 71834 389000 72514 389056
rect 72570 389000 72575 389056
rect 71516 388998 72575 389000
rect 71516 388996 71522 388998
rect 71773 388995 71839 388998
rect 72509 388995 72575 388998
rect 76005 389058 76071 389061
rect 76741 389058 76807 389061
rect 78857 389060 78923 389061
rect 76005 389056 76807 389058
rect 76005 389000 76010 389056
rect 76066 389000 76746 389056
rect 76802 389000 76807 389056
rect 76005 388998 76807 389000
rect 76005 388995 76071 388998
rect 76741 388995 76807 388998
rect 78806 388996 78812 389060
rect 78876 389058 78923 389060
rect 80053 389060 80119 389061
rect 80053 389058 80100 389060
rect 78876 389056 78968 389058
rect 78918 389000 78968 389056
rect 78876 388998 78968 389000
rect 79972 389056 80100 389058
rect 80164 389058 80170 389060
rect 80973 389058 81039 389061
rect 80164 389056 81039 389058
rect 79972 389000 80058 389056
rect 80164 389000 80978 389056
rect 81034 389000 81039 389056
rect 79972 388998 80100 389000
rect 78876 388996 78923 388998
rect 78857 388995 78923 388996
rect 80053 388996 80100 388998
rect 80164 388998 81039 389000
rect 80164 388996 80170 388998
rect 80053 388995 80119 388996
rect 80973 388995 81039 388998
rect 88333 389058 88399 389061
rect 88742 389058 88748 389060
rect 88333 389056 88748 389058
rect 88333 389000 88338 389056
rect 88394 389000 88748 389056
rect 88333 388998 88748 389000
rect 88333 388995 88399 388998
rect 88742 388996 88748 388998
rect 88812 389058 88818 389060
rect 89253 389058 89319 389061
rect 88812 389056 89319 389058
rect 88812 389000 89258 389056
rect 89314 389000 89319 389056
rect 88812 388998 89319 389000
rect 88812 388996 88818 388998
rect 89253 388995 89319 388998
rect 99649 389058 99715 389061
rect 100150 389058 100156 389060
rect 99649 389056 100156 389058
rect 99649 389000 99654 389056
rect 99710 389000 100156 389056
rect 99649 388998 100156 389000
rect 99649 388995 99715 388998
rect 100150 388996 100156 388998
rect 100220 389058 100226 389060
rect 100477 389058 100543 389061
rect 100753 389060 100819 389061
rect 100220 389056 100543 389058
rect 100220 389000 100482 389056
rect 100538 389000 100543 389056
rect 100220 388998 100543 389000
rect 100220 388996 100226 388998
rect 100477 388995 100543 388998
rect 100702 388996 100708 389060
rect 100772 389058 100819 389060
rect 100772 389056 100864 389058
rect 100814 389000 100864 389056
rect 100772 388998 100864 389000
rect 100772 388996 100819 388998
rect 104934 388996 104940 389060
rect 105004 389058 105010 389060
rect 105261 389058 105327 389061
rect 105004 389056 105327 389058
rect 105004 389000 105266 389056
rect 105322 389000 105327 389056
rect 105004 388998 105327 389000
rect 105004 388996 105010 388998
rect 100753 388995 100819 388996
rect 105261 388995 105327 388998
rect 124765 389058 124831 389061
rect 125726 389058 125732 389060
rect 124765 389056 125732 389058
rect 124765 389000 124770 389056
rect 124826 389000 125732 389056
rect 124765 388998 125732 389000
rect 124765 388995 124831 388998
rect 125726 388996 125732 388998
rect 125796 388996 125802 389060
rect 57094 388860 57100 388924
rect 57164 388922 57170 388924
rect 71865 388922 71931 388925
rect 57164 388920 71931 388922
rect 57164 388864 71870 388920
rect 71926 388864 71931 388920
rect 57164 388862 71931 388864
rect 57164 388860 57170 388862
rect 71865 388859 71931 388862
rect 14457 388786 14523 388789
rect 81433 388786 81499 388789
rect 14457 388784 81499 388786
rect 14457 388728 14462 388784
rect 14518 388728 81438 388784
rect 81494 388728 81499 388784
rect 14457 388726 81499 388728
rect 14457 388723 14523 388726
rect 81433 388723 81499 388726
rect 77293 387970 77359 387973
rect 78438 387970 78444 387972
rect 77293 387968 78444 387970
rect 77293 387912 77298 387968
rect 77354 387912 78444 387968
rect 77293 387910 78444 387912
rect 77293 387907 77359 387910
rect 78438 387908 78444 387910
rect 78508 387908 78514 387972
rect 70894 387772 70900 387836
rect 70964 387834 70970 387836
rect 71221 387834 71287 387837
rect 70964 387832 71287 387834
rect 70964 387776 71226 387832
rect 71282 387776 71287 387832
rect 70964 387774 71287 387776
rect 70964 387772 70970 387774
rect 71221 387771 71287 387774
rect 91277 387834 91343 387837
rect 91502 387834 91508 387836
rect 91277 387832 91508 387834
rect 91277 387776 91282 387832
rect 91338 387776 91508 387832
rect 91277 387774 91508 387776
rect 91277 387771 91343 387774
rect 91502 387772 91508 387774
rect 91572 387772 91578 387836
rect 94405 387834 94471 387837
rect 102777 387834 102843 387837
rect 94405 387832 102843 387834
rect 94405 387776 94410 387832
rect 94466 387776 102782 387832
rect 102838 387776 102843 387832
rect 94405 387774 102843 387776
rect 94405 387771 94471 387774
rect 102777 387771 102843 387774
rect 73153 387698 73219 387701
rect 73470 387698 73476 387700
rect 73153 387696 73476 387698
rect 73153 387640 73158 387696
rect 73214 387640 73476 387696
rect 73153 387638 73476 387640
rect 73153 387635 73219 387638
rect 73470 387636 73476 387638
rect 73540 387636 73546 387700
rect 73470 387500 73476 387564
rect 73540 387562 73546 387564
rect 75269 387562 75335 387565
rect 73540 387560 75335 387562
rect 73540 387504 75274 387560
rect 75330 387504 75335 387560
rect 73540 387502 75335 387504
rect 73540 387500 73546 387502
rect 75269 387499 75335 387502
rect 92381 387018 92447 387021
rect 102174 387018 102180 387020
rect 92381 387016 102180 387018
rect 92381 386960 92386 387016
rect 92442 386960 102180 387016
rect 92381 386958 102180 386960
rect 92381 386955 92447 386958
rect 102174 386956 102180 386958
rect 102244 386956 102250 387020
rect 72918 385732 72924 385796
rect 72988 385794 72994 385796
rect 77477 385794 77543 385797
rect 72988 385792 77543 385794
rect 72988 385736 77482 385792
rect 77538 385736 77543 385792
rect 72988 385734 77543 385736
rect 72988 385732 72994 385734
rect 77477 385731 77543 385734
rect 48037 385658 48103 385661
rect 81249 385658 81315 385661
rect 48037 385656 81315 385658
rect 48037 385600 48042 385656
rect 48098 385600 81254 385656
rect 81310 385600 81315 385656
rect 48037 385598 81315 385600
rect 48037 385595 48103 385598
rect 81249 385595 81315 385598
rect 89621 385658 89687 385661
rect 97206 385658 97212 385660
rect 89621 385656 97212 385658
rect 89621 385600 89626 385656
rect 89682 385600 97212 385656
rect 89621 385598 97212 385600
rect 89621 385595 89687 385598
rect 97206 385596 97212 385598
rect 97276 385596 97282 385660
rect -960 384284 480 384524
rect 52177 384298 52243 384301
rect 78806 384298 78812 384300
rect 52177 384296 78812 384298
rect 52177 384240 52182 384296
rect 52238 384240 78812 384296
rect 52177 384238 78812 384240
rect 52177 384235 52243 384238
rect 78806 384236 78812 384238
rect 78876 384236 78882 384300
rect 93761 384298 93827 384301
rect 105118 384298 105124 384300
rect 93761 384296 105124 384298
rect 93761 384240 93766 384296
rect 93822 384240 105124 384296
rect 93761 384238 105124 384240
rect 93761 384235 93827 384238
rect 105118 384236 105124 384238
rect 105188 384236 105194 384300
rect 108246 384236 108252 384300
rect 108316 384298 108322 384300
rect 117313 384298 117379 384301
rect 108316 384296 117379 384298
rect 108316 384240 117318 384296
rect 117374 384240 117379 384296
rect 108316 384238 117379 384240
rect 108316 384236 108322 384238
rect 117313 384235 117379 384238
rect 79869 383754 79935 383757
rect 85798 383754 85804 383756
rect 79869 383752 85804 383754
rect 79869 383696 79874 383752
rect 79930 383696 85804 383752
rect 79869 383694 85804 383696
rect 79869 383691 79935 383694
rect 85798 383692 85804 383694
rect 85868 383692 85874 383756
rect 68134 383556 68140 383620
rect 68204 383618 68210 383620
rect 91369 383618 91435 383621
rect 91737 383618 91803 383621
rect 68204 383616 91803 383618
rect 68204 383560 91374 383616
rect 91430 383560 91742 383616
rect 91798 383560 91803 383616
rect 68204 383558 91803 383560
rect 68204 383556 68210 383558
rect 91369 383555 91435 383558
rect 91737 383555 91803 383558
rect 94037 382258 94103 382261
rect 94998 382258 95004 382260
rect 94037 382256 95004 382258
rect 94037 382200 94042 382256
rect 94098 382200 95004 382256
rect 94037 382198 95004 382200
rect 94037 382195 94103 382198
rect 94998 382196 95004 382198
rect 95068 382196 95074 382260
rect 95182 380972 95188 381036
rect 95252 381034 95258 381036
rect 100702 381034 100708 381036
rect 95252 380974 100708 381034
rect 95252 380972 95258 380974
rect 100702 380972 100708 380974
rect 100772 380972 100778 381036
rect 73061 380218 73127 380221
rect 78622 380218 78628 380220
rect 73061 380216 78628 380218
rect 73061 380160 73066 380216
rect 73122 380160 78628 380216
rect 73061 380158 78628 380160
rect 73061 380155 73127 380158
rect 78622 380156 78628 380158
rect 78692 380156 78698 380220
rect 86861 380218 86927 380221
rect 96838 380218 96844 380220
rect 86861 380216 96844 380218
rect 86861 380160 86866 380216
rect 86922 380160 96844 380216
rect 86861 380158 96844 380160
rect 86861 380155 86927 380158
rect 96838 380156 96844 380158
rect 96908 380156 96914 380220
rect 79317 378722 79383 378725
rect 87454 378722 87460 378724
rect 79317 378720 87460 378722
rect 79317 378664 79322 378720
rect 79378 378664 87460 378720
rect 79317 378662 87460 378664
rect 79317 378659 79383 378662
rect 87454 378660 87460 378662
rect 87524 378660 87530 378724
rect 583520 378450 584960 378540
rect 583342 378390 584960 378450
rect 583342 378314 583402 378390
rect 583520 378314 584960 378390
rect 583342 378300 584960 378314
rect 583342 378254 583586 378300
rect 583526 378181 583586 378254
rect 583477 378176 583586 378181
rect 583477 378120 583482 378176
rect 583538 378120 583586 378176
rect 583477 378118 583586 378120
rect 583477 378115 583543 378118
rect 84101 376002 84167 376005
rect 91318 376002 91324 376004
rect 84101 376000 91324 376002
rect 84101 375944 84106 376000
rect 84162 375944 91324 376000
rect 84101 375942 91324 375944
rect 84101 375939 84167 375942
rect 91318 375940 91324 375942
rect 91388 375940 91394 376004
rect 91502 375940 91508 376004
rect 91572 376002 91578 376004
rect 97165 376002 97231 376005
rect 91572 376000 97231 376002
rect 91572 375944 97170 376000
rect 97226 375944 97231 376000
rect 91572 375942 97231 375944
rect 91572 375940 91578 375942
rect 97165 375939 97231 375942
rect 97901 376002 97967 376005
rect 108982 376002 108988 376004
rect 97901 376000 108988 376002
rect 97901 375944 97906 376000
rect 97962 375944 108988 376000
rect 97901 375942 108988 375944
rect 97901 375939 97967 375942
rect 108982 375940 108988 375942
rect 109052 375940 109058 376004
rect 96521 374642 96587 374645
rect 106406 374642 106412 374644
rect 96521 374640 106412 374642
rect 96521 374584 96526 374640
rect 96582 374584 106412 374640
rect 96521 374582 106412 374584
rect 96521 374579 96587 374582
rect 106406 374580 106412 374582
rect 106476 374580 106482 374644
rect 91001 373282 91067 373285
rect 100886 373282 100892 373284
rect 91001 373280 100892 373282
rect 91001 373224 91006 373280
rect 91062 373224 100892 373280
rect 91001 373222 100892 373224
rect 91001 373219 91067 373222
rect 100886 373220 100892 373222
rect 100956 373220 100962 373284
rect -960 371378 480 371468
rect 3417 371378 3483 371381
rect -960 371376 3483 371378
rect -960 371320 3422 371376
rect 3478 371320 3483 371376
rect -960 371318 3483 371320
rect -960 371228 480 371318
rect 3417 371315 3483 371318
rect 77201 365666 77267 365669
rect 83958 365666 83964 365668
rect 77201 365664 83964 365666
rect 77201 365608 77206 365664
rect 77262 365608 83964 365664
rect 77201 365606 83964 365608
rect 77201 365603 77267 365606
rect 83958 365604 83964 365606
rect 84028 365604 84034 365668
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect 70301 364442 70367 364445
rect 74574 364442 74580 364444
rect 70301 364440 74580 364442
rect 70301 364384 70306 364440
rect 70362 364384 74580 364440
rect 70301 364382 74580 364384
rect 70301 364379 70367 364382
rect 74574 364380 74580 364382
rect 74644 364380 74650 364444
rect -960 358458 480 358548
rect 3325 358458 3391 358461
rect -960 358456 3391 358458
rect -960 358400 3330 358456
rect 3386 358400 3391 358456
rect -960 358398 3391 358400
rect -960 358308 480 358398
rect 3325 358395 3391 358398
rect 93669 353970 93735 353973
rect 104198 353970 104204 353972
rect 93669 353968 104204 353970
rect 93669 353912 93674 353968
rect 93730 353912 104204 353968
rect 93669 353910 104204 353912
rect 93669 353907 93735 353910
rect 104198 353908 104204 353910
rect 104268 353908 104274 353972
rect 88006 351868 88012 351932
rect 88076 351930 88082 351932
rect 92473 351930 92539 351933
rect 88076 351928 92539 351930
rect 88076 351872 92478 351928
rect 92534 351872 92539 351928
rect 88076 351870 92539 351872
rect 88076 351868 88082 351870
rect 92473 351867 92539 351870
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 83549 339556 83615 339557
rect 82854 339492 82860 339556
rect 82924 339554 82930 339556
rect 83549 339554 83596 339556
rect 82924 339552 83596 339554
rect 83660 339554 83666 339556
rect 82924 339496 83554 339552
rect 82924 339494 83596 339496
rect 82924 339492 82930 339494
rect 83549 339492 83596 339494
rect 83660 339494 83742 339554
rect 83660 339492 83666 339494
rect 83549 339491 83615 339492
rect 583520 338452 584960 338692
rect 115197 335474 115263 335477
rect 237966 335474 237972 335476
rect 115197 335472 237972 335474
rect 115197 335416 115202 335472
rect 115258 335416 237972 335472
rect 115197 335414 237972 335416
rect 115197 335411 115263 335414
rect 237966 335412 237972 335414
rect 238036 335412 238042 335476
rect 98126 332556 98132 332620
rect 98196 332618 98202 332620
rect 98494 332618 98500 332620
rect 98196 332558 98500 332618
rect 98196 332556 98202 332558
rect 98494 332556 98500 332558
rect 98564 332618 98570 332620
rect 99281 332618 99347 332621
rect 98564 332616 99347 332618
rect 98564 332560 99286 332616
rect 99342 332560 99347 332616
rect 98564 332558 99347 332560
rect 98564 332556 98570 332558
rect 99281 332555 99347 332558
rect -960 332196 480 332436
rect 84009 330442 84075 330445
rect 92606 330442 92612 330444
rect 84009 330440 92612 330442
rect 84009 330384 84014 330440
rect 84070 330384 92612 330440
rect 84009 330382 92612 330384
rect 84009 330379 84075 330382
rect 92606 330380 92612 330382
rect 92676 330380 92682 330444
rect 96705 330306 96771 330309
rect 97809 330306 97875 330309
rect 96705 330304 97875 330306
rect 96705 330248 96710 330304
rect 96766 330248 97814 330304
rect 97870 330248 97875 330304
rect 96705 330246 97875 330248
rect 96705 330243 96771 330246
rect 97809 330243 97875 330246
rect 97809 329898 97875 329901
rect 242014 329898 242020 329900
rect 97809 329896 242020 329898
rect 97809 329840 97814 329896
rect 97870 329840 242020 329896
rect 97809 329838 242020 329840
rect 97809 329835 97875 329838
rect 242014 329836 242020 329838
rect 242084 329836 242090 329900
rect 12341 328538 12407 328541
rect 201493 328538 201559 328541
rect 12341 328536 201559 328538
rect 12341 328480 12346 328536
rect 12402 328480 201498 328536
rect 201554 328480 201559 328536
rect 12341 328478 201559 328480
rect 12341 328475 12407 328478
rect 201493 328475 201559 328478
rect 98085 327722 98151 327725
rect 111926 327722 111932 327724
rect 98085 327720 111932 327722
rect 98085 327664 98090 327720
rect 98146 327664 111932 327720
rect 98085 327662 111932 327664
rect 98085 327659 98151 327662
rect 111926 327660 111932 327662
rect 111996 327660 112002 327724
rect 75269 327042 75335 327045
rect 82854 327042 82860 327044
rect 75269 327040 82860 327042
rect 75269 326984 75274 327040
rect 75330 326984 82860 327040
rect 75269 326982 82860 326984
rect 75269 326979 75335 326982
rect 82854 326980 82860 326982
rect 82924 326980 82930 327044
rect 89529 326362 89595 326365
rect 99966 326362 99972 326364
rect 89529 326360 99972 326362
rect 89529 326304 89534 326360
rect 89590 326304 99972 326360
rect 89529 326302 99972 326304
rect 89529 326299 89595 326302
rect 99966 326300 99972 326302
rect 100036 326300 100042 326364
rect 580901 325274 580967 325277
rect 583520 325274 584960 325364
rect 580901 325272 584960 325274
rect 580901 325216 580906 325272
rect 580962 325216 584960 325272
rect 580901 325214 584960 325216
rect 580901 325211 580967 325214
rect 583520 325124 584960 325214
rect 79409 323642 79475 323645
rect 86166 323642 86172 323644
rect 79409 323640 86172 323642
rect 79409 323584 79414 323640
rect 79470 323584 86172 323640
rect 79409 323582 86172 323584
rect 79409 323579 79475 323582
rect 86166 323580 86172 323582
rect 86236 323580 86242 323644
rect 86718 322900 86724 322964
rect 86788 322962 86794 322964
rect 90357 322962 90423 322965
rect 86788 322960 90423 322962
rect 86788 322904 90362 322960
rect 90418 322904 90423 322960
rect 86788 322902 90423 322904
rect 86788 322900 86794 322902
rect 90357 322899 90423 322902
rect 75678 321540 75684 321604
rect 75748 321602 75754 321604
rect 256049 321602 256115 321605
rect 75748 321600 256115 321602
rect 75748 321544 256054 321600
rect 256110 321544 256115 321600
rect 75748 321542 256115 321544
rect 75748 321540 75754 321542
rect 256049 321539 256115 321542
rect 90950 321404 90956 321468
rect 91020 321466 91026 321468
rect 95233 321466 95299 321469
rect 91020 321464 95299 321466
rect 91020 321408 95238 321464
rect 95294 321408 95299 321464
rect 91020 321406 95299 321408
rect 91020 321404 91026 321406
rect 95233 321403 95299 321406
rect 80697 320786 80763 320789
rect 89846 320786 89852 320788
rect 80697 320784 89852 320786
rect 80697 320728 80702 320784
rect 80758 320728 89852 320784
rect 80697 320726 89852 320728
rect 80697 320723 80763 320726
rect 89846 320724 89852 320726
rect 89916 320724 89922 320788
rect 142797 320242 142863 320245
rect 210366 320242 210372 320244
rect 142797 320240 210372 320242
rect 142797 320184 142802 320240
rect 142858 320184 210372 320240
rect 142797 320182 210372 320184
rect 142797 320179 142863 320182
rect 210366 320180 210372 320182
rect 210436 320180 210442 320244
rect 88241 319562 88307 319565
rect 98310 319562 98316 319564
rect 88241 319560 98316 319562
rect 88241 319504 88246 319560
rect 88302 319504 98316 319560
rect 88241 319502 98316 319504
rect 88241 319499 88307 319502
rect 98310 319500 98316 319502
rect 98380 319500 98386 319564
rect 81341 319426 81407 319429
rect 115974 319426 115980 319428
rect 81341 319424 115980 319426
rect -960 319290 480 319380
rect 81341 319368 81346 319424
rect 81402 319368 115980 319424
rect 81341 319366 115980 319368
rect 81341 319363 81407 319366
rect 115974 319364 115980 319366
rect 116044 319426 116050 319428
rect 262254 319426 262260 319428
rect 116044 319366 262260 319426
rect 116044 319364 116050 319366
rect 262254 319364 262260 319366
rect 262324 319364 262330 319428
rect 3417 319290 3483 319293
rect -960 319288 3483 319290
rect -960 319232 3422 319288
rect 3478 319232 3483 319288
rect -960 319230 3483 319232
rect -960 319140 480 319230
rect 3417 319227 3483 319230
rect 94814 318820 94820 318884
rect 94884 318882 94890 318884
rect 232497 318882 232563 318885
rect 94884 318880 232563 318882
rect 94884 318824 232502 318880
rect 232558 318824 232563 318880
rect 94884 318822 232563 318824
rect 94884 318820 94890 318822
rect 232497 318819 232563 318822
rect 77017 318746 77083 318749
rect 77334 318746 77340 318748
rect 77017 318744 77340 318746
rect 77017 318688 77022 318744
rect 77078 318688 77340 318744
rect 77017 318686 77340 318688
rect 77017 318683 77083 318686
rect 77334 318684 77340 318686
rect 77404 318684 77410 318748
rect 78581 318338 78647 318341
rect 87086 318338 87092 318340
rect 78581 318336 87092 318338
rect 78581 318280 78586 318336
rect 78642 318280 87092 318336
rect 78581 318278 87092 318280
rect 78581 318275 78647 318278
rect 87086 318276 87092 318278
rect 87156 318276 87162 318340
rect 103421 318338 103487 318341
rect 114686 318338 114692 318340
rect 103421 318336 114692 318338
rect 103421 318280 103426 318336
rect 103482 318280 114692 318336
rect 103421 318278 114692 318280
rect 103421 318275 103487 318278
rect 114686 318276 114692 318278
rect 114756 318276 114762 318340
rect 116577 318338 116643 318341
rect 122097 318338 122163 318341
rect 258390 318338 258396 318340
rect 116577 318336 258396 318338
rect 116577 318280 116582 318336
rect 116638 318280 122102 318336
rect 122158 318280 258396 318336
rect 116577 318278 258396 318280
rect 116577 318275 116643 318278
rect 122097 318275 122163 318278
rect 258390 318276 258396 318278
rect 258460 318276 258466 318340
rect 81525 318202 81591 318205
rect 116025 318202 116091 318205
rect 253054 318202 253060 318204
rect 81525 318200 253060 318202
rect 81525 318144 81530 318200
rect 81586 318144 116030 318200
rect 116086 318144 253060 318200
rect 81525 318142 253060 318144
rect 81525 318139 81591 318142
rect 116025 318139 116091 318142
rect 253054 318140 253060 318142
rect 253124 318140 253130 318204
rect 79869 318066 79935 318069
rect 260046 318066 260052 318068
rect 79869 318064 260052 318066
rect 79869 318008 79874 318064
rect 79930 318008 260052 318064
rect 79869 318006 260052 318008
rect 79869 318003 79935 318006
rect 260046 318004 260052 318006
rect 260116 318004 260122 318068
rect 70209 317522 70275 317525
rect 75862 317522 75868 317524
rect 70209 317520 75868 317522
rect 70209 317464 70214 317520
rect 70270 317464 75868 317520
rect 70209 317462 75868 317464
rect 70209 317459 70275 317462
rect 75862 317460 75868 317462
rect 75932 317460 75938 317524
rect 69749 317386 69815 317389
rect 70301 317386 70367 317389
rect 69749 317384 70367 317386
rect 69749 317328 69754 317384
rect 69810 317328 70306 317384
rect 70362 317328 70367 317384
rect 69749 317326 70367 317328
rect 69749 317323 69815 317326
rect 70301 317323 70367 317326
rect 87045 316706 87111 316709
rect 98126 316706 98132 316708
rect 87045 316704 98132 316706
rect 87045 316648 87050 316704
rect 87106 316648 98132 316704
rect 87045 316646 98132 316648
rect 87045 316643 87111 316646
rect 98126 316644 98132 316646
rect 98196 316644 98202 316708
rect 125409 316706 125475 316709
rect 249149 316706 249215 316709
rect 125409 316704 249215 316706
rect 125409 316648 125414 316704
rect 125470 316648 249154 316704
rect 249210 316648 249215 316704
rect 125409 316646 249215 316648
rect 125409 316643 125475 316646
rect 249149 316643 249215 316646
rect 69749 316162 69815 316165
rect 266629 316162 266695 316165
rect 69749 316160 266695 316162
rect 69749 316104 69754 316160
rect 69810 316104 266634 316160
rect 266690 316104 266695 316160
rect 69749 316102 266695 316104
rect 69749 316099 69815 316102
rect 266629 316099 266695 316102
rect 77109 314938 77175 314941
rect 258390 314938 258396 314940
rect 77109 314936 258396 314938
rect 77109 314880 77114 314936
rect 77170 314880 258396 314936
rect 77109 314878 258396 314880
rect 77109 314875 77175 314878
rect 258390 314876 258396 314878
rect 258460 314876 258466 314940
rect 39297 314802 39363 314805
rect 224033 314802 224099 314805
rect 39297 314800 224099 314802
rect 39297 314744 39302 314800
rect 39358 314744 224038 314800
rect 224094 314744 224099 314800
rect 39297 314742 224099 314744
rect 39297 314739 39363 314742
rect 224033 314739 224099 314742
rect 35157 313442 35223 313445
rect 220905 313442 220971 313445
rect 35157 313440 220971 313442
rect 35157 313384 35162 313440
rect 35218 313384 220910 313440
rect 220966 313384 220971 313440
rect 35157 313382 220971 313384
rect 35157 313379 35223 313382
rect 220905 313379 220971 313382
rect 72417 313306 72483 313309
rect 263685 313306 263751 313309
rect 72417 313304 263751 313306
rect 72417 313248 72422 313304
rect 72478 313248 263690 313304
rect 263746 313248 263751 313304
rect 72417 313246 263751 313248
rect 72417 313243 72483 313246
rect 263685 313243 263751 313246
rect 89437 312490 89503 312493
rect 89437 312488 103530 312490
rect 89437 312432 89442 312488
rect 89498 312432 103530 312488
rect 89437 312430 103530 312432
rect 89437 312427 89503 312430
rect 66478 312156 66484 312220
rect 66548 312218 66554 312220
rect 67265 312218 67331 312221
rect 66548 312216 67331 312218
rect 66548 312160 67270 312216
rect 67326 312160 67331 312216
rect 66548 312158 67331 312160
rect 66548 312156 66554 312158
rect 67265 312155 67331 312158
rect 66662 312020 66668 312084
rect 66732 312082 66738 312084
rect 66897 312082 66963 312085
rect 66732 312080 66963 312082
rect 66732 312024 66902 312080
rect 66958 312024 66963 312080
rect 66732 312022 66963 312024
rect 103470 312082 103530 312430
rect 119981 312218 120047 312221
rect 240133 312218 240199 312221
rect 119981 312216 240199 312218
rect 119981 312160 119986 312216
rect 120042 312160 240138 312216
rect 240194 312160 240199 312216
rect 119981 312158 240199 312160
rect 119981 312155 120047 312158
rect 240133 312155 240199 312158
rect 121453 312082 121519 312085
rect 254025 312082 254091 312085
rect 103470 312080 254091 312082
rect 103470 312024 121458 312080
rect 121514 312024 254030 312080
rect 254086 312024 254091 312080
rect 103470 312022 254091 312024
rect 66732 312020 66738 312022
rect 66897 312019 66963 312022
rect 121453 312019 121519 312022
rect 254025 312019 254091 312022
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 30281 311946 30347 311949
rect 203609 311946 203675 311949
rect 30281 311944 203675 311946
rect 30281 311888 30286 311944
rect 30342 311888 203614 311944
rect 203670 311888 203675 311944
rect 583520 311932 584960 312022
rect 30281 311886 203675 311888
rect 30281 311883 30347 311886
rect 203609 311883 203675 311886
rect 191097 310858 191163 310861
rect 201534 310858 201540 310860
rect 191097 310856 201540 310858
rect 191097 310800 191102 310856
rect 191158 310800 201540 310856
rect 191097 310798 201540 310800
rect 191097 310795 191163 310798
rect 201534 310796 201540 310798
rect 201604 310796 201610 310860
rect 37181 310722 37247 310725
rect 204897 310722 204963 310725
rect 37181 310720 204963 310722
rect 37181 310664 37186 310720
rect 37242 310664 204902 310720
rect 204958 310664 204963 310720
rect 37181 310662 204963 310664
rect 37181 310659 37247 310662
rect 204897 310659 204963 310662
rect 34421 310586 34487 310589
rect 204253 310586 204319 310589
rect 34421 310584 204319 310586
rect 34421 310528 34426 310584
rect 34482 310528 204258 310584
rect 204314 310528 204319 310584
rect 34421 310526 204319 310528
rect 34421 310523 34487 310526
rect 204253 310523 204319 310526
rect 285673 310450 285739 310453
rect 286317 310450 286383 310453
rect 285673 310448 286383 310450
rect 285673 310392 285678 310448
rect 285734 310392 286322 310448
rect 286378 310392 286383 310448
rect 285673 310390 286383 310392
rect 285673 310387 285739 310390
rect 286317 310387 286383 310390
rect 187049 309498 187115 309501
rect 208393 309498 208459 309501
rect 187049 309496 208459 309498
rect 187049 309440 187054 309496
rect 187110 309440 208398 309496
rect 208454 309440 208459 309496
rect 187049 309438 208459 309440
rect 187049 309435 187115 309438
rect 208393 309435 208459 309438
rect 189717 309362 189783 309365
rect 285673 309362 285739 309365
rect 189717 309360 285739 309362
rect 189717 309304 189722 309360
rect 189778 309304 285678 309360
rect 285734 309304 285739 309360
rect 189717 309302 285739 309304
rect 189717 309299 189783 309302
rect 285673 309299 285739 309302
rect 17861 309226 17927 309229
rect 201769 309226 201835 309229
rect 17861 309224 201835 309226
rect 17861 309168 17866 309224
rect 17922 309168 201774 309224
rect 201830 309168 201835 309224
rect 17861 309166 201835 309168
rect 17861 309163 17927 309166
rect 201769 309163 201835 309166
rect 92289 308410 92355 308413
rect 92289 308408 122850 308410
rect 92289 308352 92294 308408
rect 92350 308352 122850 308408
rect 92289 308350 122850 308352
rect 92289 308347 92355 308350
rect 122790 307866 122850 308350
rect 201534 308212 201540 308276
rect 201604 308274 201610 308276
rect 202505 308274 202571 308277
rect 201604 308272 202571 308274
rect 201604 308216 202510 308272
rect 202566 308216 202571 308272
rect 201604 308214 202571 308216
rect 201604 308212 201610 308214
rect 202505 308211 202571 308214
rect 155217 308138 155283 308141
rect 219985 308138 220051 308141
rect 155217 308136 220051 308138
rect 155217 308080 155222 308136
rect 155278 308080 219990 308136
rect 220046 308080 220051 308136
rect 155217 308078 220051 308080
rect 155217 308075 155283 308078
rect 219985 308075 220051 308078
rect 137277 308002 137343 308005
rect 218053 308002 218119 308005
rect 137277 308000 218119 308002
rect 137277 307944 137282 308000
rect 137338 307944 218058 308000
rect 218114 307944 218119 308000
rect 137277 307942 218119 307944
rect 137277 307939 137343 307942
rect 218053 307939 218119 307942
rect 124213 307866 124279 307869
rect 258073 307866 258139 307869
rect 122790 307864 258139 307866
rect 122790 307808 124218 307864
rect 124274 307808 258078 307864
rect 258134 307808 258139 307864
rect 122790 307806 258139 307808
rect 124213 307803 124279 307806
rect 258073 307803 258139 307806
rect 244917 307050 244983 307053
rect 254526 307050 254532 307052
rect 244917 307048 254532 307050
rect 244917 306992 244922 307048
rect 244978 306992 254532 307048
rect 244917 306990 254532 306992
rect 244917 306987 244983 306990
rect 254526 306988 254532 306990
rect 254596 306988 254602 307052
rect 1301 306778 1367 306781
rect 196985 306778 197051 306781
rect 1301 306776 197051 306778
rect 1301 306720 1306 306776
rect 1362 306720 196990 306776
rect 197046 306720 197051 306776
rect 1301 306718 197051 306720
rect 1301 306715 1367 306718
rect 196985 306715 197051 306718
rect 188337 306642 188403 306645
rect 209773 306642 209839 306645
rect 188337 306640 209839 306642
rect 188337 306584 188342 306640
rect 188398 306584 209778 306640
rect 209834 306584 209839 306640
rect 188337 306582 209839 306584
rect 188337 306579 188403 306582
rect 209773 306579 209839 306582
rect 197302 306444 197308 306508
rect 197372 306506 197378 306508
rect 262489 306506 262555 306509
rect 197372 306504 262555 306506
rect 197372 306448 262494 306504
rect 262550 306448 262555 306504
rect 197372 306446 262555 306448
rect 197372 306444 197378 306446
rect 262489 306443 262555 306446
rect -960 306234 480 306324
rect 3233 306234 3299 306237
rect -960 306232 3299 306234
rect -960 306176 3238 306232
rect 3294 306176 3299 306232
rect -960 306174 3299 306176
rect -960 306084 480 306174
rect 3233 306171 3299 306174
rect 180149 305282 180215 305285
rect 214833 305282 214899 305285
rect 180149 305280 214899 305282
rect 180149 305224 180154 305280
rect 180210 305224 214838 305280
rect 214894 305224 214899 305280
rect 180149 305222 214899 305224
rect 180149 305219 180215 305222
rect 214833 305219 214899 305222
rect 177297 305146 177363 305149
rect 215477 305146 215543 305149
rect 177297 305144 215543 305146
rect 177297 305088 177302 305144
rect 177358 305088 215482 305144
rect 215538 305088 215543 305144
rect 177297 305086 215543 305088
rect 177297 305083 177363 305086
rect 215477 305083 215543 305086
rect 151169 305010 151235 305013
rect 203425 305010 203491 305013
rect 151169 305008 203491 305010
rect 151169 304952 151174 305008
rect 151230 304952 203430 305008
rect 203486 304952 203491 305008
rect 151169 304950 203491 304952
rect 151169 304947 151235 304950
rect 203425 304947 203491 304950
rect 73521 304194 73587 304197
rect 80646 304194 80652 304196
rect 73521 304192 80652 304194
rect 73521 304136 73526 304192
rect 73582 304136 80652 304192
rect 73521 304134 80652 304136
rect 73521 304131 73587 304134
rect 80646 304132 80652 304134
rect 80716 304194 80722 304196
rect 140129 304194 140195 304197
rect 80716 304192 140195 304194
rect 80716 304136 140134 304192
rect 140190 304136 140195 304192
rect 80716 304134 140195 304136
rect 80716 304132 80722 304134
rect 140129 304131 140195 304134
rect 249149 304194 249215 304197
rect 265157 304194 265223 304197
rect 249149 304192 265223 304194
rect 249149 304136 249154 304192
rect 249210 304136 265162 304192
rect 265218 304136 265223 304192
rect 249149 304134 265223 304136
rect 249149 304131 249215 304134
rect 265157 304131 265223 304134
rect 246113 304058 246179 304061
rect 276013 304058 276079 304061
rect 246113 304056 276079 304058
rect 246113 304000 246118 304056
rect 246174 304000 276018 304056
rect 276074 304000 276079 304056
rect 246113 303998 276079 304000
rect 246113 303995 246179 303998
rect 276013 303995 276079 303998
rect 159357 303922 159423 303925
rect 215293 303922 215359 303925
rect 159357 303920 215359 303922
rect 159357 303864 159362 303920
rect 159418 303864 215298 303920
rect 215354 303864 215359 303920
rect 159357 303862 215359 303864
rect 159357 303859 159423 303862
rect 215293 303859 215359 303862
rect 239254 303860 239260 303924
rect 239324 303922 239330 303924
rect 249333 303922 249399 303925
rect 239324 303920 249399 303922
rect 239324 303864 249338 303920
rect 249394 303864 249399 303920
rect 239324 303862 249399 303864
rect 239324 303860 239330 303862
rect 249333 303859 249399 303862
rect 182817 303786 182883 303789
rect 234613 303786 234679 303789
rect 182817 303784 234679 303786
rect 182817 303728 182822 303784
rect 182878 303728 234618 303784
rect 234674 303728 234679 303784
rect 182817 303726 234679 303728
rect 182817 303723 182883 303726
rect 234613 303723 234679 303726
rect 81249 303650 81315 303653
rect 83406 303650 83412 303652
rect 81249 303648 83412 303650
rect 81249 303592 81254 303648
rect 81310 303592 83412 303648
rect 81249 303590 83412 303592
rect 81249 303587 81315 303590
rect 83406 303588 83412 303590
rect 83476 303588 83482 303652
rect 213678 303588 213684 303652
rect 213748 303650 213754 303652
rect 213913 303650 213979 303653
rect 213748 303648 213979 303650
rect 213748 303592 213918 303648
rect 213974 303592 213979 303648
rect 213748 303590 213979 303592
rect 213748 303588 213754 303590
rect 213913 303587 213979 303590
rect 219934 303588 219940 303652
rect 220004 303650 220010 303652
rect 226977 303650 227043 303653
rect 220004 303648 227043 303650
rect 220004 303592 226982 303648
rect 227038 303592 227043 303648
rect 220004 303590 227043 303592
rect 220004 303588 220010 303590
rect 226977 303587 227043 303590
rect 237966 303588 237972 303652
rect 238036 303650 238042 303652
rect 240041 303650 240107 303653
rect 238036 303648 240107 303650
rect 238036 303592 240046 303648
rect 240102 303592 240107 303648
rect 238036 303590 240107 303592
rect 238036 303588 238042 303590
rect 240041 303587 240107 303590
rect 240685 303652 240751 303653
rect 240685 303648 240732 303652
rect 240796 303650 240802 303652
rect 240685 303592 240690 303648
rect 240685 303588 240732 303592
rect 240796 303590 240842 303650
rect 240796 303588 240802 303590
rect 242014 303588 242020 303652
rect 242084 303650 242090 303652
rect 242985 303650 243051 303653
rect 242084 303648 243051 303650
rect 242084 303592 242990 303648
rect 243046 303592 243051 303648
rect 242084 303590 243051 303592
rect 242084 303588 242090 303590
rect 240685 303587 240751 303588
rect 242985 303587 243051 303590
rect 249977 303650 250043 303653
rect 256877 303650 256943 303653
rect 249977 303648 256943 303650
rect 249977 303592 249982 303648
rect 250038 303592 256882 303648
rect 256938 303592 256943 303648
rect 249977 303590 256943 303592
rect 249977 303587 250043 303590
rect 256877 303587 256943 303590
rect 31017 302834 31083 302837
rect 195973 302834 196039 302837
rect 31017 302832 196039 302834
rect 31017 302776 31022 302832
rect 31078 302776 195978 302832
rect 196034 302776 196039 302832
rect 31017 302774 196039 302776
rect 31017 302771 31083 302774
rect 195973 302771 196039 302774
rect 247677 302834 247743 302837
rect 258257 302834 258323 302837
rect 247677 302832 258323 302834
rect 247677 302776 247682 302832
rect 247738 302776 258262 302832
rect 258318 302776 258323 302832
rect 247677 302774 258323 302776
rect 247677 302771 247743 302774
rect 258257 302771 258323 302774
rect 117957 302562 118023 302565
rect 248505 302562 248571 302565
rect 117957 302560 248571 302562
rect 117957 302504 117962 302560
rect 118018 302504 248510 302560
rect 248566 302504 248571 302560
rect 117957 302502 248571 302504
rect 117957 302499 118023 302502
rect 248505 302499 248571 302502
rect 189901 302426 189967 302429
rect 200205 302426 200271 302429
rect 189901 302424 200271 302426
rect 189901 302368 189906 302424
rect 189962 302368 200210 302424
rect 200266 302368 200271 302424
rect 189901 302366 200271 302368
rect 189901 302363 189967 302366
rect 200205 302363 200271 302366
rect 193438 302228 193444 302292
rect 193508 302290 193514 302292
rect 198273 302290 198339 302293
rect 193508 302288 198339 302290
rect 193508 302232 198278 302288
rect 198334 302232 198339 302288
rect 193508 302230 198339 302232
rect 193508 302228 193514 302230
rect 198273 302227 198339 302230
rect 251909 302290 251975 302293
rect 255313 302290 255379 302293
rect 251909 302288 255379 302290
rect 251909 302232 251914 302288
rect 251970 302232 255318 302288
rect 255374 302232 255379 302288
rect 251909 302230 255379 302232
rect 251909 302227 251975 302230
rect 255313 302227 255379 302230
rect 193254 301820 193260 301884
rect 193324 301882 193330 301884
rect 207841 301882 207907 301885
rect 193324 301880 207907 301882
rect 193324 301824 207846 301880
rect 207902 301824 207907 301880
rect 193324 301822 207907 301824
rect 193324 301820 193330 301822
rect 207841 301819 207907 301822
rect 251817 301746 251883 301749
rect 254158 301746 254164 301748
rect 251817 301744 254164 301746
rect 251817 301688 251822 301744
rect 251878 301688 254164 301744
rect 251817 301686 254164 301688
rect 251817 301683 251883 301686
rect 254158 301684 254164 301686
rect 254228 301684 254234 301748
rect 198733 301474 198799 301477
rect 180750 301472 198799 301474
rect 180750 301416 198738 301472
rect 198794 301416 198799 301472
rect 180750 301414 198799 301416
rect 16481 301338 16547 301341
rect 180750 301338 180810 301414
rect 198733 301411 198799 301414
rect 16481 301336 180810 301338
rect 16481 301280 16486 301336
rect 16542 301280 180810 301336
rect 16481 301278 180810 301280
rect 188705 301338 188771 301341
rect 188705 301336 195990 301338
rect 188705 301280 188710 301336
rect 188766 301280 195990 301336
rect 188705 301278 195990 301280
rect 16481 301275 16547 301278
rect 188705 301275 188771 301278
rect 188521 301202 188587 301205
rect 194225 301202 194291 301205
rect 188521 301200 194291 301202
rect 188521 301144 188526 301200
rect 188582 301144 194230 301200
rect 194286 301144 194291 301200
rect 188521 301142 194291 301144
rect 195930 301202 195990 301278
rect 224166 301276 224172 301340
rect 224236 301338 224242 301340
rect 224769 301338 224835 301341
rect 224236 301336 224835 301338
rect 224236 301280 224774 301336
rect 224830 301280 224835 301336
rect 224236 301278 224835 301280
rect 224236 301276 224242 301278
rect 224769 301275 224835 301278
rect 233182 301276 233188 301340
rect 233252 301338 233258 301340
rect 233785 301338 233851 301341
rect 233252 301336 233851 301338
rect 233252 301280 233790 301336
rect 233846 301280 233851 301336
rect 233252 301278 233851 301280
rect 233252 301276 233258 301278
rect 233785 301275 233851 301278
rect 234654 301276 234660 301340
rect 234724 301338 234730 301340
rect 235625 301338 235691 301341
rect 234724 301336 235691 301338
rect 234724 301280 235630 301336
rect 235686 301280 235691 301336
rect 234724 301278 235691 301280
rect 234724 301276 234730 301278
rect 235625 301275 235691 301278
rect 236494 301276 236500 301340
rect 236564 301338 236570 301340
rect 236913 301338 236979 301341
rect 236564 301336 236979 301338
rect 236564 301280 236918 301336
rect 236974 301280 236979 301336
rect 236564 301278 236979 301280
rect 236564 301276 236570 301278
rect 236913 301275 236979 301278
rect 238150 301276 238156 301340
rect 238220 301338 238226 301340
rect 239489 301338 239555 301341
rect 238220 301336 239555 301338
rect 238220 301280 239494 301336
rect 239550 301280 239555 301336
rect 238220 301278 239555 301280
rect 238220 301276 238226 301278
rect 239489 301275 239555 301278
rect 200573 301202 200639 301205
rect 195930 301200 200639 301202
rect 195930 301144 200578 301200
rect 200634 301144 200639 301200
rect 195930 301142 200639 301144
rect 188521 301139 188587 301142
rect 194225 301139 194291 301142
rect 200573 301139 200639 301142
rect 212390 301140 212396 301204
rect 212460 301202 212466 301204
rect 212460 301142 252908 301202
rect 212460 301140 212466 301142
rect 215886 301004 215892 301068
rect 215956 301066 215962 301068
rect 218421 301066 218487 301069
rect 215956 301064 218487 301066
rect 215956 301008 218426 301064
rect 218482 301008 218487 301064
rect 215956 301006 218487 301008
rect 215956 301004 215962 301006
rect 218421 301003 218487 301006
rect 218646 301004 218652 301068
rect 218716 301066 218722 301068
rect 244549 301066 244615 301069
rect 218716 301064 244615 301066
rect 218716 301008 244554 301064
rect 244610 301008 244615 301064
rect 218716 301006 244615 301008
rect 218716 301004 218722 301006
rect 244549 301003 244615 301006
rect 253473 301066 253539 301069
rect 277393 301066 277459 301069
rect 253473 301064 277459 301066
rect 253473 301008 253478 301064
rect 253534 301008 277398 301064
rect 277454 301008 277459 301064
rect 253473 301006 277459 301008
rect 253473 301003 253539 301006
rect 277393 301003 277459 301006
rect 190453 300930 190519 300933
rect 190453 300928 193660 300930
rect 190453 300872 190458 300928
rect 190514 300872 193660 300928
rect 190453 300870 193660 300872
rect 190453 300867 190519 300870
rect 194542 300868 194548 300932
rect 194612 300930 194618 300932
rect 194685 300930 194751 300933
rect 197353 300930 197419 300933
rect 194612 300928 194751 300930
rect 194612 300872 194690 300928
rect 194746 300872 194751 300928
rect 194612 300870 194751 300872
rect 194612 300868 194618 300870
rect 194685 300867 194751 300870
rect 197310 300928 197419 300930
rect 197310 300872 197358 300928
rect 197414 300872 197419 300928
rect 197310 300867 197419 300872
rect 198774 300868 198780 300932
rect 198844 300930 198850 300932
rect 199285 300930 199351 300933
rect 198844 300928 199351 300930
rect 198844 300872 199290 300928
rect 199346 300872 199351 300928
rect 198844 300870 199351 300872
rect 198844 300868 198850 300870
rect 199285 300867 199351 300870
rect 204846 300868 204852 300932
rect 204916 300930 204922 300932
rect 205633 300930 205699 300933
rect 204916 300928 205699 300930
rect 204916 300872 205638 300928
rect 205694 300872 205699 300928
rect 204916 300870 205699 300872
rect 204916 300868 204922 300870
rect 205633 300867 205699 300870
rect 205766 300868 205772 300932
rect 205836 300930 205842 300932
rect 206277 300930 206343 300933
rect 207105 300932 207171 300933
rect 207054 300930 207060 300932
rect 205836 300928 206343 300930
rect 205836 300872 206282 300928
rect 206338 300872 206343 300928
rect 205836 300870 206343 300872
rect 207014 300870 207060 300930
rect 207124 300928 207171 300932
rect 211521 300930 211587 300933
rect 207166 300872 207171 300928
rect 205836 300868 205842 300870
rect 206277 300867 206343 300870
rect 207054 300868 207060 300870
rect 207124 300868 207171 300872
rect 207105 300867 207171 300868
rect 211478 300928 211587 300930
rect 211478 300872 211526 300928
rect 211582 300872 211587 300928
rect 211478 300867 211587 300872
rect 214414 300868 214420 300932
rect 214484 300930 214490 300932
rect 217041 300930 217107 300933
rect 214484 300928 217107 300930
rect 214484 300872 217046 300928
rect 217102 300872 217107 300928
rect 214484 300870 217107 300872
rect 214484 300868 214490 300870
rect 217041 300867 217107 300870
rect 217174 300868 217180 300932
rect 217244 300930 217250 300932
rect 218973 300930 219039 300933
rect 217244 300928 219039 300930
rect 217244 300872 218978 300928
rect 219034 300872 219039 300928
rect 217244 300870 219039 300872
rect 217244 300868 217250 300870
rect 218973 300867 219039 300870
rect 219198 300868 219204 300932
rect 219268 300930 219274 300932
rect 219433 300930 219499 300933
rect 219268 300928 219499 300930
rect 219268 300872 219438 300928
rect 219494 300872 219499 300928
rect 219268 300870 219499 300872
rect 219268 300868 219274 300870
rect 219433 300867 219499 300870
rect 220854 300868 220860 300932
rect 220924 300930 220930 300932
rect 221641 300930 221707 300933
rect 222377 300932 222443 300933
rect 222326 300930 222332 300932
rect 220924 300928 221707 300930
rect 220924 300872 221646 300928
rect 221702 300872 221707 300928
rect 220924 300870 221707 300872
rect 222286 300870 222332 300930
rect 222396 300928 222443 300932
rect 222438 300872 222443 300928
rect 220924 300868 220930 300870
rect 221641 300867 221707 300870
rect 222326 300868 222332 300870
rect 222396 300868 222443 300872
rect 222377 300867 222443 300868
rect 224125 300930 224191 300933
rect 225965 300932 226031 300933
rect 226517 300932 226583 300933
rect 224350 300930 224356 300932
rect 224125 300928 224356 300930
rect 224125 300872 224130 300928
rect 224186 300872 224356 300928
rect 224125 300870 224356 300872
rect 224125 300867 224191 300870
rect 224350 300868 224356 300870
rect 224420 300868 224426 300932
rect 225965 300928 226012 300932
rect 226076 300930 226082 300932
rect 225965 300872 225970 300928
rect 225965 300868 226012 300872
rect 226076 300870 226122 300930
rect 226517 300928 226564 300932
rect 226628 300930 226634 300932
rect 226517 300872 226522 300928
rect 226076 300868 226082 300870
rect 226517 300868 226564 300872
rect 226628 300870 226674 300930
rect 226628 300868 226634 300870
rect 226742 300868 226748 300932
rect 226812 300930 226818 300932
rect 227253 300930 227319 300933
rect 226812 300928 227319 300930
rect 226812 300872 227258 300928
rect 227314 300872 227319 300928
rect 226812 300870 227319 300872
rect 226812 300868 226818 300870
rect 225965 300867 226031 300868
rect 226517 300867 226583 300868
rect 227253 300867 227319 300870
rect 229686 300868 229692 300932
rect 229756 300930 229762 300932
rect 229829 300930 229895 300933
rect 229756 300928 229895 300930
rect 229756 300872 229834 300928
rect 229890 300872 229895 300928
rect 229756 300870 229895 300872
rect 229756 300868 229762 300870
rect 229829 300867 229895 300870
rect 230422 300868 230428 300932
rect 230492 300930 230498 300932
rect 230565 300930 230631 300933
rect 230492 300928 230631 300930
rect 230492 300872 230570 300928
rect 230626 300872 230631 300928
rect 230492 300870 230631 300872
rect 230492 300868 230498 300870
rect 230565 300867 230631 300870
rect 230790 300868 230796 300932
rect 230860 300930 230866 300932
rect 231209 300930 231275 300933
rect 230860 300928 231275 300930
rect 230860 300872 231214 300928
rect 231270 300872 231275 300928
rect 230860 300870 231275 300872
rect 230860 300868 230866 300870
rect 231209 300867 231275 300870
rect 232037 300932 232103 300933
rect 232037 300928 232084 300932
rect 232148 300930 232154 300932
rect 232037 300872 232042 300928
rect 232037 300868 232084 300872
rect 232148 300870 232194 300930
rect 232148 300868 232154 300870
rect 232262 300868 232268 300932
rect 232332 300930 232338 300932
rect 232497 300930 232563 300933
rect 232332 300928 232563 300930
rect 232332 300872 232502 300928
rect 232558 300872 232563 300928
rect 232332 300870 232563 300872
rect 232332 300868 232338 300870
rect 232037 300867 232103 300868
rect 232497 300867 232563 300870
rect 233325 300932 233391 300933
rect 233325 300928 233372 300932
rect 233436 300930 233442 300932
rect 233325 300872 233330 300928
rect 233325 300868 233372 300872
rect 233436 300870 233482 300930
rect 233436 300868 233442 300870
rect 234838 300868 234844 300932
rect 234908 300930 234914 300932
rect 234981 300930 235047 300933
rect 234908 300928 235047 300930
rect 234908 300872 234986 300928
rect 235042 300872 235047 300928
rect 234908 300870 235047 300872
rect 234908 300868 234914 300870
rect 233325 300867 233391 300868
rect 234981 300867 235047 300870
rect 236637 300932 236703 300933
rect 236637 300928 236684 300932
rect 236748 300930 236754 300932
rect 236637 300872 236642 300928
rect 236637 300868 236684 300872
rect 236748 300870 236794 300930
rect 236748 300868 236754 300870
rect 238702 300868 238708 300932
rect 238772 300930 238778 300932
rect 238845 300930 238911 300933
rect 238772 300928 238911 300930
rect 238772 300872 238850 300928
rect 238906 300872 238911 300928
rect 238772 300870 238911 300872
rect 238772 300868 238778 300870
rect 236637 300867 236703 300868
rect 238845 300867 238911 300870
rect 240910 300868 240916 300932
rect 240980 300930 240986 300932
rect 241421 300930 241487 300933
rect 240980 300928 241487 300930
rect 240980 300872 241426 300928
rect 241482 300872 241487 300928
rect 240980 300870 241487 300872
rect 240980 300868 240986 300870
rect 241421 300867 241487 300870
rect 241646 300868 241652 300932
rect 241716 300930 241722 300932
rect 241973 300930 242039 300933
rect 241716 300928 242039 300930
rect 241716 300872 241978 300928
rect 242034 300872 242039 300928
rect 241716 300870 242039 300872
rect 241716 300868 241722 300870
rect 241973 300867 242039 300870
rect 242934 300868 242940 300932
rect 243004 300930 243010 300932
rect 243261 300930 243327 300933
rect 243004 300928 243327 300930
rect 243004 300872 243266 300928
rect 243322 300872 243327 300928
rect 243004 300870 243327 300872
rect 243004 300868 243010 300870
rect 243261 300867 243327 300870
rect 244406 300868 244412 300932
rect 244476 300930 244482 300932
rect 245101 300930 245167 300933
rect 244476 300928 245167 300930
rect 244476 300872 245106 300928
rect 245162 300872 245167 300928
rect 244476 300870 245167 300872
rect 244476 300868 244482 300870
rect 245101 300867 245167 300870
rect 245694 300868 245700 300932
rect 245764 300930 245770 300932
rect 246389 300930 246455 300933
rect 247769 300932 247835 300933
rect 248505 300932 248571 300933
rect 247718 300930 247724 300932
rect 245764 300928 246455 300930
rect 245764 300872 246394 300928
rect 246450 300872 246455 300928
rect 245764 300870 246455 300872
rect 247678 300870 247724 300930
rect 247788 300928 247835 300932
rect 247830 300872 247835 300928
rect 245764 300868 245770 300870
rect 246389 300867 246455 300870
rect 247718 300868 247724 300870
rect 247788 300868 247835 300872
rect 248454 300868 248460 300932
rect 248524 300930 248571 300932
rect 248524 300928 248616 300930
rect 248566 300872 248616 300928
rect 248524 300870 248616 300872
rect 248524 300868 248571 300870
rect 251214 300868 251220 300932
rect 251284 300930 251290 300932
rect 251541 300930 251607 300933
rect 251284 300928 251607 300930
rect 251284 300872 251546 300928
rect 251602 300872 251607 300928
rect 251284 300870 251607 300872
rect 251284 300868 251290 300870
rect 247769 300867 247835 300868
rect 248505 300867 248571 300868
rect 251541 300867 251607 300870
rect 252461 300932 252527 300933
rect 252461 300928 252508 300932
rect 252572 300930 252578 300932
rect 252461 300872 252466 300928
rect 252461 300868 252508 300872
rect 252572 300870 252618 300930
rect 252572 300868 252578 300870
rect 252461 300867 252527 300868
rect 86166 300732 86172 300796
rect 86236 300794 86242 300796
rect 89713 300794 89779 300797
rect 86236 300792 89779 300794
rect 86236 300736 89718 300792
rect 89774 300736 89779 300792
rect 86236 300734 89779 300736
rect 86236 300732 86242 300734
rect 89713 300731 89779 300734
rect 196566 300732 196572 300796
rect 196636 300794 196642 300796
rect 197310 300794 197370 300867
rect 196636 300734 197370 300794
rect 196636 300732 196642 300734
rect 208526 300732 208532 300796
rect 208596 300794 208602 300796
rect 211478 300794 211538 300867
rect 208596 300734 211538 300794
rect 208596 300732 208602 300734
rect 252878 300661 252938 300764
rect 191097 300658 191163 300661
rect 197302 300658 197308 300660
rect 191097 300656 197308 300658
rect 191097 300600 191102 300656
rect 191158 300600 197308 300656
rect 191097 300598 197308 300600
rect 191097 300595 191163 300598
rect 197302 300596 197308 300598
rect 197372 300596 197378 300660
rect 210366 300596 210372 300660
rect 210436 300658 210442 300660
rect 210436 300598 238770 300658
rect 252878 300656 252987 300661
rect 252878 300600 252926 300656
rect 252982 300600 252987 300656
rect 252878 300598 252987 300600
rect 210436 300596 210442 300598
rect 238710 300250 238770 300598
rect 252921 300595 252987 300598
rect 255446 300386 255452 300388
rect 253460 300326 255452 300386
rect 255446 300324 255452 300326
rect 255516 300324 255522 300388
rect 256734 300250 256740 300252
rect 238710 300190 256740 300250
rect 256734 300188 256740 300190
rect 256804 300188 256810 300252
rect 255405 299978 255471 299981
rect 253460 299976 255471 299978
rect 253460 299920 255410 299976
rect 255466 299920 255471 299976
rect 253460 299918 255471 299920
rect 255405 299915 255471 299918
rect 190545 299842 190611 299845
rect 190545 299840 193660 299842
rect 190545 299784 190550 299840
rect 190606 299784 193660 299840
rect 190545 299782 193660 299784
rect 190545 299779 190611 299782
rect 71865 299570 71931 299573
rect 73061 299570 73127 299573
rect 133229 299570 133295 299573
rect 71865 299568 133295 299570
rect 71865 299512 71870 299568
rect 71926 299512 73066 299568
rect 73122 299512 133234 299568
rect 133290 299512 133295 299568
rect 71865 299510 133295 299512
rect 71865 299507 71931 299510
rect 73061 299507 73127 299510
rect 133229 299507 133295 299510
rect 255262 299508 255268 299572
rect 255332 299570 255338 299572
rect 280245 299570 280311 299573
rect 255332 299568 280311 299570
rect 255332 299512 280250 299568
rect 280306 299512 280311 299568
rect 255332 299510 280311 299512
rect 255332 299508 255338 299510
rect 280245 299507 280311 299510
rect 256550 299434 256556 299436
rect 253460 299374 256556 299434
rect 256550 299372 256556 299374
rect 256620 299372 256626 299436
rect 254526 299026 254532 299028
rect 253460 298966 254532 299026
rect 254526 298964 254532 298966
rect 254596 299026 254602 299028
rect 255129 299026 255195 299029
rect 254596 299024 255195 299026
rect 254596 298968 255134 299024
rect 255190 298968 255195 299024
rect 254596 298966 255195 298968
rect 254596 298964 254602 298966
rect 255129 298963 255195 298966
rect 12249 298890 12315 298893
rect 193438 298890 193444 298892
rect 12249 298888 193444 298890
rect 12249 298832 12254 298888
rect 12310 298832 193444 298888
rect 12249 298830 193444 298832
rect 12249 298827 12315 298830
rect 193438 298828 193444 298830
rect 193508 298828 193514 298892
rect 71037 298754 71103 298757
rect 72734 298754 72740 298756
rect 71037 298752 72740 298754
rect 71037 298696 71042 298752
rect 71098 298696 72740 298752
rect 71037 298694 72740 298696
rect 71037 298691 71103 298694
rect 72734 298692 72740 298694
rect 72804 298754 72810 298756
rect 160093 298754 160159 298757
rect 72804 298752 160159 298754
rect 72804 298696 160098 298752
rect 160154 298696 160159 298752
rect 72804 298694 160159 298696
rect 72804 298692 72810 298694
rect 160093 298691 160159 298694
rect 255446 298692 255452 298756
rect 255516 298754 255522 298756
rect 281533 298754 281599 298757
rect 255516 298752 281599 298754
rect 255516 298696 281538 298752
rect 281594 298696 281599 298752
rect 255516 298694 281599 298696
rect 255516 298692 255522 298694
rect 281533 298691 281599 298694
rect 580257 298754 580323 298757
rect 583520 298754 584960 298844
rect 580257 298752 584960 298754
rect 580257 298696 580262 298752
rect 580318 298696 584960 298752
rect 580257 298694 584960 298696
rect 580257 298691 580323 298694
rect 191281 298618 191347 298621
rect 255262 298618 255268 298620
rect 191281 298616 193660 298618
rect 191281 298560 191286 298616
rect 191342 298560 193660 298616
rect 191281 298558 193660 298560
rect 253460 298558 255268 298618
rect 191281 298555 191347 298558
rect 255262 298556 255268 298558
rect 255332 298556 255338 298620
rect 583520 298604 584960 298694
rect 254526 298210 254532 298212
rect 253460 298150 254532 298210
rect 254526 298148 254532 298150
rect 254596 298148 254602 298212
rect 266353 298074 266419 298077
rect 266905 298074 266971 298077
rect 253430 298072 266971 298074
rect 253430 298016 266358 298072
rect 266414 298016 266910 298072
rect 266966 298016 266971 298072
rect 253430 298014 266971 298016
rect 253430 297772 253490 298014
rect 266353 298011 266419 298014
rect 266905 298011 266971 298014
rect 191189 297530 191255 297533
rect 191189 297528 193660 297530
rect 191189 297472 191194 297528
rect 191250 297472 193660 297528
rect 191189 297470 193660 297472
rect 191189 297467 191255 297470
rect 4061 297394 4127 297397
rect 190361 297394 190427 297397
rect 4061 297392 190427 297394
rect 4061 297336 4066 297392
rect 4122 297336 190366 297392
rect 190422 297336 190427 297392
rect 4061 297334 190427 297336
rect 4061 297331 4127 297334
rect 190361 297331 190427 297334
rect 266905 297394 266971 297397
rect 309777 297394 309843 297397
rect 266905 297392 309843 297394
rect 266905 297336 266910 297392
rect 266966 297336 309782 297392
rect 309838 297336 309843 297392
rect 266905 297334 309843 297336
rect 266905 297331 266971 297334
rect 309777 297331 309843 297334
rect 255497 297258 255563 297261
rect 253460 297256 255563 297258
rect 253460 297200 255502 297256
rect 255558 297200 255563 297256
rect 253460 297198 255563 297200
rect 255497 297195 255563 297198
rect 255589 296850 255655 296853
rect 253460 296848 255655 296850
rect 253460 296792 255594 296848
rect 255650 296792 255655 296848
rect 253460 296790 255655 296792
rect 255589 296787 255655 296790
rect 186957 296714 187023 296717
rect 193254 296714 193260 296716
rect 186957 296712 193260 296714
rect 186957 296656 186962 296712
rect 187018 296656 193260 296712
rect 186957 296654 193260 296656
rect 186957 296651 187023 296654
rect 193254 296652 193260 296654
rect 193324 296652 193330 296716
rect 192477 296578 192543 296581
rect 193070 296578 193076 296580
rect 192477 296576 193076 296578
rect 192477 296520 192482 296576
rect 192538 296520 193076 296576
rect 192477 296518 193076 296520
rect 192477 296515 192543 296518
rect 193070 296516 193076 296518
rect 193140 296516 193146 296580
rect 253933 296442 253999 296445
rect 253460 296440 253999 296442
rect 253460 296384 253938 296440
rect 253994 296384 253999 296440
rect 253460 296382 253999 296384
rect 253933 296379 253999 296382
rect 190453 296306 190519 296309
rect 190453 296304 193660 296306
rect 190453 296248 190458 296304
rect 190514 296248 193660 296304
rect 190453 296246 193660 296248
rect 190453 296243 190519 296246
rect 255681 296034 255747 296037
rect 253460 296032 255747 296034
rect 253460 295976 255686 296032
rect 255742 295976 255747 296032
rect 253460 295974 255747 295976
rect 255681 295971 255747 295974
rect 255497 295490 255563 295493
rect 253460 295488 255563 295490
rect 253460 295432 255502 295488
rect 255558 295432 255563 295488
rect 253460 295430 255563 295432
rect 255497 295427 255563 295430
rect 191598 295156 191604 295220
rect 191668 295218 191674 295220
rect 191668 295158 193660 295218
rect 191668 295156 191674 295158
rect 255589 295082 255655 295085
rect 253460 295080 255655 295082
rect 253460 295024 255594 295080
rect 255650 295024 255655 295080
rect 253460 295022 255655 295024
rect 255589 295019 255655 295022
rect 84193 294674 84259 294677
rect 94446 294674 94452 294676
rect 84193 294672 94452 294674
rect 84193 294616 84198 294672
rect 84254 294616 94452 294672
rect 84193 294614 94452 294616
rect 84193 294611 84259 294614
rect 94446 294612 94452 294614
rect 94516 294612 94522 294676
rect 101254 294612 101260 294676
rect 101324 294674 101330 294676
rect 114093 294674 114159 294677
rect 255497 294674 255563 294677
rect 101324 294672 114159 294674
rect 101324 294616 114098 294672
rect 114154 294616 114159 294672
rect 101324 294614 114159 294616
rect 253460 294672 255563 294674
rect 253460 294616 255502 294672
rect 255558 294616 255563 294672
rect 253460 294614 255563 294616
rect 101324 294612 101330 294614
rect 114093 294611 114159 294614
rect 255497 294611 255563 294614
rect 26141 294538 26207 294541
rect 189901 294538 189967 294541
rect 26141 294536 189967 294538
rect 26141 294480 26146 294536
rect 26202 294480 189906 294536
rect 189962 294480 189967 294536
rect 26141 294478 189967 294480
rect 26141 294475 26207 294478
rect 189901 294475 189967 294478
rect 256550 294476 256556 294540
rect 256620 294538 256626 294540
rect 278773 294538 278839 294541
rect 256620 294536 278839 294538
rect 256620 294480 278778 294536
rect 278834 294480 278839 294536
rect 256620 294478 278839 294480
rect 256620 294476 256626 294478
rect 278773 294475 278839 294478
rect 254158 294266 254164 294268
rect 253460 294206 254164 294266
rect 254158 294204 254164 294206
rect 254228 294266 254234 294268
rect 255957 294266 256023 294269
rect 254228 294264 256023 294266
rect 254228 294208 255962 294264
rect 256018 294208 256023 294264
rect 254228 294206 256023 294208
rect 254228 294204 254234 294206
rect 255957 294203 256023 294206
rect 190545 293994 190611 293997
rect 190545 293992 193660 293994
rect 190545 293936 190550 293992
rect 190606 293936 193660 293992
rect 190545 293934 193660 293936
rect 190545 293931 190611 293934
rect 253933 293858 253999 293861
rect 253460 293856 253999 293858
rect 253460 293800 253938 293856
rect 253994 293800 253999 293856
rect 253460 293798 253999 293800
rect 253933 293795 253999 293798
rect 93025 293316 93091 293317
rect 92974 293314 92980 293316
rect -960 293178 480 293268
rect 92934 293254 92980 293314
rect 93044 293312 93091 293316
rect 255589 293314 255655 293317
rect 93086 293256 93091 293312
rect 92974 293252 92980 293254
rect 93044 293252 93091 293256
rect 253460 293312 255655 293314
rect 253460 293256 255594 293312
rect 255650 293256 255655 293312
rect 253460 293254 255655 293256
rect 93025 293251 93091 293252
rect 255589 293251 255655 293254
rect 3417 293178 3483 293181
rect -960 293176 3483 293178
rect -960 293120 3422 293176
rect 3478 293120 3483 293176
rect -960 293118 3483 293120
rect -960 293028 480 293118
rect 3417 293115 3483 293118
rect 83406 293116 83412 293180
rect 83476 293178 83482 293180
rect 86953 293178 87019 293181
rect 83476 293176 87019 293178
rect 83476 293120 86958 293176
rect 87014 293120 87019 293176
rect 83476 293118 87019 293120
rect 83476 293116 83482 293118
rect 86953 293115 87019 293118
rect 173249 293178 173315 293181
rect 191373 293178 191439 293181
rect 173249 293176 191439 293178
rect 173249 293120 173254 293176
rect 173310 293120 191378 293176
rect 191434 293120 191439 293176
rect 173249 293118 191439 293120
rect 173249 293115 173315 293118
rect 191373 293115 191439 293118
rect 193121 292906 193187 292909
rect 255497 292906 255563 292909
rect 193121 292904 193660 292906
rect 193121 292848 193126 292904
rect 193182 292848 193660 292904
rect 193121 292846 193660 292848
rect 253460 292904 255563 292906
rect 253460 292848 255502 292904
rect 255558 292848 255563 292904
rect 253460 292846 255563 292848
rect 193121 292843 193187 292846
rect 255497 292843 255563 292846
rect 253606 292708 253612 292772
rect 253676 292770 253682 292772
rect 256969 292770 257035 292773
rect 253676 292768 257035 292770
rect 253676 292712 256974 292768
rect 257030 292712 257035 292768
rect 253676 292710 257035 292712
rect 253676 292708 253682 292710
rect 256969 292707 257035 292710
rect 69013 292634 69079 292637
rect 70158 292634 70164 292636
rect 69013 292632 70164 292634
rect 69013 292576 69018 292632
rect 69074 292576 70164 292632
rect 69013 292574 70164 292576
rect 69013 292571 69079 292574
rect 70158 292572 70164 292574
rect 70228 292634 70234 292636
rect 107009 292634 107075 292637
rect 70228 292632 107075 292634
rect 70228 292576 107014 292632
rect 107070 292576 107075 292632
rect 70228 292574 107075 292576
rect 70228 292572 70234 292574
rect 107009 292571 107075 292574
rect 255497 292498 255563 292501
rect 253460 292496 255563 292498
rect 253460 292440 255502 292496
rect 255558 292440 255563 292496
rect 253460 292438 255563 292440
rect 255497 292435 255563 292438
rect 100702 291892 100708 291956
rect 100772 291954 100778 291956
rect 101857 291954 101923 291957
rect 100772 291952 101923 291954
rect 100772 291896 101862 291952
rect 101918 291896 101923 291952
rect 100772 291894 101923 291896
rect 100772 291892 100778 291894
rect 101857 291891 101923 291894
rect 253430 291818 253490 292060
rect 264973 291818 265039 291821
rect 253430 291816 265039 291818
rect 253430 291760 264978 291816
rect 265034 291760 265039 291816
rect 253430 291758 265039 291760
rect 264973 291755 265039 291758
rect 191097 291682 191163 291685
rect 191097 291680 193660 291682
rect 191097 291624 191102 291680
rect 191158 291624 193660 291680
rect 191097 291622 193660 291624
rect 191097 291619 191163 291622
rect 255589 291546 255655 291549
rect 253460 291544 255655 291546
rect 253460 291488 255594 291544
rect 255650 291488 255655 291544
rect 253460 291486 255655 291488
rect 255589 291483 255655 291486
rect 76465 291274 76531 291277
rect 77109 291274 77175 291277
rect 103697 291274 103763 291277
rect 76465 291272 103763 291274
rect 76465 291216 76470 291272
rect 76526 291216 77114 291272
rect 77170 291216 103702 291272
rect 103758 291216 103763 291272
rect 76465 291214 103763 291216
rect 76465 291211 76531 291214
rect 77109 291211 77175 291214
rect 103697 291211 103763 291214
rect 66437 291138 66503 291141
rect 66897 291138 66963 291141
rect 188429 291138 188495 291141
rect 254117 291138 254183 291141
rect 66437 291136 188495 291138
rect 66437 291080 66442 291136
rect 66498 291080 66902 291136
rect 66958 291080 188434 291136
rect 188490 291080 188495 291136
rect 66437 291078 188495 291080
rect 253460 291136 254183 291138
rect 253460 291080 254122 291136
rect 254178 291080 254183 291136
rect 253460 291078 254183 291080
rect 66437 291075 66503 291078
rect 66897 291075 66963 291078
rect 188429 291075 188495 291078
rect 254117 291075 254183 291078
rect 256734 290730 256740 290732
rect 253460 290670 256740 290730
rect 256734 290668 256740 290670
rect 256804 290668 256810 290732
rect 193213 290594 193279 290597
rect 193213 290592 193660 290594
rect 193213 290536 193218 290592
rect 193274 290536 193660 290592
rect 193213 290534 193660 290536
rect 193213 290531 193279 290534
rect 57605 290458 57671 290461
rect 66437 290458 66503 290461
rect 57605 290456 66503 290458
rect 57605 290400 57610 290456
rect 57666 290400 66442 290456
rect 66498 290400 66503 290456
rect 57605 290398 66503 290400
rect 57605 290395 57671 290398
rect 66437 290395 66503 290398
rect 255497 290322 255563 290325
rect 253460 290320 255563 290322
rect 253460 290264 255502 290320
rect 255558 290264 255563 290320
rect 253460 290262 255563 290264
rect 255497 290259 255563 290262
rect 253013 290186 253079 290189
rect 253013 290184 253122 290186
rect 253013 290128 253018 290184
rect 253074 290128 253122 290184
rect 253013 290123 253122 290128
rect 77201 289914 77267 289917
rect 137461 289914 137527 289917
rect 77201 289912 137527 289914
rect 77201 289856 77206 289912
rect 77262 289856 137466 289912
rect 137522 289856 137527 289912
rect 253062 289884 253122 290123
rect 77201 289854 137527 289856
rect 77201 289851 77267 289854
rect 137461 289851 137527 289854
rect 54937 289778 55003 289781
rect 55121 289778 55187 289781
rect 189717 289778 189783 289781
rect 252921 289778 252987 289781
rect 54937 289776 189783 289778
rect 54937 289720 54942 289776
rect 54998 289720 55126 289776
rect 55182 289720 189722 289776
rect 189778 289720 189783 289776
rect 54937 289718 189783 289720
rect 54937 289715 55003 289718
rect 55121 289715 55187 289718
rect 189717 289715 189783 289718
rect 252878 289776 252987 289778
rect 252878 289720 252926 289776
rect 252982 289720 252987 289776
rect 252878 289715 252987 289720
rect 191005 289370 191071 289373
rect 191005 289368 193660 289370
rect 191005 289312 191010 289368
rect 191066 289312 193660 289368
rect 252878 289340 252938 289715
rect 191005 289310 193660 289312
rect 191005 289307 191071 289310
rect 82721 289100 82787 289101
rect 82670 289036 82676 289100
rect 82740 289098 82787 289100
rect 255589 289098 255655 289101
rect 583109 289098 583175 289101
rect 82740 289096 82832 289098
rect 82782 289040 82832 289096
rect 82740 289038 82832 289040
rect 255589 289096 583175 289098
rect 255589 289040 255594 289096
rect 255650 289040 583114 289096
rect 583170 289040 583175 289096
rect 255589 289038 583175 289040
rect 82740 289036 82787 289038
rect 82721 289035 82787 289036
rect 255589 289035 255655 289038
rect 583109 289035 583175 289038
rect 255497 288962 255563 288965
rect 253460 288960 255563 288962
rect 253460 288904 255502 288960
rect 255558 288904 255563 288960
rect 253460 288902 255563 288904
rect 255497 288899 255563 288902
rect 86769 288554 86835 288557
rect 110505 288554 110571 288557
rect 86769 288552 110571 288554
rect 86769 288496 86774 288552
rect 86830 288496 110510 288552
rect 110566 288496 110571 288552
rect 86769 288494 110571 288496
rect 86769 288491 86835 288494
rect 110505 288491 110571 288494
rect 135897 288554 135963 288557
rect 149789 288554 149855 288557
rect 256785 288554 256851 288557
rect 135897 288552 149855 288554
rect 135897 288496 135902 288552
rect 135958 288496 149794 288552
rect 149850 288496 149855 288552
rect 135897 288494 149855 288496
rect 253460 288552 256851 288554
rect 253460 288496 256790 288552
rect 256846 288496 256851 288552
rect 253460 288494 256851 288496
rect 135897 288491 135963 288494
rect 149789 288491 149855 288494
rect 256785 288491 256851 288494
rect 80329 288418 80395 288421
rect 81341 288418 81407 288421
rect 80329 288416 81407 288418
rect 80329 288360 80334 288416
rect 80390 288360 81346 288416
rect 81402 288360 81407 288416
rect 80329 288358 81407 288360
rect 80329 288355 80395 288358
rect 81341 288355 81407 288358
rect 89529 288418 89595 288421
rect 90214 288418 90220 288420
rect 89529 288416 90220 288418
rect 89529 288360 89534 288416
rect 89590 288360 90220 288416
rect 89529 288358 90220 288360
rect 89529 288355 89595 288358
rect 90214 288356 90220 288358
rect 90284 288356 90290 288420
rect 191741 288282 191807 288285
rect 191741 288280 193660 288282
rect 191741 288224 191746 288280
rect 191802 288224 193660 288280
rect 191741 288222 193660 288224
rect 191741 288219 191807 288222
rect 255497 288146 255563 288149
rect 253460 288144 255563 288146
rect 253460 288088 255502 288144
rect 255558 288088 255563 288144
rect 253460 288086 255563 288088
rect 255497 288083 255563 288086
rect 172421 287738 172487 287741
rect 191281 287738 191347 287741
rect 172421 287736 191347 287738
rect 172421 287680 172426 287736
rect 172482 287680 191286 287736
rect 191342 287680 191347 287736
rect 172421 287678 191347 287680
rect 172421 287675 172487 287678
rect 191281 287675 191347 287678
rect 254209 287602 254275 287605
rect 253460 287600 254275 287602
rect 253460 287544 254214 287600
rect 254270 287544 254275 287600
rect 253460 287542 254275 287544
rect 254209 287539 254275 287542
rect 93761 287466 93827 287469
rect 97993 287466 98059 287469
rect 93761 287464 98059 287466
rect 93761 287408 93766 287464
rect 93822 287408 97998 287464
rect 98054 287408 98059 287464
rect 93761 287406 98059 287408
rect 93761 287403 93827 287406
rect 97993 287403 98059 287406
rect 89253 287330 89319 287333
rect 97942 287330 97948 287332
rect 89253 287328 97948 287330
rect 89253 287272 89258 287328
rect 89314 287272 97948 287328
rect 89253 287270 97948 287272
rect 89253 287267 89319 287270
rect 97942 287268 97948 287270
rect 98012 287268 98018 287332
rect 80329 287194 80395 287197
rect 113173 287194 113239 287197
rect 255497 287194 255563 287197
rect 80329 287192 113239 287194
rect 80329 287136 80334 287192
rect 80390 287136 113178 287192
rect 113234 287136 113239 287192
rect 80329 287134 113239 287136
rect 253460 287192 255563 287194
rect 253460 287136 255502 287192
rect 255558 287136 255563 287192
rect 253460 287134 255563 287136
rect 80329 287131 80395 287134
rect 113173 287131 113239 287134
rect 255497 287131 255563 287134
rect 193998 286516 194058 287028
rect 255405 286786 255471 286789
rect 253460 286784 255471 286786
rect 253460 286728 255410 286784
rect 255466 286728 255471 286784
rect 253460 286726 255471 286728
rect 255405 286723 255471 286726
rect 193990 286452 193996 286516
rect 194060 286452 194066 286516
rect 94129 286378 94195 286381
rect 131113 286378 131179 286381
rect 160737 286378 160803 286381
rect 255589 286378 255655 286381
rect 94129 286376 160803 286378
rect 94129 286320 94134 286376
rect 94190 286320 131118 286376
rect 131174 286320 160742 286376
rect 160798 286320 160803 286376
rect 94129 286318 160803 286320
rect 253460 286376 255655 286378
rect 253460 286320 255594 286376
rect 255650 286320 255655 286376
rect 253460 286318 255655 286320
rect 94129 286315 94195 286318
rect 131113 286315 131179 286318
rect 160737 286315 160803 286318
rect 255589 286315 255655 286318
rect 78121 286242 78187 286245
rect 79501 286242 79567 286245
rect 78121 286240 79567 286242
rect 78121 286184 78126 286240
rect 78182 286184 79506 286240
rect 79562 286184 79567 286240
rect 78121 286182 79567 286184
rect 78121 286179 78187 286182
rect 79501 286179 79567 286182
rect 71313 286106 71379 286109
rect 71630 286106 71636 286108
rect 71313 286104 71636 286106
rect 71313 286048 71318 286104
rect 71374 286048 71636 286104
rect 71313 286046 71636 286048
rect 71313 286043 71379 286046
rect 71630 286044 71636 286046
rect 71700 286044 71706 286108
rect 93025 286106 93091 286109
rect 93669 286106 93735 286109
rect 93025 286104 93735 286106
rect 93025 286048 93030 286104
rect 93086 286048 93674 286104
rect 93730 286048 93735 286104
rect 93025 286046 93735 286048
rect 93025 286043 93091 286046
rect 93669 286043 93735 286046
rect 52085 285970 52151 285973
rect 75269 285970 75335 285973
rect 52085 285968 75335 285970
rect 52085 285912 52090 285968
rect 52146 285912 75274 285968
rect 75330 285912 75335 285968
rect 52085 285910 75335 285912
rect 52085 285907 52151 285910
rect 75269 285907 75335 285910
rect 191649 285970 191715 285973
rect 191649 285968 193660 285970
rect 191649 285912 191654 285968
rect 191710 285912 193660 285968
rect 191649 285910 193660 285912
rect 191649 285907 191715 285910
rect 50838 285772 50844 285836
rect 50908 285834 50914 285836
rect 69105 285834 69171 285837
rect 69749 285834 69815 285837
rect 50908 285832 69815 285834
rect 50908 285776 69110 285832
rect 69166 285776 69754 285832
rect 69810 285776 69815 285832
rect 50908 285774 69815 285776
rect 50908 285772 50914 285774
rect 69105 285771 69171 285774
rect 69749 285771 69815 285774
rect 69197 285698 69263 285701
rect 69606 285698 69612 285700
rect 69197 285696 69612 285698
rect 69197 285640 69202 285696
rect 69258 285640 69612 285696
rect 69197 285638 69612 285640
rect 69197 285635 69263 285638
rect 69606 285636 69612 285638
rect 69676 285636 69682 285700
rect 82445 285698 82511 285701
rect 82670 285698 82676 285700
rect 82445 285696 82676 285698
rect 82445 285640 82450 285696
rect 82506 285640 82676 285696
rect 82445 285638 82676 285640
rect 82445 285635 82511 285638
rect 82670 285636 82676 285638
rect 82740 285636 82746 285700
rect 88742 285636 88748 285700
rect 88812 285698 88818 285700
rect 89621 285698 89687 285701
rect 88812 285696 89687 285698
rect 88812 285640 89626 285696
rect 89682 285640 89687 285696
rect 88812 285638 89687 285640
rect 253430 285698 253490 285940
rect 262397 285698 262463 285701
rect 253430 285696 262463 285698
rect 253430 285640 262402 285696
rect 262458 285640 262463 285696
rect 253430 285638 262463 285640
rect 88812 285636 88818 285638
rect 89621 285635 89687 285638
rect 262397 285635 262463 285638
rect 91369 285562 91435 285565
rect 92289 285562 92355 285565
rect 91369 285560 92355 285562
rect 91369 285504 91374 285560
rect 91430 285504 92294 285560
rect 92350 285504 92355 285560
rect 91369 285502 92355 285504
rect 91369 285499 91435 285502
rect 92289 285499 92355 285502
rect 255497 285426 255563 285429
rect 253460 285424 255563 285426
rect 253460 285368 255502 285424
rect 255558 285368 255563 285424
rect 253460 285366 255563 285368
rect 255497 285363 255563 285366
rect 583520 285276 584960 285516
rect 255313 285018 255379 285021
rect 253460 285016 255379 285018
rect 253460 284960 255318 285016
rect 255374 284960 255379 285016
rect 253460 284958 255379 284960
rect 255313 284955 255379 284958
rect 256049 285018 256115 285021
rect 259821 285018 259887 285021
rect 256049 285016 259887 285018
rect 256049 284960 256054 285016
rect 256110 284960 259826 285016
rect 259882 284960 259887 285016
rect 256049 284958 259887 284960
rect 256049 284955 256115 284958
rect 259821 284955 259887 284958
rect 97942 284820 97948 284884
rect 98012 284882 98018 284884
rect 145649 284882 145715 284885
rect 98012 284880 145715 284882
rect 98012 284824 145654 284880
rect 145710 284824 145715 284880
rect 98012 284822 145715 284824
rect 98012 284820 98018 284822
rect 145649 284819 145715 284822
rect 158069 284882 158135 284885
rect 191189 284882 191255 284885
rect 158069 284880 191255 284882
rect 158069 284824 158074 284880
rect 158130 284824 191194 284880
rect 191250 284824 191255 284880
rect 158069 284822 191255 284824
rect 158069 284819 158135 284822
rect 191189 284819 191255 284822
rect 191557 284746 191623 284749
rect 191557 284744 193660 284746
rect 191557 284688 191562 284744
rect 191618 284688 193660 284744
rect 191557 284686 193660 284688
rect 191557 284683 191623 284686
rect 255405 284610 255471 284613
rect 253460 284608 255471 284610
rect 253460 284552 255410 284608
rect 255466 284552 255471 284608
rect 253460 284550 255471 284552
rect 255405 284547 255471 284550
rect 91369 284474 91435 284477
rect 100109 284474 100175 284477
rect 91369 284472 100175 284474
rect 91369 284416 91374 284472
rect 91430 284416 100114 284472
rect 100170 284416 100175 284472
rect 91369 284414 100175 284416
rect 91369 284411 91435 284414
rect 100109 284411 100175 284414
rect 61745 284338 61811 284341
rect 64689 284338 64755 284341
rect 134609 284338 134675 284341
rect 61745 284336 134675 284338
rect 61745 284280 61750 284336
rect 61806 284280 64694 284336
rect 64750 284280 134614 284336
rect 134670 284280 134675 284336
rect 61745 284278 134675 284280
rect 61745 284275 61811 284278
rect 64689 284275 64755 284278
rect 134609 284275 134675 284278
rect 71957 284202 72023 284205
rect 72366 284202 72372 284204
rect 71957 284200 72372 284202
rect 71957 284144 71962 284200
rect 72018 284144 72372 284200
rect 71957 284142 72372 284144
rect 71957 284139 72023 284142
rect 72366 284140 72372 284142
rect 72436 284140 72442 284204
rect 91318 284140 91324 284204
rect 91388 284202 91394 284204
rect 91461 284202 91527 284205
rect 91388 284200 91527 284202
rect 91388 284144 91466 284200
rect 91522 284144 91527 284200
rect 91388 284142 91527 284144
rect 91388 284140 91394 284142
rect 91461 284139 91527 284142
rect 102777 284202 102843 284205
rect 105813 284202 105879 284205
rect 255589 284202 255655 284205
rect 102777 284200 105879 284202
rect 102777 284144 102782 284200
rect 102838 284144 105818 284200
rect 105874 284144 105879 284200
rect 102777 284142 105879 284144
rect 253460 284200 255655 284202
rect 253460 284144 255594 284200
rect 255650 284144 255655 284200
rect 253460 284142 255655 284144
rect 102777 284139 102843 284142
rect 105813 284139 105879 284142
rect 255589 284139 255655 284142
rect 95182 283732 95188 283796
rect 95252 283794 95258 283796
rect 96015 283794 96081 283797
rect 96470 283794 96476 283796
rect 95252 283792 96476 283794
rect 95252 283736 96020 283792
rect 96076 283736 96476 283792
rect 95252 283734 96476 283736
rect 95252 283732 95258 283734
rect 96015 283731 96081 283734
rect 96470 283732 96476 283734
rect 96540 283732 96546 283796
rect 256601 283794 256667 283797
rect 253460 283792 256667 283794
rect 253460 283736 256606 283792
rect 256662 283736 256667 283792
rect 253460 283734 256667 283736
rect 256601 283731 256667 283734
rect 68870 283596 68876 283660
rect 68940 283658 68946 283660
rect 69197 283658 69263 283661
rect 68940 283656 69263 283658
rect 68940 283600 69202 283656
rect 69258 283600 69263 283656
rect 68940 283598 69263 283600
rect 68940 283596 68946 283598
rect 69197 283595 69263 283598
rect 69974 283596 69980 283660
rect 70044 283658 70050 283660
rect 70761 283658 70827 283661
rect 70044 283656 70827 283658
rect 70044 283600 70766 283656
rect 70822 283600 70827 283656
rect 70044 283598 70827 283600
rect 70044 283596 70050 283598
rect 70761 283595 70827 283598
rect 84694 283596 84700 283660
rect 84764 283658 84770 283660
rect 85389 283658 85455 283661
rect 84764 283656 85455 283658
rect 84764 283600 85394 283656
rect 85450 283600 85455 283656
rect 84764 283598 85455 283600
rect 84764 283596 84770 283598
rect 85389 283595 85455 283598
rect 191005 283658 191071 283661
rect 191005 283656 193660 283658
rect 191005 283600 191010 283656
rect 191066 283600 193660 283656
rect 191005 283598 193660 283600
rect 191005 283595 191071 283598
rect 73153 283524 73219 283525
rect 73102 283522 73108 283524
rect 73062 283462 73108 283522
rect 73172 283520 73219 283524
rect 73214 283464 73219 283520
rect 73102 283460 73108 283462
rect 73172 283460 73219 283464
rect 73153 283459 73219 283460
rect 89805 283524 89871 283525
rect 92565 283524 92631 283525
rect 89805 283520 89852 283524
rect 89916 283522 89922 283524
rect 89805 283464 89810 283520
rect 89805 283460 89852 283464
rect 89916 283462 89962 283522
rect 92565 283520 92612 283524
rect 92676 283522 92682 283524
rect 92565 283464 92570 283520
rect 89916 283460 89922 283462
rect 92565 283460 92612 283464
rect 92676 283462 92722 283522
rect 92676 283460 92682 283462
rect 89805 283459 89871 283460
rect 92565 283459 92631 283460
rect 61653 283250 61719 283253
rect 74349 283250 74415 283253
rect 75729 283252 75795 283253
rect 61653 283248 74415 283250
rect 61653 283192 61658 283248
rect 61714 283192 74354 283248
rect 74410 283192 74415 283248
rect 61653 283190 74415 283192
rect 61653 283187 61719 283190
rect 74349 283187 74415 283190
rect 75678 283188 75684 283252
rect 75748 283250 75795 283252
rect 255405 283250 255471 283253
rect 75748 283248 75840 283250
rect 75790 283192 75840 283248
rect 75748 283190 75840 283192
rect 253460 283248 255471 283250
rect 253460 283192 255410 283248
rect 255466 283192 255471 283248
rect 253460 283190 255471 283192
rect 75748 283188 75795 283190
rect 75729 283187 75795 283188
rect 255405 283187 255471 283190
rect 66805 282978 66871 282981
rect 66805 282976 68908 282978
rect 66805 282920 66810 282976
rect 66866 282920 68908 282976
rect 66805 282918 68908 282920
rect 66805 282915 66871 282918
rect 70342 282916 70348 282980
rect 70412 282978 70418 282980
rect 70945 282978 71011 282981
rect 70412 282976 71011 282978
rect 70412 282920 70950 282976
rect 71006 282920 71011 282976
rect 70412 282918 71011 282920
rect 70412 282916 70418 282918
rect 70945 282915 71011 282918
rect 80881 282978 80947 282981
rect 81249 282978 81315 282981
rect 87873 282980 87939 282981
rect 83958 282978 83964 282980
rect 80881 282976 83964 282978
rect 80881 282920 80886 282976
rect 80942 282920 81254 282976
rect 81310 282920 83964 282976
rect 80881 282918 83964 282920
rect 80881 282915 80947 282918
rect 81249 282915 81315 282918
rect 83958 282916 83964 282918
rect 84028 282916 84034 282980
rect 87822 282916 87828 282980
rect 87892 282978 87939 282980
rect 88517 282978 88583 282981
rect 88742 282978 88748 282980
rect 87892 282976 87984 282978
rect 87934 282920 87984 282976
rect 87892 282918 87984 282920
rect 88517 282976 88748 282978
rect 88517 282920 88522 282976
rect 88578 282920 88748 282976
rect 88517 282918 88748 282920
rect 87892 282916 87939 282918
rect 87873 282915 87939 282916
rect 88517 282915 88583 282918
rect 88742 282916 88748 282918
rect 88812 282916 88818 282980
rect 97901 282978 97967 282981
rect 98862 282978 98868 282980
rect 97901 282976 98868 282978
rect 97901 282920 97906 282976
rect 97962 282920 98868 282976
rect 97901 282918 98868 282920
rect 97901 282915 97967 282918
rect 98862 282916 98868 282918
rect 98932 282916 98938 282980
rect 127709 282978 127775 282981
rect 178033 282978 178099 282981
rect 127709 282976 178099 282978
rect 127709 282920 127714 282976
rect 127770 282920 178038 282976
rect 178094 282920 178099 282976
rect 127709 282918 178099 282920
rect 127709 282915 127775 282918
rect 178033 282915 178099 282918
rect 258165 282842 258231 282845
rect 253460 282840 258231 282842
rect 253460 282784 258170 282840
rect 258226 282784 258231 282840
rect 253460 282782 258231 282784
rect 258165 282779 258231 282782
rect 69013 282706 69079 282709
rect 100753 282708 100819 282709
rect 100702 282706 100708 282708
rect 69013 282704 69122 282706
rect 69013 282648 69018 282704
rect 69074 282648 69122 282704
rect 69013 282643 69122 282648
rect 98716 282646 100708 282706
rect 100772 282704 100819 282708
rect 100814 282648 100819 282704
rect 100702 282644 100708 282646
rect 100772 282644 100819 282648
rect 100753 282643 100819 282644
rect 69062 282132 69122 282643
rect 192385 282434 192451 282437
rect 193029 282434 193095 282437
rect 255405 282434 255471 282437
rect 192385 282432 193660 282434
rect 192385 282376 192390 282432
rect 192446 282376 193034 282432
rect 193090 282376 193660 282432
rect 192385 282374 193660 282376
rect 253460 282432 255471 282434
rect 253460 282376 255410 282432
rect 255466 282376 255471 282432
rect 253460 282374 255471 282376
rect 192385 282371 192451 282374
rect 193029 282371 193095 282374
rect 255405 282371 255471 282374
rect 255497 282026 255563 282029
rect 253460 282024 255563 282026
rect 253460 281968 255502 282024
rect 255558 281968 255563 282024
rect 253460 281966 255563 281968
rect 255497 281963 255563 281966
rect 98686 281618 98746 281860
rect 133965 281618 134031 281621
rect 138657 281618 138723 281621
rect 98686 281616 138723 281618
rect 98686 281560 133970 281616
rect 134026 281560 138662 281616
rect 138718 281560 138723 281616
rect 98686 281558 138723 281560
rect 133965 281555 134031 281558
rect 138657 281555 138723 281558
rect 255405 281482 255471 281485
rect 253460 281480 255471 281482
rect 253460 281424 255410 281480
rect 255466 281424 255471 281480
rect 253460 281422 255471 281424
rect 255405 281419 255471 281422
rect 191741 281346 191807 281349
rect 252829 281346 252895 281349
rect 191741 281344 193660 281346
rect 68878 281213 68938 281316
rect 191741 281288 191746 281344
rect 191802 281288 193660 281344
rect 191741 281286 193660 281288
rect 252829 281344 252938 281346
rect 252829 281288 252834 281344
rect 252890 281288 252938 281344
rect 191741 281283 191807 281286
rect 252829 281283 252938 281288
rect 68829 281208 68938 281213
rect 68829 281152 68834 281208
rect 68890 281152 68938 281208
rect 68829 281150 68938 281152
rect 68829 281147 68895 281150
rect 100753 281074 100819 281077
rect 98716 281072 100819 281074
rect 98716 281016 100758 281072
rect 100814 281016 100819 281072
rect 252878 281044 252938 281283
rect 98716 281014 100819 281016
rect 100753 281011 100819 281014
rect 134517 280802 134583 280805
rect 177297 280802 177363 280805
rect 134517 280800 177363 280802
rect 134517 280744 134522 280800
rect 134578 280744 177302 280800
rect 177358 280744 177363 280800
rect 134517 280742 177363 280744
rect 134517 280739 134583 280742
rect 177297 280739 177363 280742
rect 259637 280666 259703 280669
rect 253460 280664 259703 280666
rect 253460 280608 259642 280664
rect 259698 280608 259703 280664
rect 253460 280606 259703 280608
rect 259637 280603 259703 280606
rect 68001 280530 68067 280533
rect 68001 280528 68908 280530
rect 68001 280472 68006 280528
rect 68062 280472 68908 280528
rect 68001 280470 68908 280472
rect 68001 280467 68067 280470
rect 101489 280258 101555 280261
rect 255405 280258 255471 280261
rect 98716 280256 101555 280258
rect -960 279972 480 280212
rect 98716 280200 101494 280256
rect 101550 280200 101555 280256
rect 98716 280198 101555 280200
rect 253460 280256 255471 280258
rect 253460 280200 255410 280256
rect 255466 280200 255471 280256
rect 253460 280198 255471 280200
rect 101489 280195 101555 280198
rect 255405 280195 255471 280198
rect 190453 280122 190519 280125
rect 256601 280122 256667 280125
rect 190453 280120 193660 280122
rect 190453 280064 190458 280120
rect 190514 280064 193660 280120
rect 190453 280062 193660 280064
rect 253430 280120 256667 280122
rect 253430 280064 256606 280120
rect 256662 280064 256667 280120
rect 253430 280062 256667 280064
rect 190453 280059 190519 280062
rect 253430 279820 253490 280062
rect 256601 280059 256667 280062
rect 68553 279714 68619 279717
rect 68553 279712 68908 279714
rect 68553 279656 68558 279712
rect 68614 279656 68908 279712
rect 68553 279654 68908 279656
rect 68553 279651 68619 279654
rect 100753 279442 100819 279445
rect 98716 279440 100819 279442
rect 98716 279384 100758 279440
rect 100814 279384 100819 279440
rect 98716 279382 100819 279384
rect 100753 279379 100819 279382
rect 255313 279306 255379 279309
rect 253460 279304 255379 279306
rect 253460 279248 255318 279304
rect 255374 279248 255379 279304
rect 253460 279246 255379 279248
rect 255313 279243 255379 279246
rect 190361 279034 190427 279037
rect 190361 279032 193660 279034
rect 190361 278976 190366 279032
rect 190422 278976 193660 279032
rect 190361 278974 193660 278976
rect 190361 278971 190427 278974
rect 66529 278898 66595 278901
rect 261109 278898 261175 278901
rect 66529 278896 68908 278898
rect 66529 278840 66534 278896
rect 66590 278840 68908 278896
rect 66529 278838 68908 278840
rect 253460 278896 261175 278898
rect 253460 278840 261114 278896
rect 261170 278840 261175 278896
rect 253460 278838 261175 278840
rect 66529 278835 66595 278838
rect 261109 278835 261175 278838
rect 101254 278626 101260 278628
rect 98716 278566 101260 278626
rect 101254 278564 101260 278566
rect 101324 278564 101330 278628
rect 254025 278490 254091 278493
rect 253460 278488 254091 278490
rect 253460 278432 254030 278488
rect 254086 278432 254091 278488
rect 253460 278430 254091 278432
rect 254025 278427 254091 278430
rect 66805 278082 66871 278085
rect 255497 278082 255563 278085
rect 66805 278080 68908 278082
rect 66805 278024 66810 278080
rect 66866 278024 68908 278080
rect 66805 278022 68908 278024
rect 253460 278080 255563 278082
rect 253460 278024 255502 278080
rect 255558 278024 255563 278080
rect 253460 278022 255563 278024
rect 66805 278019 66871 278022
rect 255497 278019 255563 278022
rect 99373 277810 99439 277813
rect 98716 277808 99439 277810
rect 98716 277752 99378 277808
rect 99434 277752 99439 277808
rect 98716 277750 99439 277752
rect 99373 277747 99439 277750
rect 191649 277810 191715 277813
rect 191649 277808 193660 277810
rect 191649 277752 191654 277808
rect 191710 277752 193660 277808
rect 191649 277750 193660 277752
rect 191649 277747 191715 277750
rect 59077 277674 59143 277677
rect 66294 277674 66300 277676
rect 59077 277672 66300 277674
rect 59077 277616 59082 277672
rect 59138 277616 66300 277672
rect 59077 277614 66300 277616
rect 59077 277611 59143 277614
rect 66294 277612 66300 277614
rect 66364 277612 66370 277676
rect 255405 277538 255471 277541
rect 253460 277536 255471 277538
rect 253460 277480 255410 277536
rect 255466 277480 255471 277536
rect 253460 277478 255471 277480
rect 255405 277475 255471 277478
rect 98862 277340 98868 277404
rect 98932 277402 98938 277404
rect 140865 277402 140931 277405
rect 98932 277400 140931 277402
rect 98932 277344 140870 277400
rect 140926 277344 140931 277400
rect 98932 277342 140931 277344
rect 98932 277340 98938 277342
rect 140865 277339 140931 277342
rect 66805 277266 66871 277269
rect 66805 277264 68908 277266
rect 66805 277208 66810 277264
rect 66866 277208 68908 277264
rect 66805 277206 68908 277208
rect 66805 277203 66871 277206
rect 255405 277130 255471 277133
rect 253460 277128 255471 277130
rect 253460 277072 255410 277128
rect 255466 277072 255471 277128
rect 253460 277070 255471 277072
rect 255405 277067 255471 277070
rect 100753 276994 100819 276997
rect 266445 276994 266511 276997
rect 98716 276992 100819 276994
rect 98716 276936 100758 276992
rect 100814 276936 100819 276992
rect 98716 276934 100819 276936
rect 100753 276931 100819 276934
rect 253430 276992 267750 276994
rect 253430 276936 266450 276992
rect 266506 276936 267750 276992
rect 253430 276934 267750 276936
rect 140865 276722 140931 276725
rect 155401 276722 155467 276725
rect 140865 276720 155467 276722
rect 140865 276664 140870 276720
rect 140926 276664 155406 276720
rect 155462 276664 155467 276720
rect 253430 276692 253490 276934
rect 266445 276931 266511 276934
rect 267690 276722 267750 276934
rect 276105 276722 276171 276725
rect 267690 276720 276171 276722
rect 140865 276662 155467 276664
rect 140865 276659 140931 276662
rect 155401 276659 155467 276662
rect 66897 276450 66963 276453
rect 66897 276448 68908 276450
rect 66897 276392 66902 276448
rect 66958 276392 68908 276448
rect 66897 276390 68908 276392
rect 66897 276387 66963 276390
rect 102225 276178 102291 276181
rect 98716 276176 102291 276178
rect 98716 276120 102230 276176
rect 102286 276120 102291 276176
rect 98716 276118 102291 276120
rect 102225 276115 102291 276118
rect 126237 276042 126303 276045
rect 193630 276042 193690 276692
rect 267690 276664 276110 276720
rect 276166 276664 276171 276720
rect 267690 276662 276171 276664
rect 276105 276659 276171 276662
rect 255497 276314 255563 276317
rect 253460 276312 255563 276314
rect 253460 276256 255502 276312
rect 255558 276256 255563 276312
rect 253460 276254 255563 276256
rect 255497 276251 255563 276254
rect 126237 276040 193690 276042
rect 126237 275984 126242 276040
rect 126298 275984 193690 276040
rect 126237 275982 193690 275984
rect 126237 275979 126303 275982
rect 255405 275906 255471 275909
rect 253460 275904 255471 275906
rect 253460 275848 255410 275904
rect 255466 275848 255471 275904
rect 253460 275846 255471 275848
rect 255405 275843 255471 275846
rect 66621 275634 66687 275637
rect 66621 275632 68908 275634
rect 66621 275576 66626 275632
rect 66682 275576 68908 275632
rect 66621 275574 68908 275576
rect 66621 275571 66687 275574
rect 64689 274818 64755 274821
rect 66294 274818 66300 274820
rect 64689 274816 66300 274818
rect 64689 274760 64694 274816
rect 64750 274760 66300 274816
rect 64689 274758 66300 274760
rect 64689 274755 64755 274758
rect 66294 274756 66300 274758
rect 66364 274818 66370 274820
rect 98686 274818 98746 275332
rect 66364 274758 68908 274818
rect 98686 274758 108314 274818
rect 66364 274756 66370 274758
rect 100845 274546 100911 274549
rect 98716 274544 100911 274546
rect 98716 274488 100850 274544
rect 100906 274488 100911 274544
rect 98716 274486 100911 274488
rect 108254 274546 108314 274758
rect 184054 274620 184060 274684
rect 184124 274682 184130 274684
rect 193630 274682 193690 275468
rect 255405 275362 255471 275365
rect 253460 275360 255471 275362
rect 253460 275304 255410 275360
rect 255466 275304 255471 275360
rect 253460 275302 255471 275304
rect 255405 275299 255471 275302
rect 252878 274821 252938 274924
rect 252829 274816 252938 274821
rect 252829 274760 252834 274816
rect 252890 274760 252938 274816
rect 252829 274758 252938 274760
rect 252829 274755 252895 274758
rect 184124 274622 193690 274682
rect 184124 274620 184130 274622
rect 144913 274546 144979 274549
rect 146201 274546 146267 274549
rect 255313 274546 255379 274549
rect 108254 274544 146267 274546
rect 108254 274488 144918 274544
rect 144974 274488 146206 274544
rect 146262 274488 146267 274544
rect 108254 274486 146267 274488
rect 253460 274544 255379 274546
rect 253460 274488 255318 274544
rect 255374 274488 255379 274544
rect 253460 274486 255379 274488
rect 100845 274483 100911 274486
rect 144913 274483 144979 274486
rect 146201 274483 146267 274486
rect 255313 274483 255379 274486
rect 191649 274410 191715 274413
rect 191649 274408 193660 274410
rect 191649 274352 191654 274408
rect 191710 274352 193660 274408
rect 191649 274350 193660 274352
rect 191649 274347 191715 274350
rect 255497 274138 255563 274141
rect 253460 274136 255563 274138
rect 253460 274080 255502 274136
rect 255558 274080 255563 274136
rect 253460 274078 255563 274080
rect 255497 274075 255563 274078
rect 68878 273458 68938 273972
rect 146201 273866 146267 273869
rect 170581 273866 170647 273869
rect 146201 273864 170647 273866
rect 146201 273808 146206 273864
rect 146262 273808 170586 273864
rect 170642 273808 170647 273864
rect 146201 273806 170647 273808
rect 146201 273803 146267 273806
rect 170581 273803 170647 273806
rect 100753 273730 100819 273733
rect 98716 273728 100819 273730
rect 98716 273672 100758 273728
rect 100814 273672 100819 273728
rect 98716 273670 100819 273672
rect 100753 273667 100819 273670
rect 64830 273398 68938 273458
rect 253430 273458 253490 273564
rect 264053 273458 264119 273461
rect 253430 273456 264119 273458
rect 253430 273400 264058 273456
rect 264114 273400 264119 273456
rect 253430 273398 264119 273400
rect 60549 273322 60615 273325
rect 61745 273322 61811 273325
rect 64830 273322 64890 273398
rect 264053 273395 264119 273398
rect 60549 273320 64890 273322
rect 60549 273264 60554 273320
rect 60610 273264 61750 273320
rect 61806 273264 64890 273320
rect 60549 273262 64890 273264
rect 60549 273259 60615 273262
rect 61745 273259 61811 273262
rect 66805 273186 66871 273189
rect 191557 273186 191623 273189
rect 255405 273186 255471 273189
rect 66805 273184 68908 273186
rect 66805 273128 66810 273184
rect 66866 273128 68908 273184
rect 66805 273126 68908 273128
rect 191557 273184 193660 273186
rect 191557 273128 191562 273184
rect 191618 273128 193660 273184
rect 191557 273126 193660 273128
rect 253460 273184 255471 273186
rect 253460 273128 255410 273184
rect 255466 273128 255471 273184
rect 253460 273126 255471 273128
rect 66805 273123 66871 273126
rect 191557 273123 191623 273126
rect 255405 273123 255471 273126
rect 265157 273050 265223 273053
rect 253430 273048 267750 273050
rect 253430 272992 265162 273048
rect 265218 272992 267750 273048
rect 253430 272990 267750 272992
rect 100753 272914 100819 272917
rect 98716 272912 100819 272914
rect 98716 272856 100758 272912
rect 100814 272856 100819 272912
rect 98716 272854 100819 272856
rect 100753 272851 100819 272854
rect 253430 272748 253490 272990
rect 265157 272987 265223 272990
rect 267690 272506 267750 272990
rect 271873 272506 271939 272509
rect 267690 272504 271939 272506
rect 267690 272448 271878 272504
rect 271934 272448 271939 272504
rect 267690 272446 271939 272448
rect 271873 272443 271939 272446
rect 60365 271962 60431 271965
rect 66069 271962 66135 271965
rect 68878 271962 68938 272340
rect 253430 272234 253490 272340
rect 261201 272234 261267 272237
rect 253430 272232 261267 272234
rect 253430 272176 261206 272232
rect 261262 272176 261267 272232
rect 253430 272174 261267 272176
rect 261201 272171 261267 272174
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 101121 272098 101187 272101
rect 98716 272096 101187 272098
rect 98716 272040 101126 272096
rect 101182 272040 101187 272096
rect 98716 272038 101187 272040
rect 101121 272035 101187 272038
rect 191649 272098 191715 272101
rect 191649 272096 193660 272098
rect 191649 272040 191654 272096
rect 191710 272040 193660 272096
rect 583520 272084 584960 272174
rect 191649 272038 193660 272040
rect 191649 272035 191715 272038
rect 256601 271962 256667 271965
rect 60365 271960 68938 271962
rect 60365 271904 60370 271960
rect 60426 271904 66074 271960
rect 66130 271904 68938 271960
rect 60365 271902 68938 271904
rect 253460 271960 256667 271962
rect 253460 271904 256606 271960
rect 256662 271904 256667 271960
rect 253460 271902 256667 271904
rect 60365 271899 60431 271902
rect 66069 271899 66135 271902
rect 256601 271899 256667 271902
rect 68878 271010 68938 271524
rect 256601 271418 256667 271421
rect 253460 271416 256667 271418
rect 253460 271360 256606 271416
rect 256662 271360 256667 271416
rect 253460 271358 256667 271360
rect 256601 271355 256667 271358
rect 99281 271282 99347 271285
rect 98716 271280 99347 271282
rect 98716 271252 99286 271280
rect 64830 270950 68938 271010
rect 98686 271224 99286 271252
rect 99342 271224 99347 271280
rect 98686 271222 99347 271224
rect 60641 270602 60707 270605
rect 64830 270602 64890 270950
rect 66253 270738 66319 270741
rect 98177 270738 98243 270741
rect 98686 270738 98746 271222
rect 99281 271219 99347 271222
rect 106181 271146 106247 271149
rect 114502 271146 114508 271148
rect 106181 271144 114508 271146
rect 106181 271088 106186 271144
rect 106242 271088 114508 271144
rect 106181 271086 114508 271088
rect 106181 271083 106247 271086
rect 114502 271084 114508 271086
rect 114572 271084 114578 271148
rect 258073 271010 258139 271013
rect 253460 271008 258139 271010
rect 66253 270736 68908 270738
rect 66253 270680 66258 270736
rect 66314 270680 68908 270736
rect 66253 270678 68908 270680
rect 98177 270736 98746 270738
rect 98177 270680 98182 270736
rect 98238 270680 98746 270736
rect 98177 270678 98746 270680
rect 66253 270675 66319 270678
rect 98177 270675 98243 270678
rect 60641 270600 64890 270602
rect 60641 270544 60646 270600
rect 60702 270544 64890 270600
rect 60641 270542 64890 270544
rect 189717 270602 189783 270605
rect 193630 270602 193690 270980
rect 253460 270952 258078 271008
rect 258134 270952 258139 271008
rect 253460 270950 258139 270952
rect 258073 270947 258139 270950
rect 260833 270874 260899 270877
rect 189717 270600 193690 270602
rect 189717 270544 189722 270600
rect 189778 270544 193690 270600
rect 253430 270872 260899 270874
rect 253430 270816 260838 270872
rect 260894 270816 260899 270872
rect 253430 270814 260899 270816
rect 253430 270572 253490 270814
rect 260833 270811 260899 270814
rect 189717 270542 193690 270544
rect 60641 270539 60707 270542
rect 189717 270539 189783 270542
rect 99465 270466 99531 270469
rect 100293 270466 100359 270469
rect 98716 270464 100359 270466
rect 98716 270408 99470 270464
rect 99526 270408 100298 270464
rect 100354 270408 100359 270464
rect 98716 270406 100359 270408
rect 99465 270403 99531 270406
rect 100293 270403 100359 270406
rect 255497 270194 255563 270197
rect 253460 270192 255563 270194
rect 253460 270136 255502 270192
rect 255558 270136 255563 270192
rect 253460 270134 255563 270136
rect 255497 270131 255563 270134
rect 39849 269786 39915 269789
rect 64638 269786 64644 269788
rect 39849 269784 64644 269786
rect 39849 269728 39854 269784
rect 39910 269728 64644 269784
rect 39849 269726 64644 269728
rect 39849 269723 39915 269726
rect 64638 269724 64644 269726
rect 64708 269786 64714 269788
rect 68878 269786 68938 269892
rect 143533 269786 143599 269789
rect 162209 269786 162275 269789
rect 64708 269726 68938 269786
rect 142110 269784 162275 269786
rect 142110 269728 143538 269784
rect 143594 269728 162214 269784
rect 162270 269728 162275 269784
rect 142110 269726 162275 269728
rect 64708 269724 64714 269726
rect 98686 269378 98746 269620
rect 142110 269378 142170 269726
rect 143533 269723 143599 269726
rect 162209 269723 162275 269726
rect 191649 269786 191715 269789
rect 255405 269786 255471 269789
rect 191649 269784 193660 269786
rect 191649 269728 191654 269784
rect 191710 269728 193660 269784
rect 191649 269726 193660 269728
rect 253460 269784 255471 269786
rect 253460 269728 255410 269784
rect 255466 269728 255471 269784
rect 253460 269726 255471 269728
rect 191649 269723 191715 269726
rect 255405 269723 255471 269726
rect 98686 269318 142170 269378
rect 259729 269242 259795 269245
rect 253460 269240 259795 269242
rect 253460 269184 259734 269240
rect 259790 269184 259795 269240
rect 253460 269182 259795 269184
rect 259729 269179 259795 269182
rect 68878 268562 68938 269076
rect 100753 268834 100819 268837
rect 255313 268834 255379 268837
rect 98716 268832 100819 268834
rect 98716 268776 100758 268832
rect 100814 268776 100819 268832
rect 98716 268774 100819 268776
rect 253460 268832 255379 268834
rect 253460 268776 255318 268832
rect 255374 268776 255379 268832
rect 253460 268774 255379 268776
rect 100753 268771 100819 268774
rect 255313 268771 255379 268774
rect 191649 268698 191715 268701
rect 191649 268696 193660 268698
rect 191649 268640 191654 268696
rect 191710 268640 193660 268696
rect 191649 268638 193660 268640
rect 191649 268635 191715 268638
rect 64830 268502 68938 268562
rect 102777 268562 102843 268565
rect 108246 268562 108252 268564
rect 102777 268560 108252 268562
rect 102777 268504 102782 268560
rect 102838 268504 108252 268560
rect 102777 268502 108252 268504
rect 50889 268426 50955 268429
rect 63033 268426 63099 268429
rect 64830 268426 64890 268502
rect 102777 268499 102843 268502
rect 108246 268500 108252 268502
rect 108316 268500 108322 268564
rect 50889 268424 64890 268426
rect 50889 268368 50894 268424
rect 50950 268368 63038 268424
rect 63094 268368 64890 268424
rect 50889 268366 64890 268368
rect 98729 268426 98795 268429
rect 176009 268426 176075 268429
rect 255405 268426 255471 268429
rect 98729 268424 176075 268426
rect 98729 268368 98734 268424
rect 98790 268368 176014 268424
rect 176070 268368 176075 268424
rect 98729 268366 176075 268368
rect 253460 268424 255471 268426
rect 253460 268368 255410 268424
rect 255466 268368 255471 268424
rect 253460 268366 255471 268368
rect 50889 268363 50955 268366
rect 63033 268363 63099 268366
rect 98729 268363 98795 268366
rect 176009 268363 176075 268366
rect 255405 268363 255471 268366
rect 66805 268290 66871 268293
rect 66805 268288 68908 268290
rect 66805 268232 66810 268288
rect 66866 268232 68908 268288
rect 66805 268230 68908 268232
rect 66805 268227 66871 268230
rect 263961 268154 264027 268157
rect 253430 268152 264027 268154
rect 253430 268096 263966 268152
rect 264022 268096 264027 268152
rect 253430 268094 264027 268096
rect 101213 268018 101279 268021
rect 98716 268016 101279 268018
rect 98716 267960 101218 268016
rect 101274 267960 101279 268016
rect 253430 267988 253490 268094
rect 263961 268091 264027 268094
rect 98716 267958 101279 267960
rect 101213 267955 101279 267958
rect 191281 267474 191347 267477
rect 259494 267474 259500 267476
rect 191281 267472 193660 267474
rect -960 267202 480 267292
rect 3509 267202 3575 267205
rect -960 267200 3575 267202
rect -960 267144 3514 267200
rect 3570 267144 3575 267200
rect -960 267142 3575 267144
rect -960 267052 480 267142
rect 3509 267139 3575 267142
rect 68878 266930 68938 267444
rect 191281 267416 191286 267472
rect 191342 267416 193660 267472
rect 252908 267444 259500 267474
rect 191281 267414 193660 267416
rect 252878 267414 259500 267444
rect 191281 267411 191347 267414
rect 252878 267341 252938 267414
rect 259494 267412 259500 267414
rect 259564 267412 259570 267476
rect 252878 267336 252987 267341
rect 252878 267280 252926 267336
rect 252982 267280 252987 267336
rect 252878 267278 252987 267280
rect 252921 267275 252987 267278
rect 100753 267202 100819 267205
rect 98716 267200 100819 267202
rect 98716 267144 100758 267200
rect 100814 267144 100819 267200
rect 98716 267142 100819 267144
rect 100753 267139 100819 267142
rect 110638 267004 110644 267068
rect 110708 267066 110714 267068
rect 136633 267066 136699 267069
rect 153929 267066 153995 267069
rect 255497 267066 255563 267069
rect 110708 267064 153995 267066
rect 110708 267008 136638 267064
rect 136694 267008 153934 267064
rect 153990 267008 153995 267064
rect 110708 267006 153995 267008
rect 253460 267064 255563 267066
rect 253460 267008 255502 267064
rect 255558 267008 255563 267064
rect 253460 267006 255563 267008
rect 110708 267004 110714 267006
rect 136633 267003 136699 267006
rect 153929 267003 153995 267006
rect 255497 267003 255563 267006
rect 64830 266870 68938 266930
rect 49601 266522 49667 266525
rect 64830 266522 64890 266870
rect 66805 266658 66871 266661
rect 255405 266658 255471 266661
rect 66805 266656 68908 266658
rect 66805 266600 66810 266656
rect 66866 266600 68908 266656
rect 66805 266598 68908 266600
rect 253460 266656 255471 266658
rect 253460 266600 255410 266656
rect 255466 266600 255471 266656
rect 253460 266598 255471 266600
rect 66805 266595 66871 266598
rect 255405 266595 255471 266598
rect 49601 266520 64890 266522
rect 49601 266464 49606 266520
rect 49662 266464 64890 266520
rect 49601 266462 64890 266464
rect 49601 266459 49667 266462
rect 108246 266386 108252 266388
rect 98716 266326 108252 266386
rect 108246 266324 108252 266326
rect 108316 266324 108322 266388
rect 191005 266386 191071 266389
rect 191005 266384 193660 266386
rect 191005 266328 191010 266384
rect 191066 266328 193660 266384
rect 191005 266326 193660 266328
rect 191005 266323 191071 266326
rect 254025 266250 254091 266253
rect 253460 266248 254091 266250
rect 253460 266192 254030 266248
rect 254086 266192 254091 266248
rect 253460 266190 254091 266192
rect 254025 266187 254091 266190
rect 255313 265842 255379 265845
rect 253460 265840 255379 265842
rect 68878 265298 68938 265812
rect 253460 265784 255318 265840
rect 255374 265784 255379 265840
rect 253460 265782 255379 265784
rect 255313 265779 255379 265782
rect 100845 265570 100911 265573
rect 98716 265568 100911 265570
rect 98716 265512 100850 265568
rect 100906 265512 100911 265568
rect 98716 265510 100911 265512
rect 100845 265507 100911 265510
rect 263685 265434 263751 265437
rect 268326 265434 268332 265436
rect 263685 265432 268332 265434
rect 263685 265376 263690 265432
rect 263746 265376 268332 265432
rect 263685 265374 268332 265376
rect 263685 265371 263751 265374
rect 268326 265372 268332 265374
rect 268396 265372 268402 265436
rect 258390 265298 258396 265300
rect 64830 265238 68938 265298
rect 253460 265238 258396 265298
rect 50521 265026 50587 265029
rect 50889 265026 50955 265029
rect 64830 265026 64890 265238
rect 258390 265236 258396 265238
rect 258460 265236 258466 265300
rect 65701 265164 65767 265165
rect 65701 265162 65748 265164
rect 65656 265160 65748 265162
rect 65812 265162 65818 265164
rect 191557 265162 191623 265165
rect 65656 265104 65706 265160
rect 65656 265102 65748 265104
rect 65701 265100 65748 265102
rect 65812 265102 68938 265162
rect 65812 265100 65818 265102
rect 65701 265099 65767 265100
rect 50521 265024 64890 265026
rect 50521 264968 50526 265024
rect 50582 264968 50894 265024
rect 50950 264968 64890 265024
rect 68878 264996 68938 265102
rect 191557 265160 193660 265162
rect 191557 265104 191562 265160
rect 191618 265104 193660 265160
rect 191557 265102 193660 265104
rect 191557 265099 191623 265102
rect 110638 265026 110644 265028
rect 50521 264966 64890 264968
rect 100710 264966 110644 265026
rect 50521 264963 50587 264966
rect 50889 264963 50955 264966
rect 100710 264890 100770 264966
rect 110638 264964 110644 264966
rect 110708 264964 110714 265028
rect 255497 264890 255563 264893
rect 98686 264830 100770 264890
rect 253460 264888 255563 264890
rect 253460 264832 255502 264888
rect 255558 264832 255563 264888
rect 253460 264830 255563 264832
rect 98686 264724 98746 264830
rect 255497 264827 255563 264830
rect 255313 264482 255379 264485
rect 253460 264480 255379 264482
rect 253460 264424 255318 264480
rect 255374 264424 255379 264480
rect 253460 264422 255379 264424
rect 255313 264419 255379 264422
rect 62021 263666 62087 263669
rect 64781 263666 64847 263669
rect 68878 263666 68938 264180
rect 256049 264074 256115 264077
rect 253460 264072 256115 264074
rect 100753 263938 100819 263941
rect 98716 263936 100819 263938
rect 98716 263880 100758 263936
rect 100814 263880 100819 263936
rect 98716 263878 100819 263880
rect 100753 263875 100819 263878
rect 62021 263664 68938 263666
rect 62021 263608 62026 263664
rect 62082 263608 64786 263664
rect 64842 263608 68938 263664
rect 62021 263606 68938 263608
rect 62021 263603 62087 263606
rect 64781 263603 64847 263606
rect 160686 263604 160692 263668
rect 160756 263666 160762 263668
rect 193630 263666 193690 264044
rect 253460 264016 256054 264072
rect 256110 264016 256115 264072
rect 253460 264014 256115 264016
rect 256049 264011 256115 264014
rect 160756 263606 193690 263666
rect 160756 263604 160762 263606
rect 66897 263394 66963 263397
rect 253430 263394 253490 263500
rect 66897 263392 68908 263394
rect 66897 263336 66902 263392
rect 66958 263336 68908 263392
rect 66897 263334 68908 263336
rect 253430 263334 258090 263394
rect 66897 263331 66963 263334
rect 101673 263122 101739 263125
rect 255405 263122 255471 263125
rect 98716 263120 101739 263122
rect 98716 263064 101678 263120
rect 101734 263064 101739 263120
rect 98716 263062 101739 263064
rect 253460 263120 255471 263122
rect 253460 263064 255410 263120
rect 255466 263064 255471 263120
rect 253460 263062 255471 263064
rect 101673 263059 101739 263062
rect 255405 263059 255471 263062
rect 258030 262986 258090 263334
rect 276197 262986 276263 262989
rect 280797 262986 280863 262989
rect 258030 262984 280863 262986
rect 258030 262928 276202 262984
rect 276258 262928 280802 262984
rect 280858 262928 280863 262984
rect 258030 262926 280863 262928
rect 276197 262923 276263 262926
rect 280797 262923 280863 262926
rect 108430 262788 108436 262852
rect 108500 262850 108506 262852
rect 128445 262850 128511 262853
rect 108500 262848 128511 262850
rect 108500 262792 128450 262848
rect 128506 262792 128511 262848
rect 108500 262790 128511 262792
rect 108500 262788 108506 262790
rect 128445 262787 128511 262790
rect 155309 262850 155375 262853
rect 180241 262850 180307 262853
rect 155309 262848 180307 262850
rect 155309 262792 155314 262848
rect 155370 262792 180246 262848
rect 180302 262792 180307 262848
rect 155309 262790 180307 262792
rect 155309 262787 155375 262790
rect 180241 262787 180307 262790
rect 191649 262850 191715 262853
rect 191649 262848 193660 262850
rect 191649 262792 191654 262848
rect 191710 262792 193660 262848
rect 191649 262790 193660 262792
rect 191649 262787 191715 262790
rect 261109 262714 261175 262717
rect 253460 262712 261175 262714
rect 253460 262656 261114 262712
rect 261170 262656 261175 262712
rect 253460 262654 261175 262656
rect 261109 262651 261175 262654
rect 66529 262578 66595 262581
rect 66529 262576 68908 262578
rect 66529 262520 66534 262576
rect 66590 262520 68908 262576
rect 66529 262518 68908 262520
rect 66529 262515 66595 262518
rect 100753 262306 100819 262309
rect 255405 262306 255471 262309
rect 98716 262304 100819 262306
rect 98716 262248 100758 262304
rect 100814 262248 100819 262304
rect 98716 262246 100819 262248
rect 253460 262304 255471 262306
rect 253460 262248 255410 262304
rect 255466 262248 255471 262304
rect 253460 262246 255471 262248
rect 100753 262243 100819 262246
rect 255405 262243 255471 262246
rect 255497 261900 255563 261901
rect 255446 261898 255452 261900
rect 253460 261838 255452 261898
rect 255516 261896 255563 261900
rect 255558 261840 255563 261896
rect 255446 261836 255452 261838
rect 255516 261836 255563 261840
rect 255497 261835 255563 261836
rect 66110 261700 66116 261764
rect 66180 261762 66186 261764
rect 191649 261762 191715 261765
rect 66180 261702 68908 261762
rect 191649 261760 193660 261762
rect 191649 261704 191654 261760
rect 191710 261704 193660 261760
rect 191649 261702 193660 261704
rect 66180 261700 66186 261702
rect 191649 261699 191715 261702
rect 100937 261490 101003 261493
rect 101397 261490 101463 261493
rect 98716 261488 101463 261490
rect 98716 261432 100942 261488
rect 100998 261432 101402 261488
rect 101458 261432 101463 261488
rect 98716 261430 101463 261432
rect 100937 261427 101003 261430
rect 101397 261427 101463 261430
rect 131849 261490 131915 261493
rect 182909 261490 182975 261493
rect 131849 261488 182975 261490
rect 131849 261432 131854 261488
rect 131910 261432 182914 261488
rect 182970 261432 182975 261488
rect 131849 261430 182975 261432
rect 131849 261427 131915 261430
rect 182909 261427 182975 261430
rect 255313 261354 255379 261357
rect 253460 261352 255379 261354
rect 253460 261296 255318 261352
rect 255374 261296 255379 261352
rect 253460 261294 255379 261296
rect 255313 261291 255379 261294
rect 66253 260946 66319 260949
rect 255405 260946 255471 260949
rect 66253 260944 68908 260946
rect 66253 260888 66258 260944
rect 66314 260888 68908 260944
rect 66253 260886 68908 260888
rect 253460 260944 255471 260946
rect 253460 260888 255410 260944
rect 255466 260888 255471 260944
rect 253460 260886 255471 260888
rect 66253 260883 66319 260886
rect 108246 260748 108252 260812
rect 108316 260810 108322 260812
rect 147673 260810 147739 260813
rect 255270 260812 255330 260886
rect 255405 260883 255471 260886
rect 108316 260808 147739 260810
rect 108316 260752 147678 260808
rect 147734 260752 147739 260808
rect 108316 260750 147739 260752
rect 108316 260748 108322 260750
rect 147673 260747 147739 260750
rect 255262 260748 255268 260812
rect 255332 260748 255338 260812
rect 100753 260674 100819 260677
rect 98716 260672 100819 260674
rect 98716 260616 100758 260672
rect 100814 260616 100819 260672
rect 98716 260614 100819 260616
rect 100753 260611 100819 260614
rect 191281 260538 191347 260541
rect 256734 260538 256740 260540
rect 191281 260536 193660 260538
rect 191281 260480 191286 260536
rect 191342 260480 193660 260536
rect 191281 260478 193660 260480
rect 253460 260478 256740 260538
rect 191281 260475 191347 260478
rect 256734 260476 256740 260478
rect 256804 260476 256810 260540
rect 66805 260130 66871 260133
rect 147673 260130 147739 260133
rect 173341 260130 173407 260133
rect 66805 260128 68908 260130
rect 66805 260072 66810 260128
rect 66866 260072 68908 260128
rect 66805 260070 68908 260072
rect 147673 260128 173407 260130
rect 147673 260072 147678 260128
rect 147734 260072 173346 260128
rect 173402 260072 173407 260128
rect 147673 260070 173407 260072
rect 66805 260067 66871 260070
rect 147673 260067 147739 260070
rect 173341 260067 173407 260070
rect 101213 259858 101279 259861
rect 98716 259856 101279 259858
rect 98716 259800 101218 259856
rect 101274 259800 101279 259856
rect 98716 259798 101279 259800
rect 253430 259858 253490 260100
rect 262254 259858 262260 259860
rect 253430 259798 262260 259858
rect 101213 259795 101279 259798
rect 262254 259796 262260 259798
rect 262324 259796 262330 259860
rect 255405 259586 255471 259589
rect 253460 259584 255471 259586
rect 253460 259528 255410 259584
rect 255466 259528 255471 259584
rect 253460 259526 255471 259528
rect 255405 259523 255471 259526
rect 46841 258770 46907 258773
rect 64638 258770 64644 258772
rect 46841 258768 64644 258770
rect 46841 258712 46846 258768
rect 46902 258712 64644 258768
rect 46841 258710 64644 258712
rect 46841 258707 46907 258710
rect 64638 258708 64644 258710
rect 64708 258770 64714 258772
rect 68878 258770 68938 259284
rect 100753 259042 100819 259045
rect 98716 259040 100819 259042
rect 98716 258984 100758 259040
rect 100814 258984 100819 259040
rect 98716 258982 100819 258984
rect 100753 258979 100819 258982
rect 193397 258906 193463 258909
rect 193630 258906 193690 259420
rect 255497 259178 255563 259181
rect 253460 259176 255563 259178
rect 253460 259120 255502 259176
rect 255558 259120 255563 259176
rect 253460 259118 255563 259120
rect 255497 259115 255563 259118
rect 193397 258904 193690 258906
rect 193397 258848 193402 258904
rect 193458 258848 193690 258904
rect 193397 258846 193690 258848
rect 582373 258906 582439 258909
rect 583520 258906 584960 258996
rect 582373 258904 584960 258906
rect 582373 258848 582378 258904
rect 582434 258848 584960 258904
rect 582373 258846 584960 258848
rect 193397 258843 193463 258846
rect 582373 258843 582439 258846
rect 64708 258710 68938 258770
rect 64708 258708 64714 258710
rect 111006 258708 111012 258772
rect 111076 258770 111082 258772
rect 129733 258770 129799 258773
rect 185761 258770 185827 258773
rect 111076 258768 185827 258770
rect 111076 258712 129738 258768
rect 129794 258712 185766 258768
rect 185822 258712 185827 258768
rect 583520 258756 584960 258846
rect 111076 258710 185827 258712
rect 111076 258708 111082 258710
rect 129733 258707 129799 258710
rect 185761 258707 185827 258710
rect 253430 258634 253490 258740
rect 263542 258634 263548 258636
rect 253430 258574 263548 258634
rect 263542 258572 263548 258574
rect 263612 258572 263618 258636
rect 66437 258090 66503 258093
rect 66437 258088 66546 258090
rect 66437 258032 66442 258088
rect 66498 258032 66546 258088
rect 66437 258027 66546 258032
rect 66486 257954 66546 258027
rect 67909 257954 67975 257957
rect 68878 257954 68938 258468
rect 100753 258226 100819 258229
rect 98716 258224 100819 258226
rect 98716 258168 100758 258224
rect 100814 258168 100819 258224
rect 98716 258166 100819 258168
rect 100753 258163 100819 258166
rect 178534 258164 178540 258228
rect 178604 258226 178610 258228
rect 253430 258226 253490 258332
rect 262254 258226 262260 258228
rect 178604 258166 193660 258226
rect 253430 258166 262260 258226
rect 178604 258164 178610 258166
rect 262254 258164 262260 258166
rect 262324 258164 262330 258228
rect 255497 257954 255563 257957
rect 66486 257952 68938 257954
rect 66486 257896 67914 257952
rect 67970 257896 68938 257952
rect 66486 257894 68938 257896
rect 253460 257952 255563 257954
rect 253460 257896 255502 257952
rect 255558 257896 255563 257952
rect 253460 257894 255563 257896
rect 67909 257891 67975 257894
rect 255497 257891 255563 257894
rect 66805 257682 66871 257685
rect 66805 257680 68908 257682
rect 66805 257624 66810 257680
rect 66866 257624 68908 257680
rect 66805 257622 68908 257624
rect 66805 257619 66871 257622
rect 100753 257410 100819 257413
rect 259494 257410 259500 257412
rect 98716 257408 100819 257410
rect 98716 257352 100758 257408
rect 100814 257352 100819 257408
rect 98716 257350 100819 257352
rect 253460 257350 259500 257410
rect 100753 257347 100819 257350
rect 259494 257348 259500 257350
rect 259564 257348 259570 257412
rect 138013 257274 138079 257277
rect 180333 257274 180399 257277
rect 138013 257272 180399 257274
rect 138013 257216 138018 257272
rect 138074 257216 180338 257272
rect 180394 257216 180399 257272
rect 138013 257214 180399 257216
rect 138013 257211 138079 257214
rect 180333 257211 180399 257214
rect 267774 257212 267780 257276
rect 267844 257274 267850 257276
rect 268101 257274 268167 257277
rect 267844 257272 268167 257274
rect 267844 257216 268106 257272
rect 268162 257216 268167 257272
rect 267844 257214 268167 257216
rect 267844 257212 267850 257214
rect 268101 257211 268167 257214
rect 191649 257138 191715 257141
rect 191649 257136 193660 257138
rect 191649 257080 191654 257136
rect 191710 257080 193660 257136
rect 191649 257078 193660 257080
rect 191649 257075 191715 257078
rect 255313 257002 255379 257005
rect 253460 257000 255379 257002
rect 253460 256944 255318 257000
rect 255374 256944 255379 257000
rect 253460 256942 255379 256944
rect 255313 256939 255379 256942
rect 66253 256866 66319 256869
rect 66253 256864 68908 256866
rect 66253 256808 66258 256864
rect 66314 256808 68908 256864
rect 66253 256806 68908 256808
rect 66253 256803 66319 256806
rect 99966 256668 99972 256732
rect 100036 256730 100042 256732
rect 100385 256730 100451 256733
rect 100036 256728 100451 256730
rect 100036 256672 100390 256728
rect 100446 256672 100451 256728
rect 100036 256670 100451 256672
rect 100036 256668 100042 256670
rect 100385 256667 100451 256670
rect 255497 256594 255563 256597
rect 253460 256592 255563 256594
rect 66805 256050 66871 256053
rect 98686 256050 98746 256564
rect 253460 256536 255502 256592
rect 255558 256536 255563 256592
rect 253460 256534 255563 256536
rect 255497 256531 255563 256534
rect 255405 256186 255471 256189
rect 253460 256184 255471 256186
rect 253460 256128 255410 256184
rect 255466 256128 255471 256184
rect 253460 256126 255471 256128
rect 255405 256123 255471 256126
rect 66805 256048 68908 256050
rect 66805 255992 66810 256048
rect 66866 255992 68908 256048
rect 66805 255990 68908 255992
rect 98686 255990 103530 256050
rect 66805 255987 66871 255990
rect 101029 255778 101095 255781
rect 98164 255776 101095 255778
rect 98164 255748 101034 255776
rect 98134 255720 101034 255748
rect 101090 255720 101095 255776
rect 98134 255718 101095 255720
rect 98134 255372 98194 255718
rect 101029 255715 101095 255718
rect 98126 255308 98132 255372
rect 98196 255308 98202 255372
rect 103470 255370 103530 255990
rect 146293 255914 146359 255917
rect 169293 255914 169359 255917
rect 146293 255912 169359 255914
rect 146293 255856 146298 255912
rect 146354 255856 169298 255912
rect 169354 255856 169359 255912
rect 146293 255854 169359 255856
rect 146293 255851 146359 255854
rect 169293 255851 169359 255854
rect 190637 255914 190703 255917
rect 190637 255912 193660 255914
rect 190637 255856 190642 255912
rect 190698 255856 193660 255912
rect 190637 255854 193660 255856
rect 190637 255851 190703 255854
rect 253430 255642 253490 255748
rect 269062 255642 269068 255644
rect 253430 255582 269068 255642
rect 269062 255580 269068 255582
rect 269132 255580 269138 255644
rect 146293 255370 146359 255373
rect 103470 255368 146359 255370
rect 103470 255312 146298 255368
rect 146354 255312 146359 255368
rect 103470 255310 146359 255312
rect 146293 255307 146359 255310
rect 255497 255234 255563 255237
rect 253460 255232 255563 255234
rect 68878 254690 68938 255204
rect 253460 255176 255502 255232
rect 255558 255176 255563 255232
rect 253460 255174 255563 255176
rect 255497 255171 255563 255174
rect 100845 254962 100911 254965
rect 98716 254960 100911 254962
rect 98716 254904 100850 254960
rect 100906 254904 100911 254960
rect 98716 254902 100911 254904
rect 100845 254899 100911 254902
rect 191649 254826 191715 254829
rect 258390 254826 258396 254828
rect 191649 254824 193660 254826
rect 191649 254768 191654 254824
rect 191710 254768 193660 254824
rect 191649 254766 193660 254768
rect 253460 254766 258396 254826
rect 191649 254763 191715 254766
rect 258390 254764 258396 254766
rect 258460 254764 258466 254828
rect 64830 254630 68938 254690
rect 35801 254554 35867 254557
rect 35801 254552 45570 254554
rect 35801 254496 35806 254552
rect 35862 254496 45570 254552
rect 35801 254494 45570 254496
rect 35801 254491 35867 254494
rect -960 254146 480 254236
rect 3141 254146 3207 254149
rect -960 254144 3207 254146
rect -960 254088 3146 254144
rect 3202 254088 3207 254144
rect -960 254086 3207 254088
rect 45510 254146 45570 254494
rect 48129 254146 48195 254149
rect 64830 254146 64890 254630
rect 106641 254554 106707 254557
rect 108246 254554 108252 254556
rect 106641 254552 108252 254554
rect 106641 254496 106646 254552
rect 106702 254496 108252 254552
rect 106641 254494 108252 254496
rect 106641 254491 106707 254494
rect 108246 254492 108252 254494
rect 108316 254492 108322 254556
rect 66805 254418 66871 254421
rect 255589 254418 255655 254421
rect 66805 254416 68908 254418
rect 66805 254360 66810 254416
rect 66866 254360 68908 254416
rect 66805 254358 68908 254360
rect 253460 254416 255655 254418
rect 253460 254360 255594 254416
rect 255650 254360 255655 254416
rect 253460 254358 255655 254360
rect 66805 254355 66871 254358
rect 255589 254355 255655 254358
rect 100753 254146 100819 254149
rect 45510 254144 64890 254146
rect 45510 254088 48134 254144
rect 48190 254088 64890 254144
rect 45510 254086 64890 254088
rect 98716 254144 100819 254146
rect 98716 254088 100758 254144
rect 100814 254088 100819 254144
rect 98716 254086 100819 254088
rect -960 253996 480 254086
rect 3141 254083 3207 254086
rect 48129 254083 48195 254086
rect 100753 254083 100819 254086
rect 255405 254010 255471 254013
rect 253460 254008 255471 254010
rect 253460 253952 255410 254008
rect 255466 253952 255471 254008
rect 253460 253950 255471 253952
rect 255405 253947 255471 253950
rect 266302 253948 266308 254012
rect 266372 254010 266378 254012
rect 266721 254010 266787 254013
rect 266372 254008 266787 254010
rect 266372 253952 266726 254008
rect 266782 253952 266787 254008
rect 266372 253950 266787 253952
rect 266372 253948 266378 253950
rect 266721 253947 266787 253950
rect 273294 253948 273300 254012
rect 273364 254010 273370 254012
rect 273621 254010 273687 254013
rect 273364 254008 273687 254010
rect 273364 253952 273626 254008
rect 273682 253952 273687 254008
rect 273364 253950 273687 253952
rect 273364 253948 273370 253950
rect 273621 253947 273687 253950
rect 32397 253874 32463 253877
rect 66662 253874 66668 253876
rect 32397 253872 66668 253874
rect 32397 253816 32402 253872
rect 32458 253816 66668 253872
rect 32397 253814 66668 253816
rect 32397 253811 32463 253814
rect 66662 253812 66668 253814
rect 66732 253874 66738 253876
rect 66732 253814 68938 253874
rect 66732 253812 66738 253814
rect 68878 253572 68938 253814
rect 191649 253602 191715 253605
rect 191649 253600 193660 253602
rect 191649 253544 191654 253600
rect 191710 253544 193660 253600
rect 191649 253542 193660 253544
rect 191649 253539 191715 253542
rect 254710 253466 254716 253468
rect 253460 253406 254716 253466
rect 254710 253404 254716 253406
rect 254780 253404 254786 253468
rect 100753 253330 100819 253333
rect 98716 253328 100819 253330
rect 98716 253272 100758 253328
rect 100814 253272 100819 253328
rect 98716 253270 100819 253272
rect 100753 253267 100819 253270
rect 141049 253194 141115 253197
rect 188286 253194 188292 253196
rect 141049 253192 188292 253194
rect 141049 253136 141054 253192
rect 141110 253136 188292 253192
rect 141049 253134 188292 253136
rect 141049 253131 141115 253134
rect 188286 253132 188292 253134
rect 188356 253132 188362 253196
rect 275277 253194 275343 253197
rect 583477 253194 583543 253197
rect 275277 253192 583543 253194
rect 275277 253136 275282 253192
rect 275338 253136 583482 253192
rect 583538 253136 583543 253192
rect 275277 253134 583543 253136
rect 275277 253131 275343 253134
rect 583477 253131 583543 253134
rect 256141 253058 256207 253061
rect 253460 253056 256207 253058
rect 253460 253000 256146 253056
rect 256202 253000 256207 253056
rect 253460 252998 256207 253000
rect 256141 252995 256207 252998
rect 66069 252786 66135 252789
rect 66529 252786 66595 252789
rect 66069 252784 68908 252786
rect 66069 252728 66074 252784
rect 66130 252728 66534 252784
rect 66590 252728 68908 252784
rect 66069 252726 68908 252728
rect 66069 252723 66135 252726
rect 66529 252723 66595 252726
rect 255405 252650 255471 252653
rect 253460 252648 255471 252650
rect 253460 252592 255410 252648
rect 255466 252592 255471 252648
rect 253460 252590 255471 252592
rect 255405 252587 255471 252590
rect 100845 252514 100911 252517
rect 98716 252512 100911 252514
rect 98716 252456 100850 252512
rect 100906 252456 100911 252512
rect 98716 252454 100911 252456
rect 100845 252451 100911 252454
rect 191649 252514 191715 252517
rect 191649 252512 193660 252514
rect 191649 252456 191654 252512
rect 191710 252456 193660 252512
rect 191649 252454 193660 252456
rect 191649 252451 191715 252454
rect 255589 252242 255655 252245
rect 253460 252240 255655 252242
rect 253460 252184 255594 252240
rect 255650 252184 255655 252240
rect 253460 252182 255655 252184
rect 255589 252179 255655 252182
rect 66253 251970 66319 251973
rect 66253 251968 68908 251970
rect 66253 251912 66258 251968
rect 66314 251912 68908 251968
rect 66253 251910 68908 251912
rect 66253 251907 66319 251910
rect 255405 251834 255471 251837
rect 253460 251832 255471 251834
rect 253460 251776 255410 251832
rect 255466 251776 255471 251832
rect 253460 251774 255471 251776
rect 255405 251771 255471 251774
rect 106181 251698 106247 251701
rect 98716 251696 106247 251698
rect 98716 251640 106186 251696
rect 106242 251640 106247 251696
rect 98716 251638 106247 251640
rect 106181 251635 106247 251638
rect 53741 251290 53807 251293
rect 61009 251290 61075 251293
rect 53741 251288 61075 251290
rect 53741 251232 53746 251288
rect 53802 251232 61014 251288
rect 61070 251232 61075 251288
rect 53741 251230 61075 251232
rect 53741 251227 53807 251230
rect 61009 251227 61075 251230
rect 107469 251290 107535 251293
rect 174629 251290 174695 251293
rect 107469 251288 174695 251290
rect 107469 251232 107474 251288
rect 107530 251232 174634 251288
rect 174690 251232 174695 251288
rect 107469 251230 174695 251232
rect 107469 251227 107535 251230
rect 174629 251227 174695 251230
rect 190821 251290 190887 251293
rect 256233 251290 256299 251293
rect 190821 251288 193660 251290
rect 190821 251232 190826 251288
rect 190882 251232 193660 251288
rect 190821 251230 193660 251232
rect 253460 251288 256299 251290
rect 253460 251232 256238 251288
rect 256294 251232 256299 251288
rect 253460 251230 256299 251232
rect 190821 251227 190887 251230
rect 256233 251227 256299 251230
rect 66805 251154 66871 251157
rect 66805 251152 68908 251154
rect 66805 251096 66810 251152
rect 66866 251096 68908 251152
rect 66805 251094 68908 251096
rect 66805 251091 66871 251094
rect 100753 250882 100819 250885
rect 255497 250882 255563 250885
rect 98716 250880 100819 250882
rect 98716 250824 100758 250880
rect 100814 250824 100819 250880
rect 98716 250822 100819 250824
rect 253460 250880 255563 250882
rect 253460 250824 255502 250880
rect 255558 250824 255563 250880
rect 253460 250822 255563 250824
rect 100753 250819 100819 250822
rect 255497 250819 255563 250822
rect 256049 250474 256115 250477
rect 253460 250472 256115 250474
rect 253460 250416 256054 250472
rect 256110 250416 256115 250472
rect 253460 250414 256115 250416
rect 256049 250411 256115 250414
rect 66897 250338 66963 250341
rect 66897 250336 68908 250338
rect 66897 250280 66902 250336
rect 66958 250280 68908 250336
rect 66897 250278 68908 250280
rect 66897 250275 66963 250278
rect 191649 250202 191715 250205
rect 191649 250200 193660 250202
rect 191649 250144 191654 250200
rect 191710 250144 193660 250200
rect 191649 250142 193660 250144
rect 191649 250139 191715 250142
rect 101949 250066 102015 250069
rect 255405 250066 255471 250069
rect 98716 250064 102015 250066
rect 98716 250008 101954 250064
rect 102010 250008 102015 250064
rect 98716 250006 102015 250008
rect 253460 250064 255471 250066
rect 253460 250008 255410 250064
rect 255466 250008 255471 250064
rect 253460 250006 255471 250008
rect 101949 250003 102015 250006
rect 255405 250003 255471 250006
rect 255313 249522 255379 249525
rect 253460 249520 255379 249522
rect 68878 248978 68938 249492
rect 253460 249464 255318 249520
rect 255374 249464 255379 249520
rect 253460 249462 255379 249464
rect 255313 249459 255379 249462
rect 64830 248918 68938 248978
rect 61837 248570 61903 248573
rect 64830 248570 64890 248918
rect 66805 248706 66871 248709
rect 98686 248706 98746 249220
rect 117221 249114 117287 249117
rect 126329 249114 126395 249117
rect 103470 249112 126395 249114
rect 103470 249056 117226 249112
rect 117282 249056 126334 249112
rect 126390 249056 126395 249112
rect 103470 249054 126395 249056
rect 103470 248706 103530 249054
rect 117221 249051 117287 249054
rect 126329 249051 126395 249054
rect 155401 249114 155467 249117
rect 187049 249114 187115 249117
rect 255405 249114 255471 249117
rect 155401 249112 187115 249114
rect 155401 249056 155406 249112
rect 155462 249056 187054 249112
rect 187110 249056 187115 249112
rect 155401 249054 187115 249056
rect 253460 249112 255471 249114
rect 253460 249056 255410 249112
rect 255466 249056 255471 249112
rect 253460 249054 255471 249056
rect 155401 249051 155467 249054
rect 187049 249051 187115 249054
rect 255405 249051 255471 249054
rect 191649 248978 191715 248981
rect 191649 248976 193660 248978
rect 191649 248920 191654 248976
rect 191710 248920 193660 248976
rect 191649 248918 193660 248920
rect 191649 248915 191715 248918
rect 256417 248706 256483 248709
rect 66805 248704 68908 248706
rect 66805 248648 66810 248704
rect 66866 248648 68908 248704
rect 66805 248646 68908 248648
rect 98686 248646 103530 248706
rect 253460 248704 256483 248706
rect 253460 248648 256422 248704
rect 256478 248648 256483 248704
rect 253460 248646 256483 248648
rect 66805 248643 66871 248646
rect 256417 248643 256483 248646
rect 61837 248568 64890 248570
rect 61837 248512 61842 248568
rect 61898 248512 64890 248568
rect 61837 248510 64890 248512
rect 61837 248507 61903 248510
rect 101673 248434 101739 248437
rect 98716 248432 101739 248434
rect 98716 248376 101678 248432
rect 101734 248376 101739 248432
rect 98716 248374 101739 248376
rect 101673 248371 101739 248374
rect 255589 248434 255655 248437
rect 259678 248434 259684 248436
rect 255589 248432 259684 248434
rect 255589 248376 255594 248432
rect 255650 248376 259684 248432
rect 255589 248374 259684 248376
rect 255589 248371 255655 248374
rect 259678 248372 259684 248374
rect 259748 248372 259754 248436
rect 61929 248300 61995 248301
rect 61878 248298 61884 248300
rect 61838 248238 61884 248298
rect 61948 248296 61995 248300
rect 255405 248298 255471 248301
rect 61990 248240 61995 248296
rect 61878 248236 61884 248238
rect 61948 248236 61995 248240
rect 253460 248296 255471 248298
rect 253460 248240 255410 248296
rect 255466 248240 255471 248296
rect 253460 248238 255471 248240
rect 61929 248235 61995 248236
rect 255405 248235 255471 248238
rect 66897 247890 66963 247893
rect 191649 247890 191715 247893
rect 255313 247890 255379 247893
rect 66897 247888 68908 247890
rect 66897 247832 66902 247888
rect 66958 247832 68908 247888
rect 66897 247830 68908 247832
rect 191649 247888 193660 247890
rect 191649 247832 191654 247888
rect 191710 247832 193660 247888
rect 191649 247830 193660 247832
rect 253460 247888 255379 247890
rect 253460 247832 255318 247888
rect 255374 247832 255379 247888
rect 253460 247830 255379 247832
rect 66897 247827 66963 247830
rect 191649 247827 191715 247830
rect 255313 247827 255379 247830
rect 99189 247618 99255 247621
rect 98164 247616 99255 247618
rect 98164 247588 99194 247616
rect 98134 247560 99194 247588
rect 99250 247560 99255 247616
rect 98134 247558 99255 247560
rect 98134 247077 98194 247558
rect 99189 247555 99255 247558
rect 173341 247618 173407 247621
rect 193254 247618 193260 247620
rect 173341 247616 193260 247618
rect 173341 247560 173346 247616
rect 173402 247560 193260 247616
rect 173341 247558 193260 247560
rect 173341 247555 173407 247558
rect 193254 247556 193260 247558
rect 193324 247556 193330 247620
rect 258257 247346 258323 247349
rect 253460 247344 258323 247346
rect 253460 247288 258262 247344
rect 258318 247288 258323 247344
rect 253460 247286 258323 247288
rect 258257 247283 258323 247286
rect 67173 247074 67239 247077
rect 67357 247074 67423 247077
rect 67173 247072 68908 247074
rect 67173 247016 67178 247072
rect 67234 247016 67362 247072
rect 67418 247016 68908 247072
rect 67173 247014 68908 247016
rect 98085 247072 98194 247077
rect 98085 247016 98090 247072
rect 98146 247016 98194 247072
rect 98085 247014 98194 247016
rect 256141 247074 256207 247077
rect 258390 247074 258396 247076
rect 256141 247072 258396 247074
rect 256141 247016 256146 247072
rect 256202 247016 258396 247072
rect 256141 247014 258396 247016
rect 67173 247011 67239 247014
rect 67357 247011 67423 247014
rect 98085 247011 98151 247014
rect 256141 247011 256207 247014
rect 258390 247012 258396 247014
rect 258460 247012 258466 247076
rect 255405 246938 255471 246941
rect 253460 246936 255471 246938
rect 253460 246880 255410 246936
rect 255466 246880 255471 246936
rect 253460 246878 255471 246880
rect 255405 246875 255471 246878
rect 101029 246802 101095 246805
rect 98716 246800 101095 246802
rect 98716 246744 101034 246800
rect 101090 246744 101095 246800
rect 98716 246742 101095 246744
rect 101029 246739 101095 246742
rect 190637 246666 190703 246669
rect 190637 246664 193660 246666
rect 190637 246608 190642 246664
rect 190698 246608 193660 246664
rect 190637 246606 193660 246608
rect 190637 246603 190703 246606
rect 255681 246530 255747 246533
rect 253460 246528 255747 246530
rect 253460 246472 255686 246528
rect 255742 246472 255747 246528
rect 253460 246470 255747 246472
rect 255681 246467 255747 246470
rect 67357 246258 67423 246261
rect 67357 246256 68908 246258
rect 67357 246200 67362 246256
rect 67418 246200 68908 246256
rect 67357 246198 68908 246200
rect 67357 246195 67423 246198
rect 256785 246122 256851 246125
rect 253460 246120 256851 246122
rect 253460 246064 256790 246120
rect 256846 246064 256851 246120
rect 253460 246062 256851 246064
rect 256785 246059 256851 246062
rect 101121 245986 101187 245989
rect 98716 245984 101187 245986
rect 98716 245928 101126 245984
rect 101182 245928 101187 245984
rect 98716 245926 101187 245928
rect 101121 245923 101187 245926
rect 102409 245714 102475 245717
rect 103421 245714 103487 245717
rect 112621 245714 112687 245717
rect 102409 245712 112687 245714
rect 102409 245656 102414 245712
rect 102470 245656 103426 245712
rect 103482 245656 112626 245712
rect 112682 245656 112687 245712
rect 102409 245654 112687 245656
rect 102409 245651 102475 245654
rect 103421 245651 103487 245654
rect 112621 245651 112687 245654
rect 254761 245578 254827 245581
rect 253460 245576 254827 245578
rect 68878 244898 68938 245412
rect 102317 245170 102383 245173
rect 98716 245168 102383 245170
rect 98716 245112 102322 245168
rect 102378 245112 102383 245168
rect 98716 245110 102383 245112
rect 102317 245107 102383 245110
rect 64830 244838 68938 244898
rect 57697 244490 57763 244493
rect 57881 244490 57947 244493
rect 64830 244490 64890 244838
rect 67541 244626 67607 244629
rect 189809 244626 189875 244629
rect 193630 244626 193690 245548
rect 253460 245520 254766 245576
rect 254822 245520 254827 245576
rect 253460 245518 254827 245520
rect 254761 245515 254827 245518
rect 582465 245578 582531 245581
rect 583520 245578 584960 245668
rect 582465 245576 584960 245578
rect 582465 245520 582470 245576
rect 582526 245520 584960 245576
rect 582465 245518 584960 245520
rect 582465 245515 582531 245518
rect 583520 245428 584960 245518
rect 255497 245170 255563 245173
rect 253460 245168 255563 245170
rect 253460 245112 255502 245168
rect 255558 245112 255563 245168
rect 253460 245110 255563 245112
rect 255497 245107 255563 245110
rect 67541 244624 69092 244626
rect 67541 244568 67546 244624
rect 67602 244596 69092 244624
rect 189809 244624 193690 244626
rect 67602 244568 69122 244596
rect 67541 244566 69122 244568
rect 67541 244563 67607 244566
rect 57697 244488 64890 244490
rect 57697 244432 57702 244488
rect 57758 244432 57886 244488
rect 57942 244432 64890 244488
rect 57697 244430 64890 244432
rect 57697 244427 57763 244430
rect 57881 244427 57947 244430
rect 69062 244357 69122 244566
rect 189809 244568 189814 244624
rect 189870 244568 193690 244624
rect 189809 244566 193690 244568
rect 253430 244626 253490 244732
rect 253430 244566 258090 244626
rect 189809 244563 189875 244566
rect 69013 244352 69122 244357
rect 102409 244354 102475 244357
rect 69013 244296 69018 244352
rect 69074 244296 69122 244352
rect 69013 244294 69122 244296
rect 98716 244352 102475 244354
rect 98716 244296 102414 244352
rect 102470 244296 102475 244352
rect 98716 244294 102475 244296
rect 69013 244291 69079 244294
rect 102409 244291 102475 244294
rect 168966 244292 168972 244356
rect 169036 244354 169042 244356
rect 255405 244354 255471 244357
rect 169036 244294 193660 244354
rect 253460 244352 255471 244354
rect 253460 244296 255410 244352
rect 255466 244296 255471 244352
rect 253460 244294 255471 244296
rect 258030 244354 258090 244566
rect 269205 244354 269271 244357
rect 258030 244352 269271 244354
rect 258030 244296 269210 244352
rect 269266 244296 269271 244352
rect 258030 244294 269271 244296
rect 169036 244292 169042 244294
rect 255405 244291 255471 244294
rect 269205 244291 269271 244294
rect 259678 244156 259684 244220
rect 259748 244218 259754 244220
rect 574737 244218 574803 244221
rect 259748 244216 574803 244218
rect 259748 244160 574742 244216
rect 574798 244160 574803 244216
rect 259748 244158 574803 244160
rect 259748 244156 259754 244158
rect 574737 244155 574803 244158
rect 66253 243810 66319 243813
rect 66253 243808 68908 243810
rect 66253 243752 66258 243808
rect 66314 243752 68908 243808
rect 66253 243750 68908 243752
rect 66253 243747 66319 243750
rect 252878 243676 252938 243916
rect 252870 243612 252876 243676
rect 252940 243612 252946 243676
rect 102225 243538 102291 243541
rect 98716 243536 102291 243538
rect 98716 243480 102230 243536
rect 102286 243480 102291 243536
rect 98716 243478 102291 243480
rect 102225 243475 102291 243478
rect 115289 243538 115355 243541
rect 122925 243538 122991 243541
rect 115289 243536 122991 243538
rect 115289 243480 115294 243536
rect 115350 243480 122930 243536
rect 122986 243480 122991 243536
rect 115289 243478 122991 243480
rect 115289 243475 115355 243478
rect 122925 243475 122991 243478
rect 254117 243402 254183 243405
rect 253460 243400 254183 243402
rect 253460 243344 254122 243400
rect 254178 243344 254183 243400
rect 253460 243342 254183 243344
rect 254117 243339 254183 243342
rect 41229 242994 41295 242997
rect 57094 242994 57100 242996
rect 41229 242992 57100 242994
rect 41229 242936 41234 242992
rect 41290 242936 57100 242992
rect 41229 242934 57100 242936
rect 41229 242931 41295 242934
rect 57094 242932 57100 242934
rect 57164 242994 57170 242996
rect 57830 242994 57836 242996
rect 57164 242934 57836 242994
rect 57164 242932 57170 242934
rect 57830 242932 57836 242934
rect 57900 242932 57906 242996
rect 66805 242994 66871 242997
rect 189901 242994 189967 242997
rect 193630 242994 193690 243236
rect 66805 242992 68908 242994
rect 66805 242936 66810 242992
rect 66866 242936 68908 242992
rect 66805 242934 68908 242936
rect 189901 242992 193690 242994
rect 189901 242936 189906 242992
rect 189962 242936 193690 242992
rect 189901 242934 193690 242936
rect 66805 242931 66871 242934
rect 189901 242931 189967 242934
rect 252878 242861 252938 242964
rect 193254 242796 193260 242860
rect 193324 242858 193330 242860
rect 193581 242858 193647 242861
rect 193324 242856 193647 242858
rect 193324 242800 193586 242856
rect 193642 242800 193647 242856
rect 193324 242798 193647 242800
rect 252878 242856 252987 242861
rect 252878 242800 252926 242856
rect 252982 242800 252987 242856
rect 252878 242798 252987 242800
rect 193324 242796 193330 242798
rect 193581 242795 193647 242798
rect 252921 242795 252987 242798
rect 101029 242722 101095 242725
rect 98716 242720 101095 242722
rect 98716 242664 101034 242720
rect 101090 242664 101095 242720
rect 98716 242662 101095 242664
rect 101029 242659 101095 242662
rect 99557 242586 99623 242589
rect 99966 242586 99972 242588
rect 99557 242584 99972 242586
rect 99557 242528 99562 242584
rect 99618 242528 99972 242584
rect 99557 242526 99972 242528
rect 99557 242523 99623 242526
rect 99966 242524 99972 242526
rect 100036 242524 100042 242588
rect 100109 242586 100175 242589
rect 110689 242586 110755 242589
rect 100109 242584 110755 242586
rect 100109 242528 100114 242584
rect 100170 242528 110694 242584
rect 110750 242528 110755 242584
rect 100109 242526 110755 242528
rect 100109 242523 100175 242526
rect 110689 242523 110755 242526
rect 253062 242453 253122 242556
rect 253013 242448 253122 242453
rect 253013 242392 253018 242448
rect 253074 242392 253122 242448
rect 253013 242390 253122 242392
rect 253013 242387 253079 242390
rect 144269 242178 144335 242181
rect 192886 242178 192892 242180
rect 144269 242176 192892 242178
rect 62113 241634 62179 241637
rect 63401 241634 63467 241637
rect 68878 241634 68938 242148
rect 144269 242120 144274 242176
rect 144330 242120 192892 242176
rect 144269 242118 192892 242120
rect 144269 242115 144335 242118
rect 192886 242116 192892 242118
rect 192956 242116 192962 242180
rect 107469 241906 107535 241909
rect 98716 241904 107535 241906
rect 98716 241848 107474 241904
rect 107530 241848 107535 241904
rect 98716 241846 107535 241848
rect 107469 241843 107535 241846
rect 69473 241770 69539 241773
rect 70945 241772 71011 241773
rect 70158 241770 70164 241772
rect 69473 241768 70164 241770
rect 69473 241712 69478 241768
rect 69534 241712 70164 241768
rect 69473 241710 70164 241712
rect 69473 241707 69539 241710
rect 70158 241708 70164 241710
rect 70228 241708 70234 241772
rect 70894 241708 70900 241772
rect 70964 241770 71011 241772
rect 72325 241772 72391 241773
rect 72325 241770 72372 241772
rect 70964 241768 71056 241770
rect 71006 241712 71056 241768
rect 70964 241710 71056 241712
rect 72280 241768 72372 241770
rect 72280 241712 72330 241768
rect 72280 241710 72372 241712
rect 70964 241708 71011 241710
rect 70945 241707 71011 241708
rect 72325 241708 72372 241710
rect 72436 241708 72442 241772
rect 73470 241708 73476 241772
rect 73540 241770 73546 241772
rect 73889 241770 73955 241773
rect 83365 241772 83431 241773
rect 83365 241770 83412 241772
rect 73540 241768 73955 241770
rect 73540 241712 73894 241768
rect 73950 241712 73955 241768
rect 73540 241710 73955 241712
rect 83320 241768 83412 241770
rect 83320 241712 83370 241768
rect 83320 241710 83412 241712
rect 73540 241708 73546 241710
rect 72325 241707 72391 241708
rect 73889 241707 73955 241710
rect 83365 241708 83412 241710
rect 83476 241708 83482 241772
rect 84694 241708 84700 241772
rect 84764 241770 84770 241772
rect 84929 241770 84995 241773
rect 84764 241768 84995 241770
rect 84764 241712 84934 241768
rect 84990 241712 84995 241768
rect 84764 241710 84995 241712
rect 84764 241708 84770 241710
rect 83365 241707 83431 241708
rect 84929 241707 84995 241710
rect 85941 241770 86007 241773
rect 86677 241772 86743 241773
rect 88057 241772 88123 241773
rect 86166 241770 86172 241772
rect 85941 241768 86172 241770
rect 85941 241712 85946 241768
rect 86002 241712 86172 241768
rect 85941 241710 86172 241712
rect 85941 241707 86007 241710
rect 86166 241708 86172 241710
rect 86236 241708 86242 241772
rect 86677 241770 86724 241772
rect 86632 241768 86724 241770
rect 86632 241712 86682 241768
rect 86632 241710 86724 241712
rect 86677 241708 86724 241710
rect 86788 241708 86794 241772
rect 88006 241708 88012 241772
rect 88076 241770 88123 241772
rect 96429 241770 96495 241773
rect 100109 241770 100175 241773
rect 88076 241768 88168 241770
rect 88118 241712 88168 241768
rect 88076 241710 88168 241712
rect 96429 241768 100175 241770
rect 96429 241712 96434 241768
rect 96490 241712 100114 241768
rect 100170 241712 100175 241768
rect 96429 241710 100175 241712
rect 88076 241708 88123 241710
rect 86677 241707 86743 241708
rect 88057 241707 88123 241708
rect 96429 241707 96495 241710
rect 100109 241707 100175 241710
rect 70025 241636 70091 241637
rect 62113 241632 68938 241634
rect 62113 241576 62118 241632
rect 62174 241576 63406 241632
rect 63462 241576 68938 241632
rect 62113 241574 68938 241576
rect 62113 241571 62179 241574
rect 63401 241571 63467 241574
rect 69974 241572 69980 241636
rect 70044 241634 70091 241636
rect 70044 241632 70136 241634
rect 70086 241576 70136 241632
rect 70044 241574 70136 241576
rect 70044 241572 70091 241574
rect 72918 241572 72924 241636
rect 72988 241634 72994 241636
rect 75545 241634 75611 241637
rect 72988 241632 75611 241634
rect 72988 241576 75550 241632
rect 75606 241576 75611 241632
rect 72988 241574 75611 241576
rect 72988 241572 72994 241574
rect 70025 241571 70091 241572
rect 75545 241571 75611 241574
rect 91318 241572 91324 241636
rect 91388 241634 91394 241636
rect 92105 241634 92171 241637
rect 91388 241632 92171 241634
rect 91388 241576 92110 241632
rect 92166 241576 92171 241632
rect 91388 241574 92171 241576
rect 91388 241572 91394 241574
rect 92105 241571 92171 241574
rect 103421 241634 103487 241637
rect 115197 241634 115263 241637
rect 162117 241634 162183 241637
rect 103421 241632 103898 241634
rect 103421 241576 103426 241632
rect 103482 241576 103898 241632
rect 103421 241574 103898 241576
rect 103421 241571 103487 241574
rect 92887 241498 92953 241501
rect 103838 241498 103898 241574
rect 115197 241632 162183 241634
rect 115197 241576 115202 241632
rect 115258 241576 162122 241632
rect 162178 241576 162183 241632
rect 115197 241574 162183 241576
rect 115197 241571 115263 241574
rect 162117 241571 162183 241574
rect 188337 241634 188403 241637
rect 193630 241634 193690 242148
rect 252878 242042 252938 242148
rect 252510 241982 252938 242042
rect 188337 241632 193690 241634
rect 188337 241576 188342 241632
rect 188398 241576 193690 241632
rect 188337 241574 193690 241576
rect 251817 241634 251883 241637
rect 252510 241634 252570 241982
rect 284293 241770 284359 241773
rect 253460 241768 284359 241770
rect 253460 241712 284298 241768
rect 284354 241712 284359 241768
rect 253460 241710 284359 241712
rect 284293 241707 284359 241710
rect 251817 241632 252570 241634
rect 251817 241576 251822 241632
rect 251878 241576 252570 241632
rect 251817 241574 252570 241576
rect 188337 241571 188403 241574
rect 251817 241571 251883 241574
rect 104934 241498 104940 241500
rect 92887 241496 103714 241498
rect 92887 241440 92892 241496
rect 92948 241440 103714 241496
rect 92887 241438 103714 241440
rect 103838 241438 104940 241498
rect 92887 241435 92953 241438
rect 57830 241300 57836 241364
rect 57900 241362 57906 241364
rect 71037 241362 71103 241365
rect 57900 241360 71103 241362
rect 57900 241304 71042 241360
rect 71098 241304 71103 241360
rect 57900 241302 71103 241304
rect 57900 241300 57906 241302
rect 71037 241299 71103 241302
rect 81341 241362 81407 241365
rect 83958 241362 83964 241364
rect 81341 241360 83964 241362
rect 81341 241304 81346 241360
rect 81402 241304 83964 241360
rect 81341 241302 83964 241304
rect 81341 241299 81407 241302
rect 83958 241300 83964 241302
rect 84028 241300 84034 241364
rect 97717 241362 97783 241365
rect 103421 241362 103487 241365
rect 97717 241360 103487 241362
rect 97717 241304 97722 241360
rect 97778 241304 103426 241360
rect 103482 241304 103487 241360
rect 97717 241302 103487 241304
rect 103654 241362 103714 241438
rect 104934 241436 104940 241438
rect 105004 241436 105010 241500
rect 193070 241436 193076 241500
rect 193140 241498 193146 241500
rect 195973 241498 196039 241501
rect 275277 241498 275343 241501
rect 193140 241496 196039 241498
rect 193140 241440 195978 241496
rect 196034 241440 196039 241496
rect 193140 241438 196039 241440
rect 193140 241436 193146 241438
rect 195973 241435 196039 241438
rect 267690 241496 275343 241498
rect 267690 241440 275282 241496
rect 275338 241440 275343 241496
rect 267690 241438 275343 241440
rect 111006 241362 111012 241364
rect 103654 241302 111012 241362
rect 97717 241299 97783 241302
rect 103421 241299 103487 241302
rect 111006 241300 111012 241302
rect 111076 241300 111082 241364
rect 18689 241226 18755 241229
rect 93117 241226 93183 241229
rect 18689 241224 93183 241226
rect -960 241090 480 241180
rect 18689 241168 18694 241224
rect 18750 241168 93122 241224
rect 93178 241168 93183 241224
rect 18689 241166 93183 241168
rect 18689 241163 18755 241166
rect 93117 241163 93183 241166
rect 3509 241090 3575 241093
rect -960 241088 3575 241090
rect -960 241032 3514 241088
rect 3570 241032 3575 241088
rect -960 241030 3575 241032
rect -960 240940 480 241030
rect 3509 241027 3575 241030
rect 192886 240892 192892 240956
rect 192956 240954 192962 240956
rect 215937 240954 216003 240957
rect 258349 240954 258415 240957
rect 192956 240952 258415 240954
rect 192956 240896 215942 240952
rect 215998 240896 258354 240952
rect 258410 240896 258415 240952
rect 192956 240894 258415 240896
rect 192956 240892 192962 240894
rect 215937 240891 216003 240894
rect 258349 240891 258415 240894
rect 71497 240818 71563 240821
rect 176561 240818 176627 240821
rect 258390 240818 258396 240820
rect 71497 240816 258396 240818
rect 71497 240760 71502 240816
rect 71558 240760 176566 240816
rect 176622 240760 258396 240816
rect 71497 240758 258396 240760
rect 71497 240755 71563 240758
rect 176561 240755 176627 240758
rect 258390 240756 258396 240758
rect 258460 240818 258466 240820
rect 267690 240818 267750 241438
rect 275277 241435 275343 241438
rect 258460 240758 267750 240818
rect 258460 240756 258466 240758
rect 198641 240274 198707 240277
rect 201534 240274 201540 240276
rect 198641 240272 201540 240274
rect 198641 240216 198646 240272
rect 198702 240216 201540 240272
rect 198641 240214 201540 240216
rect 198641 240211 198707 240214
rect 201534 240212 201540 240214
rect 201604 240212 201610 240276
rect 79685 240138 79751 240141
rect 82077 240138 82143 240141
rect 64830 240136 82143 240138
rect 64830 240080 79690 240136
rect 79746 240080 82082 240136
rect 82138 240080 82143 240136
rect 64830 240078 82143 240080
rect 64597 240002 64663 240005
rect 64830 240002 64890 240078
rect 79685 240075 79751 240078
rect 82077 240075 82143 240078
rect 84285 240138 84351 240141
rect 84694 240138 84700 240140
rect 84285 240136 84700 240138
rect 84285 240080 84290 240136
rect 84346 240080 84700 240136
rect 84285 240078 84700 240080
rect 84285 240075 84351 240078
rect 84694 240076 84700 240078
rect 84764 240076 84770 240140
rect 91502 240076 91508 240140
rect 91572 240138 91578 240140
rect 91645 240138 91711 240141
rect 91572 240136 91711 240138
rect 91572 240080 91650 240136
rect 91706 240080 91711 240136
rect 91572 240078 91711 240080
rect 91572 240076 91578 240078
rect 91645 240075 91711 240078
rect 94313 240138 94379 240141
rect 94865 240138 94931 240141
rect 94998 240138 95004 240140
rect 94313 240136 95004 240138
rect 94313 240080 94318 240136
rect 94374 240080 94870 240136
rect 94926 240080 95004 240136
rect 94313 240078 95004 240080
rect 94313 240075 94379 240078
rect 94865 240075 94931 240078
rect 94998 240076 95004 240078
rect 95068 240076 95074 240140
rect 96797 240138 96863 240141
rect 215385 240140 215451 240141
rect 97758 240138 97764 240140
rect 96797 240136 97764 240138
rect 96797 240080 96802 240136
rect 96858 240080 97764 240136
rect 96797 240078 97764 240080
rect 96797 240075 96863 240078
rect 97758 240076 97764 240078
rect 97828 240076 97834 240140
rect 215334 240138 215340 240140
rect 215294 240078 215340 240138
rect 215404 240136 215451 240140
rect 222377 240138 222443 240141
rect 223481 240138 223547 240141
rect 215446 240080 215451 240136
rect 215334 240076 215340 240078
rect 215404 240076 215451 240080
rect 215385 240075 215451 240076
rect 219390 240136 223547 240138
rect 219390 240080 222382 240136
rect 222438 240080 223486 240136
rect 223542 240080 223547 240136
rect 219390 240078 223547 240080
rect 64597 240000 64890 240002
rect 64597 239944 64602 240000
rect 64658 239944 64890 240000
rect 64597 239942 64890 239944
rect 64597 239939 64663 239942
rect 72550 239940 72556 240004
rect 72620 240002 72626 240004
rect 72877 240002 72943 240005
rect 72620 240000 72943 240002
rect 72620 239944 72882 240000
rect 72938 239944 72943 240000
rect 72620 239942 72943 239944
rect 72620 239940 72626 239942
rect 52269 239866 52335 239869
rect 72558 239866 72618 239940
rect 72877 239939 72943 239942
rect 86861 240002 86927 240005
rect 219390 240002 219450 240078
rect 222377 240075 222443 240078
rect 223481 240075 223547 240078
rect 234705 240138 234771 240141
rect 234838 240138 234844 240140
rect 234705 240136 234844 240138
rect 234705 240080 234710 240136
rect 234766 240080 234844 240136
rect 234705 240078 234844 240080
rect 234705 240075 234771 240078
rect 234838 240076 234844 240078
rect 234908 240076 234914 240140
rect 235993 240138 236059 240141
rect 236678 240138 236684 240140
rect 235993 240136 236684 240138
rect 235993 240080 235998 240136
rect 236054 240080 236684 240136
rect 235993 240078 236684 240080
rect 235993 240075 236059 240078
rect 236678 240076 236684 240078
rect 236748 240076 236754 240140
rect 251909 240138 251975 240141
rect 254710 240138 254716 240140
rect 251909 240136 254716 240138
rect 251909 240080 251914 240136
rect 251970 240080 254716 240136
rect 251909 240078 254716 240080
rect 251909 240075 251975 240078
rect 254710 240076 254716 240078
rect 254780 240138 254786 240140
rect 583293 240138 583359 240141
rect 254780 240136 583359 240138
rect 254780 240080 583298 240136
rect 583354 240080 583359 240136
rect 254780 240078 583359 240080
rect 254780 240076 254786 240078
rect 583293 240075 583359 240078
rect 86861 240000 219450 240002
rect 86861 239944 86866 240000
rect 86922 239944 219450 240000
rect 86861 239942 219450 239944
rect 86861 239939 86927 239942
rect 52269 239864 72618 239866
rect 52269 239808 52274 239864
rect 52330 239808 72618 239864
rect 52269 239806 72618 239808
rect 89621 239866 89687 239869
rect 128537 239866 128603 239869
rect 215334 239866 215340 239868
rect 89621 239864 215340 239866
rect 89621 239808 89626 239864
rect 89682 239808 128542 239864
rect 128598 239808 215340 239864
rect 89621 239806 215340 239808
rect 52269 239803 52335 239806
rect 89621 239803 89687 239806
rect 128537 239803 128603 239806
rect 215334 239804 215340 239806
rect 215404 239804 215410 239868
rect 90265 239730 90331 239733
rect 90950 239730 90956 239732
rect 90265 239728 90956 239730
rect 90265 239672 90270 239728
rect 90326 239672 90956 239728
rect 90265 239670 90956 239672
rect 90265 239667 90331 239670
rect 90950 239668 90956 239670
rect 91020 239730 91026 239732
rect 227713 239730 227779 239733
rect 228357 239730 228423 239733
rect 91020 239728 228423 239730
rect 91020 239672 227718 239728
rect 227774 239672 228362 239728
rect 228418 239672 228423 239728
rect 91020 239670 228423 239672
rect 91020 239668 91026 239670
rect 227713 239667 227779 239670
rect 228357 239667 228423 239670
rect 245009 239594 245075 239597
rect 256734 239594 256740 239596
rect 245009 239592 256740 239594
rect 245009 239536 245014 239592
rect 245070 239536 256740 239592
rect 245009 239534 256740 239536
rect 245009 239531 245075 239534
rect 256734 239532 256740 239534
rect 256804 239532 256810 239596
rect 231117 239458 231183 239461
rect 252502 239458 252508 239460
rect 231117 239456 252508 239458
rect 231117 239400 231122 239456
rect 231178 239400 252508 239456
rect 231117 239398 252508 239400
rect 231117 239395 231183 239398
rect 252502 239396 252508 239398
rect 252572 239396 252578 239460
rect 238702 238716 238708 238780
rect 238772 238778 238778 238780
rect 238845 238778 238911 238781
rect 238772 238776 238911 238778
rect 238772 238720 238850 238776
rect 238906 238720 238911 238776
rect 238772 238718 238911 238720
rect 238772 238716 238778 238718
rect 238845 238715 238911 238718
rect 256969 238778 257035 238781
rect 259678 238778 259684 238780
rect 256969 238776 259684 238778
rect 256969 238720 256974 238776
rect 257030 238720 259684 238776
rect 256969 238718 259684 238720
rect 256969 238715 257035 238718
rect 259678 238716 259684 238718
rect 259748 238716 259754 238780
rect 67909 238642 67975 238645
rect 115381 238642 115447 238645
rect 67909 238640 115447 238642
rect 67909 238584 67914 238640
rect 67970 238584 115386 238640
rect 115442 238584 115447 238640
rect 67909 238582 115447 238584
rect 67909 238579 67975 238582
rect 115381 238579 115447 238582
rect 178677 238642 178743 238645
rect 222101 238642 222167 238645
rect 583661 238642 583727 238645
rect 178677 238640 222167 238642
rect 178677 238584 178682 238640
rect 178738 238584 222106 238640
rect 222162 238584 222167 238640
rect 178677 238582 222167 238584
rect 178677 238579 178743 238582
rect 222101 238579 222167 238582
rect 277350 238640 583727 238642
rect 277350 238584 583666 238640
rect 583722 238584 583727 238640
rect 277350 238582 583727 238584
rect 95049 238506 95115 238509
rect 106365 238506 106431 238509
rect 95049 238504 106431 238506
rect 95049 238448 95054 238504
rect 95110 238448 106370 238504
rect 106426 238448 106431 238504
rect 95049 238446 106431 238448
rect 95049 238443 95115 238446
rect 106365 238443 106431 238446
rect 156689 238506 156755 238509
rect 268009 238506 268075 238509
rect 156689 238504 268075 238506
rect 156689 238448 156694 238504
rect 156750 238448 268014 238504
rect 268070 238448 268075 238504
rect 156689 238446 268075 238448
rect 156689 238443 156755 238446
rect 268009 238443 268075 238446
rect 93710 238172 93716 238236
rect 93780 238234 93786 238236
rect 95049 238234 95115 238237
rect 93780 238232 95115 238234
rect 93780 238176 95054 238232
rect 95110 238176 95115 238232
rect 93780 238174 95115 238176
rect 93780 238172 93786 238174
rect 95049 238171 95115 238174
rect 52361 238098 52427 238101
rect 74717 238098 74783 238101
rect 52361 238096 74783 238098
rect 52361 238040 52366 238096
rect 52422 238040 74722 238096
rect 74778 238040 74783 238096
rect 52361 238038 74783 238040
rect 52361 238035 52427 238038
rect 74717 238035 74783 238038
rect 222837 238098 222903 238101
rect 242014 238098 242020 238100
rect 222837 238096 242020 238098
rect 222837 238040 222842 238096
rect 222898 238040 242020 238096
rect 222837 238038 242020 238040
rect 222837 238035 222903 238038
rect 242014 238036 242020 238038
rect 242084 238036 242090 238100
rect 254577 238098 254643 238101
rect 262254 238098 262260 238100
rect 254577 238096 262260 238098
rect 254577 238040 254582 238096
rect 254638 238040 262260 238096
rect 254577 238038 262260 238040
rect 254577 238035 254643 238038
rect 262254 238036 262260 238038
rect 262324 238098 262330 238100
rect 277350 238098 277410 238582
rect 583661 238579 583727 238582
rect 262324 238038 277410 238098
rect 262324 238036 262330 238038
rect 64638 237900 64644 237964
rect 64708 237962 64714 237964
rect 157241 237962 157307 237965
rect 64708 237960 157307 237962
rect 64708 237904 157246 237960
rect 157302 237904 157307 237960
rect 64708 237902 157307 237904
rect 64708 237900 64714 237902
rect 157241 237899 157307 237902
rect 195237 237962 195303 237965
rect 241513 237962 241579 237965
rect 256049 237962 256115 237965
rect 195237 237960 256115 237962
rect 195237 237904 195242 237960
rect 195298 237904 241518 237960
rect 241574 237904 256054 237960
rect 256110 237904 256115 237960
rect 195237 237902 256115 237904
rect 195237 237899 195303 237902
rect 241513 237899 241579 237902
rect 256049 237899 256115 237902
rect 95233 237282 95299 237285
rect 198774 237282 198780 237284
rect 95233 237280 198780 237282
rect 95233 237224 95238 237280
rect 95294 237224 198780 237280
rect 95233 237222 198780 237224
rect 95233 237219 95299 237222
rect 198774 237220 198780 237222
rect 198844 237220 198850 237284
rect 103605 237146 103671 237149
rect 84150 237144 103671 237146
rect 84150 237088 103610 237144
rect 103666 237088 103671 237144
rect 84150 237086 103671 237088
rect 79961 236874 80027 236877
rect 84150 236874 84210 237086
rect 103605 237083 103671 237086
rect 159449 237146 159515 237149
rect 159909 237146 159975 237149
rect 261017 237146 261083 237149
rect 159449 237144 261083 237146
rect 159449 237088 159454 237144
rect 159510 237088 159914 237144
rect 159970 237088 261022 237144
rect 261078 237088 261083 237144
rect 159449 237086 261083 237088
rect 159449 237083 159515 237086
rect 159909 237083 159975 237086
rect 261017 237083 261083 237086
rect 93761 237010 93827 237013
rect 95182 237010 95188 237012
rect 93761 237008 95188 237010
rect 93761 236952 93766 237008
rect 93822 236952 95188 237008
rect 93761 236950 95188 236952
rect 93761 236947 93827 236950
rect 95182 236948 95188 236950
rect 95252 236948 95258 237012
rect 79961 236872 84210 236874
rect 79961 236816 79966 236872
rect 80022 236816 84210 236872
rect 79961 236814 84210 236816
rect 79961 236811 80027 236814
rect 85573 236602 85639 236605
rect 108941 236602 109007 236605
rect 85573 236600 109007 236602
rect 85573 236544 85578 236600
rect 85634 236544 108946 236600
rect 109002 236544 109007 236600
rect 85573 236542 109007 236544
rect 85573 236539 85639 236542
rect 108941 236539 109007 236542
rect 203977 236602 204043 236605
rect 582465 236602 582531 236605
rect 203977 236600 582531 236602
rect 203977 236544 203982 236600
rect 204038 236544 582470 236600
rect 582526 236544 582531 236600
rect 203977 236542 582531 236544
rect 203977 236539 204043 236542
rect 582465 236539 582531 236542
rect 21357 236058 21423 236061
rect 76833 236058 76899 236061
rect 21357 236056 76899 236058
rect 21357 236000 21362 236056
rect 21418 236000 76838 236056
rect 76894 236000 76899 236056
rect 21357 235998 76899 236000
rect 21357 235995 21423 235998
rect 76833 235995 76899 235998
rect 78673 236058 78739 236061
rect 79961 236058 80027 236061
rect 78673 236056 80027 236058
rect 78673 236000 78678 236056
rect 78734 236000 79966 236056
rect 80022 236000 80027 236056
rect 78673 235998 80027 236000
rect 78673 235995 78739 235998
rect 79961 235995 80027 235998
rect 84193 235922 84259 235925
rect 122833 235922 122899 235925
rect 84193 235920 122899 235922
rect 84193 235864 84198 235920
rect 84254 235864 122838 235920
rect 122894 235864 122899 235920
rect 84193 235862 122899 235864
rect 84193 235859 84259 235862
rect 122790 235859 122899 235862
rect 205541 235922 205607 235925
rect 210366 235922 210372 235924
rect 205541 235920 210372 235922
rect 205541 235864 205546 235920
rect 205602 235864 210372 235920
rect 205541 235862 210372 235864
rect 205541 235859 205607 235862
rect 210366 235860 210372 235862
rect 210436 235860 210442 235924
rect 269062 235922 269068 235924
rect 258030 235862 269068 235922
rect 91001 235786 91067 235789
rect 92606 235786 92612 235788
rect 91001 235784 92612 235786
rect 91001 235728 91006 235784
rect 91062 235728 92612 235784
rect 91001 235726 92612 235728
rect 91001 235723 91067 235726
rect 92606 235724 92612 235726
rect 92676 235724 92682 235788
rect 122790 235514 122850 235859
rect 180149 235650 180215 235653
rect 161430 235648 180215 235650
rect 161430 235592 180154 235648
rect 180210 235592 180215 235648
rect 161430 235590 180215 235592
rect 161430 235514 161490 235590
rect 180149 235587 180215 235590
rect 122790 235454 161490 235514
rect 179413 235514 179479 235517
rect 195237 235514 195303 235517
rect 179413 235512 195303 235514
rect 179413 235456 179418 235512
rect 179474 235456 195242 235512
rect 195298 235456 195303 235512
rect 179413 235454 195303 235456
rect 179413 235451 179479 235454
rect 195237 235451 195303 235454
rect 256049 235514 256115 235517
rect 258030 235514 258090 235862
rect 269062 235860 269068 235862
rect 269132 235922 269138 235924
rect 582925 235922 582991 235925
rect 269132 235920 582991 235922
rect 269132 235864 582930 235920
rect 582986 235864 582991 235920
rect 269132 235862 582991 235864
rect 269132 235860 269138 235862
rect 582925 235859 582991 235862
rect 256049 235512 258090 235514
rect 256049 235456 256054 235512
rect 256110 235456 258090 235512
rect 256049 235454 258090 235456
rect 256049 235451 256115 235454
rect 160921 235378 160987 235381
rect 259729 235378 259795 235381
rect 160921 235376 259795 235378
rect 160921 235320 160926 235376
rect 160982 235320 259734 235376
rect 259790 235320 259795 235376
rect 160921 235318 259795 235320
rect 160921 235315 160987 235318
rect 259729 235315 259795 235318
rect 15101 235242 15167 235245
rect 189901 235242 189967 235245
rect 15101 235240 189967 235242
rect 15101 235184 15106 235240
rect 15162 235184 189906 235240
rect 189962 235184 189967 235240
rect 15101 235182 189967 235184
rect 15101 235179 15167 235182
rect 189901 235179 189967 235182
rect 196617 235242 196683 235245
rect 233233 235242 233299 235245
rect 266302 235242 266308 235244
rect 196617 235240 266308 235242
rect 196617 235184 196622 235240
rect 196678 235184 233238 235240
rect 233294 235184 266308 235240
rect 196617 235182 266308 235184
rect 196617 235179 196683 235182
rect 233233 235179 233299 235182
rect 266302 235180 266308 235182
rect 266372 235180 266378 235244
rect 100017 234562 100083 234565
rect 102225 234562 102291 234565
rect 125726 234562 125732 234564
rect 100017 234560 125732 234562
rect 100017 234504 100022 234560
rect 100078 234504 102230 234560
rect 102286 234504 125732 234560
rect 100017 234502 125732 234504
rect 100017 234499 100083 234502
rect 102225 234499 102291 234502
rect 125726 234500 125732 234502
rect 125796 234562 125802 234564
rect 261109 234562 261175 234565
rect 125796 234560 261175 234562
rect 125796 234504 261114 234560
rect 261170 234504 261175 234560
rect 125796 234502 261175 234504
rect 125796 234500 125802 234502
rect 261109 234499 261175 234502
rect 88333 234426 88399 234429
rect 105629 234426 105695 234429
rect 88333 234424 105695 234426
rect 88333 234368 88338 234424
rect 88394 234368 105634 234424
rect 105690 234368 105695 234424
rect 88333 234366 105695 234368
rect 88333 234363 88399 234366
rect 105629 234363 105695 234366
rect 227805 234426 227871 234429
rect 228214 234426 228220 234428
rect 227805 234424 228220 234426
rect 227805 234368 227810 234424
rect 227866 234368 228220 234424
rect 227805 234366 228220 234368
rect 227805 234363 227871 234366
rect 228214 234364 228220 234366
rect 228284 234426 228290 234428
rect 267774 234426 267780 234428
rect 228284 234366 267780 234426
rect 228284 234364 228290 234366
rect 267774 234364 267780 234366
rect 267844 234364 267850 234428
rect 180333 234018 180399 234021
rect 220997 234018 221063 234021
rect 180333 234016 221063 234018
rect 180333 233960 180338 234016
rect 180394 233960 221002 234016
rect 221058 233960 221063 234016
rect 180333 233958 221063 233960
rect 180333 233955 180399 233958
rect 220997 233955 221063 233958
rect 184197 233882 184263 233885
rect 207105 233882 207171 233885
rect 256877 233882 256943 233885
rect 184197 233880 256943 233882
rect 184197 233824 184202 233880
rect 184258 233824 207110 233880
rect 207166 233824 256882 233880
rect 256938 233824 256943 233880
rect 184197 233822 256943 233824
rect 184197 233819 184263 233822
rect 207105 233819 207171 233822
rect 256877 233819 256943 233822
rect 18597 233474 18663 233477
rect 97257 233474 97323 233477
rect 97717 233474 97783 233477
rect 18597 233472 97783 233474
rect 18597 233416 18602 233472
rect 18658 233416 97262 233472
rect 97318 233416 97722 233472
rect 97778 233416 97783 233472
rect 18597 233414 97783 233416
rect 18597 233411 18663 233414
rect 97257 233411 97323 233414
rect 97717 233411 97783 233414
rect 67633 233338 67699 233341
rect 170581 233338 170647 233341
rect 67633 233336 170647 233338
rect 67633 233280 67638 233336
rect 67694 233280 170586 233336
rect 170642 233280 170647 233336
rect 67633 233278 170647 233280
rect 67633 233275 67699 233278
rect 170581 233275 170647 233278
rect 118693 233202 118759 233205
rect 209814 233202 209820 233204
rect 118693 233200 209820 233202
rect 118693 233144 118698 233200
rect 118754 233144 209820 233200
rect 118693 233142 209820 233144
rect 118693 233139 118759 233142
rect 209814 233140 209820 233142
rect 209884 233202 209890 233204
rect 211061 233202 211127 233205
rect 209884 233200 211127 233202
rect 209884 233144 211066 233200
rect 211122 233144 211127 233200
rect 209884 233142 211127 233144
rect 209884 233140 209890 233142
rect 211061 233139 211127 233142
rect 162209 232658 162275 232661
rect 234613 232658 234679 232661
rect 162209 232656 234679 232658
rect 162209 232600 162214 232656
rect 162270 232600 234618 232656
rect 234674 232600 234679 232656
rect 162209 232598 234679 232600
rect 162209 232595 162275 232598
rect 234613 232595 234679 232598
rect 28901 232522 28967 232525
rect 187233 232522 187299 232525
rect 28901 232520 187299 232522
rect 28901 232464 28906 232520
rect 28962 232464 187238 232520
rect 187294 232464 187299 232520
rect 28901 232462 187299 232464
rect 28901 232459 28967 232462
rect 187233 232459 187299 232462
rect 190361 232522 190427 232525
rect 582925 232522 582991 232525
rect 190361 232520 582991 232522
rect 190361 232464 190366 232520
rect 190422 232464 582930 232520
rect 582986 232464 582991 232520
rect 190361 232462 582991 232464
rect 190361 232459 190427 232462
rect 582925 232459 582991 232462
rect 580165 232386 580231 232389
rect 583520 232386 584960 232476
rect 580165 232384 584960 232386
rect 580165 232328 580170 232384
rect 580226 232328 584960 232384
rect 580165 232326 584960 232328
rect 580165 232323 580231 232326
rect 583520 232236 584960 232326
rect 50889 231842 50955 231845
rect 263961 231842 264027 231845
rect 50889 231840 264027 231842
rect 50889 231784 50894 231840
rect 50950 231784 263966 231840
rect 264022 231784 264027 231840
rect 50889 231782 264027 231784
rect 50889 231779 50955 231782
rect 263961 231779 264027 231782
rect 195830 231100 195836 231164
rect 195900 231162 195906 231164
rect 254526 231162 254532 231164
rect 195900 231102 254532 231162
rect 195900 231100 195906 231102
rect 254526 231100 254532 231102
rect 254596 231100 254602 231164
rect 68870 230556 68876 230620
rect 68940 230618 68946 230620
rect 74533 230618 74599 230621
rect 68940 230616 74599 230618
rect 68940 230560 74538 230616
rect 74594 230560 74599 230616
rect 68940 230558 74599 230560
rect 68940 230556 68946 230558
rect 74533 230555 74599 230558
rect 157241 230482 157307 230485
rect 262489 230482 262555 230485
rect 157241 230480 262555 230482
rect 157241 230424 157246 230480
rect 157302 230424 262494 230480
rect 262550 230424 262555 230480
rect 157241 230422 262555 230424
rect 157241 230419 157307 230422
rect 262489 230419 262555 230422
rect 68001 229938 68067 229941
rect 128997 229938 129063 229941
rect 68001 229936 129063 229938
rect 68001 229880 68006 229936
rect 68062 229880 129002 229936
rect 129058 229880 129063 229936
rect 68001 229878 129063 229880
rect 68001 229875 68067 229878
rect 128997 229875 129063 229878
rect 108297 229802 108363 229805
rect 234705 229802 234771 229805
rect 108297 229800 234771 229802
rect 108297 229744 108302 229800
rect 108358 229744 234710 229800
rect 234766 229744 234771 229800
rect 108297 229742 234771 229744
rect 108297 229739 108363 229742
rect 234705 229739 234771 229742
rect 59169 228986 59235 228989
rect 115197 228986 115263 228989
rect 59169 228984 115263 228986
rect 59169 228928 59174 228984
rect 59230 228928 115202 228984
rect 115258 228928 115263 228984
rect 59169 228926 115263 228928
rect 59169 228923 59235 228926
rect 115197 228923 115263 228926
rect 140129 228986 140195 228989
rect 251909 228986 251975 228989
rect 140129 228984 251975 228986
rect 140129 228928 140134 228984
rect 140190 228928 251914 228984
rect 251970 228928 251975 228984
rect 140129 228926 251975 228928
rect 140129 228923 140195 228926
rect 251909 228923 251975 228926
rect 192477 228850 192543 228853
rect 208485 228850 208551 228853
rect 192477 228848 208551 228850
rect 192477 228792 192482 228848
rect 192538 228792 208490 228848
rect 208546 228792 208551 228848
rect 192477 228790 208551 228792
rect 192477 228787 192543 228790
rect 208485 228787 208551 228790
rect -960 227884 480 228124
rect 208485 227762 208551 227765
rect 208710 227762 208716 227764
rect 208485 227760 208716 227762
rect 208485 227704 208490 227760
rect 208546 227704 208716 227760
rect 208485 227702 208716 227704
rect 208485 227699 208551 227702
rect 208710 227700 208716 227702
rect 208780 227700 208786 227764
rect 251173 227762 251239 227765
rect 251909 227762 251975 227765
rect 251173 227760 251975 227762
rect 251173 227704 251178 227760
rect 251234 227704 251914 227760
rect 251970 227704 251975 227760
rect 251173 227702 251975 227704
rect 251173 227699 251239 227702
rect 251909 227699 251975 227702
rect 186221 227626 186287 227629
rect 277577 227626 277643 227629
rect 186221 227624 277643 227626
rect 186221 227568 186226 227624
rect 186282 227568 277582 227624
rect 277638 227568 277643 227624
rect 186221 227566 277643 227568
rect 186221 227563 186287 227566
rect 277577 227563 277643 227566
rect 212073 227082 212139 227085
rect 223614 227082 223620 227084
rect 212073 227080 223620 227082
rect 212073 227024 212078 227080
rect 212134 227024 223620 227080
rect 212073 227022 223620 227024
rect 212073 227019 212139 227022
rect 223614 227020 223620 227022
rect 223684 227020 223690 227084
rect 13721 226946 13787 226949
rect 220854 226946 220860 226948
rect 13721 226944 220860 226946
rect 13721 226888 13726 226944
rect 13782 226888 220860 226944
rect 13721 226886 220860 226888
rect 13721 226883 13787 226886
rect 220854 226884 220860 226886
rect 220924 226884 220930 226948
rect 223573 226538 223639 226541
rect 224350 226538 224356 226540
rect 223573 226536 224356 226538
rect 223573 226480 223578 226536
rect 223634 226480 224356 226536
rect 223573 226478 224356 226480
rect 223573 226475 223639 226478
rect 224350 226476 224356 226478
rect 224420 226476 224426 226540
rect 65926 226340 65932 226404
rect 65996 226402 66002 226404
rect 66161 226402 66227 226405
rect 171869 226402 171935 226405
rect 65996 226400 171935 226402
rect 65996 226344 66166 226400
rect 66222 226344 171874 226400
rect 171930 226344 171935 226400
rect 65996 226342 171935 226344
rect 65996 226340 66002 226342
rect 66161 226339 66227 226342
rect 171869 226339 171935 226342
rect 118785 226266 118851 226269
rect 259494 226266 259500 226268
rect 118785 226264 259500 226266
rect 118785 226208 118790 226264
rect 118846 226208 259500 226264
rect 118785 226206 259500 226208
rect 118785 226203 118851 226206
rect 259494 226204 259500 226206
rect 259564 226204 259570 226268
rect 162117 226130 162183 226133
rect 273294 226130 273300 226132
rect 162117 226128 273300 226130
rect 162117 226072 162122 226128
rect 162178 226072 273300 226128
rect 162117 226070 273300 226072
rect 162117 226067 162183 226070
rect 273294 226068 273300 226070
rect 273364 226068 273370 226132
rect 115749 225042 115815 225045
rect 118785 225042 118851 225045
rect 115749 225040 118851 225042
rect 115749 224984 115754 225040
rect 115810 224984 118790 225040
rect 118846 224984 118851 225040
rect 115749 224982 118851 224984
rect 115749 224979 115815 224982
rect 118785 224979 118851 224982
rect 162117 225042 162183 225045
rect 162761 225042 162827 225045
rect 162117 225040 162827 225042
rect 162117 224984 162122 225040
rect 162178 224984 162766 225040
rect 162822 224984 162827 225040
rect 162117 224982 162827 224984
rect 162117 224979 162183 224982
rect 162761 224979 162827 224982
rect 193765 224362 193831 224365
rect 252461 224362 252527 224365
rect 193765 224360 252527 224362
rect 193765 224304 193770 224360
rect 193826 224304 252466 224360
rect 252522 224304 252527 224360
rect 193765 224302 252527 224304
rect 193765 224299 193831 224302
rect 252461 224299 252527 224302
rect 29637 224226 29703 224229
rect 223573 224226 223639 224229
rect 29637 224224 223639 224226
rect 29637 224168 29642 224224
rect 29698 224168 223578 224224
rect 223634 224168 223639 224224
rect 29637 224166 223639 224168
rect 29637 224163 29703 224166
rect 223573 224163 223639 224166
rect 51993 223546 52059 223549
rect 52269 223546 52335 223549
rect 51993 223544 52335 223546
rect 51993 223488 51998 223544
rect 52054 223488 52274 223544
rect 52330 223488 52335 223544
rect 51993 223486 52335 223488
rect 51993 223483 52059 223486
rect 52269 223483 52335 223486
rect 153193 223546 153259 223549
rect 201534 223546 201540 223548
rect 153193 223544 201540 223546
rect 153193 223488 153198 223544
rect 153254 223488 201540 223544
rect 153193 223486 201540 223488
rect 153193 223483 153259 223486
rect 201534 223484 201540 223486
rect 201604 223546 201610 223548
rect 202781 223546 202847 223549
rect 201604 223544 202847 223546
rect 201604 223488 202786 223544
rect 202842 223488 202847 223544
rect 201604 223486 202847 223488
rect 201604 223484 201610 223486
rect 202781 223483 202847 223486
rect 186129 223002 186195 223005
rect 256049 223002 256115 223005
rect 186129 223000 256115 223002
rect 186129 222944 186134 223000
rect 186190 222944 256054 223000
rect 256110 222944 256115 223000
rect 186129 222942 256115 222944
rect 186129 222939 186195 222942
rect 256049 222939 256115 222942
rect 35801 222866 35867 222869
rect 224166 222866 224172 222868
rect 35801 222864 224172 222866
rect 35801 222808 35806 222864
rect 35862 222808 224172 222864
rect 35801 222806 224172 222808
rect 35801 222803 35867 222806
rect 224166 222804 224172 222806
rect 224236 222804 224242 222868
rect 52269 222322 52335 222325
rect 186129 222322 186195 222325
rect 52269 222320 186195 222322
rect 52269 222264 52274 222320
rect 52330 222264 186134 222320
rect 186190 222264 186195 222320
rect 52269 222262 186195 222264
rect 52269 222259 52335 222262
rect 186129 222259 186195 222262
rect 108246 221580 108252 221644
rect 108316 221642 108322 221644
rect 244273 221642 244339 221645
rect 108316 221640 244339 221642
rect 108316 221584 244278 221640
rect 244334 221584 244339 221640
rect 108316 221582 244339 221584
rect 108316 221580 108322 221582
rect 244273 221579 244339 221582
rect 24761 221506 24827 221509
rect 189809 221506 189875 221509
rect 24761 221504 189875 221506
rect 24761 221448 24766 221504
rect 24822 221448 189814 221504
rect 189870 221448 189875 221504
rect 24761 221446 189875 221448
rect 24761 221443 24827 221446
rect 189809 221443 189875 221446
rect 196617 221506 196683 221509
rect 255446 221506 255452 221508
rect 196617 221504 255452 221506
rect 196617 221448 196622 221504
rect 196678 221448 255452 221504
rect 196617 221446 255452 221448
rect 196617 221443 196683 221446
rect 255446 221444 255452 221446
rect 255516 221444 255522 221508
rect 263542 220826 263548 220828
rect 122790 220766 263548 220826
rect 112437 220282 112503 220285
rect 120717 220282 120783 220285
rect 122790 220282 122850 220766
rect 263542 220764 263548 220766
rect 263612 220764 263618 220828
rect 112437 220280 122850 220282
rect 112437 220224 112442 220280
rect 112498 220224 120722 220280
rect 120778 220224 122850 220280
rect 112437 220222 122850 220224
rect 112437 220219 112503 220222
rect 120717 220219 120783 220222
rect 115841 220146 115907 220149
rect 217174 220146 217180 220148
rect 115841 220144 217180 220146
rect 115841 220088 115846 220144
rect 115902 220088 217180 220144
rect 115841 220086 217180 220088
rect 115841 220083 115907 220086
rect 217174 220084 217180 220086
rect 217244 220084 217250 220148
rect 182909 219330 182975 219333
rect 265065 219330 265131 219333
rect 182909 219328 265131 219330
rect 182909 219272 182914 219328
rect 182970 219272 265070 219328
rect 265126 219272 265131 219328
rect 182909 219270 265131 219272
rect 182909 219267 182975 219270
rect 265065 219267 265131 219270
rect 582373 219058 582439 219061
rect 583520 219058 584960 219148
rect 582373 219056 584960 219058
rect 582373 219000 582378 219056
rect 582434 219000 584960 219056
rect 582373 218998 584960 219000
rect 582373 218995 582439 218998
rect 583520 218908 584960 218998
rect 42701 218650 42767 218653
rect 226558 218650 226564 218652
rect 42701 218648 226564 218650
rect 42701 218592 42706 218648
rect 42762 218592 226564 218648
rect 42701 218590 226564 218592
rect 42701 218587 42767 218590
rect 226558 218588 226564 218590
rect 226628 218588 226634 218652
rect 182909 218106 182975 218109
rect 183461 218106 183527 218109
rect 182909 218104 183527 218106
rect 182909 218048 182914 218104
rect 182970 218048 183466 218104
rect 183522 218048 183527 218104
rect 182909 218046 183527 218048
rect 182909 218043 182975 218046
rect 183461 218043 183527 218046
rect 175181 217426 175247 217429
rect 256141 217426 256207 217429
rect 175181 217424 256207 217426
rect 175181 217368 175186 217424
rect 175242 217368 256146 217424
rect 256202 217368 256207 217424
rect 175181 217366 256207 217368
rect 175181 217363 175247 217366
rect 256141 217363 256207 217366
rect 49509 217290 49575 217293
rect 226742 217290 226748 217292
rect 49509 217288 226748 217290
rect 49509 217232 49514 217288
rect 49570 217232 226748 217288
rect 49509 217230 226748 217232
rect 49509 217227 49575 217230
rect 226742 217228 226748 217230
rect 226812 217228 226818 217292
rect 61929 216748 61995 216749
rect 61878 216746 61884 216748
rect 61802 216686 61884 216746
rect 61948 216746 61995 216748
rect 175181 216746 175247 216749
rect 61948 216744 175247 216746
rect 61990 216688 175186 216744
rect 175242 216688 175247 216744
rect 61878 216684 61884 216686
rect 61948 216686 175247 216688
rect 61948 216684 61995 216686
rect 61929 216683 61995 216684
rect 175181 216683 175247 216686
rect 111609 216066 111675 216069
rect 215886 216066 215892 216068
rect 111609 216064 215892 216066
rect 111609 216008 111614 216064
rect 111670 216008 215892 216064
rect 111609 216006 215892 216008
rect 111609 216003 111675 216006
rect 215886 216004 215892 216006
rect 215956 216004 215962 216068
rect 72918 215868 72924 215932
rect 72988 215930 72994 215932
rect 269205 215930 269271 215933
rect 72988 215928 269271 215930
rect 72988 215872 269210 215928
rect 269266 215872 269271 215928
rect 72988 215870 269271 215872
rect 72988 215868 72994 215870
rect 269205 215867 269271 215870
rect -960 214978 480 215068
rect 3417 214978 3483 214981
rect -960 214976 3483 214978
rect -960 214920 3422 214976
rect 3478 214920 3483 214976
rect -960 214918 3483 214920
rect -960 214828 480 214918
rect 3417 214915 3483 214918
rect 117221 214570 117287 214573
rect 238150 214570 238156 214572
rect 117221 214568 238156 214570
rect 117221 214512 117226 214568
rect 117282 214512 238156 214568
rect 117221 214510 238156 214512
rect 117221 214507 117287 214510
rect 238150 214508 238156 214510
rect 238220 214508 238226 214572
rect 76557 214026 76623 214029
rect 181529 214026 181595 214029
rect 76557 214024 181595 214026
rect 76557 213968 76562 214024
rect 76618 213968 181534 214024
rect 181590 213968 181595 214024
rect 76557 213966 181595 213968
rect 76557 213963 76623 213966
rect 181529 213963 181595 213966
rect 232497 213482 232563 213485
rect 248454 213482 248460 213484
rect 232497 213480 248460 213482
rect 232497 213424 232502 213480
rect 232558 213424 248460 213480
rect 232497 213422 248460 213424
rect 232497 213419 232563 213422
rect 248454 213420 248460 213422
rect 248524 213420 248530 213484
rect 184790 213284 184796 213348
rect 184860 213346 184866 213348
rect 255262 213346 255268 213348
rect 184860 213286 255268 213346
rect 184860 213284 184866 213286
rect 255262 213284 255268 213286
rect 255332 213284 255338 213348
rect 106917 213210 106983 213213
rect 236494 213210 236500 213212
rect 106917 213208 236500 213210
rect 106917 213152 106922 213208
rect 106978 213152 236500 213208
rect 106917 213150 236500 213152
rect 106917 213147 106983 213150
rect 236494 213148 236500 213150
rect 236564 213148 236570 213212
rect 57697 212666 57763 212669
rect 184790 212666 184796 212668
rect 57697 212664 184796 212666
rect 57697 212608 57702 212664
rect 57758 212608 184796 212664
rect 57697 212606 184796 212608
rect 57697 212603 57763 212606
rect 184790 212604 184796 212606
rect 184860 212604 184866 212668
rect 188286 212468 188292 212532
rect 188356 212530 188362 212532
rect 288525 212530 288591 212533
rect 188356 212528 288591 212530
rect 188356 212472 288530 212528
rect 288586 212472 288591 212528
rect 188356 212470 288591 212472
rect 188356 212468 188362 212470
rect 288525 212467 288591 212470
rect 19241 211850 19307 211853
rect 222326 211850 222332 211852
rect 19241 211848 222332 211850
rect 19241 211792 19246 211848
rect 19302 211792 222332 211848
rect 19241 211790 222332 211792
rect 19241 211787 19307 211790
rect 222326 211788 222332 211790
rect 222396 211788 222402 211852
rect 55029 211170 55095 211173
rect 188838 211170 188844 211172
rect 55029 211168 188844 211170
rect 55029 211112 55034 211168
rect 55090 211112 188844 211168
rect 55029 211110 188844 211112
rect 55029 211107 55095 211110
rect 188838 211108 188844 211110
rect 188908 211170 188914 211172
rect 191833 211170 191899 211173
rect 230473 211170 230539 211173
rect 231117 211170 231183 211173
rect 188908 211168 191899 211170
rect 188908 211112 191838 211168
rect 191894 211112 191899 211168
rect 188908 211110 191899 211112
rect 188908 211108 188914 211110
rect 191833 211107 191899 211110
rect 219390 211168 231183 211170
rect 219390 211112 230478 211168
rect 230534 211112 231122 211168
rect 231178 211112 231183 211168
rect 219390 211110 231183 211112
rect 92381 211034 92447 211037
rect 219390 211034 219450 211110
rect 230473 211107 230539 211110
rect 231117 211107 231183 211110
rect 249701 211170 249767 211173
rect 256785 211170 256851 211173
rect 249701 211168 256851 211170
rect 249701 211112 249706 211168
rect 249762 211112 256790 211168
rect 256846 211112 256851 211168
rect 249701 211110 256851 211112
rect 249701 211107 249767 211110
rect 256785 211107 256851 211110
rect 92381 211032 219450 211034
rect 92381 210976 92386 211032
rect 92442 210976 219450 211032
rect 92381 210974 219450 210976
rect 92381 210971 92447 210974
rect 45461 210354 45527 210357
rect 219934 210354 219940 210356
rect 45461 210352 219940 210354
rect 45461 210296 45466 210352
rect 45522 210296 219940 210352
rect 45461 210294 219940 210296
rect 45461 210291 45527 210294
rect 219934 210292 219940 210294
rect 220004 210292 220010 210356
rect 181529 209674 181595 209677
rect 182081 209674 182147 209677
rect 278865 209674 278931 209677
rect 181529 209672 278931 209674
rect 181529 209616 181534 209672
rect 181590 209616 182086 209672
rect 182142 209616 278870 209672
rect 278926 209616 278931 209672
rect 181529 209614 278931 209616
rect 181529 209611 181595 209614
rect 182081 209611 182147 209614
rect 278865 209611 278931 209614
rect 69657 208450 69723 208453
rect 71630 208450 71636 208452
rect 69657 208448 71636 208450
rect 69657 208392 69662 208448
rect 69718 208392 71636 208448
rect 69657 208390 71636 208392
rect 69657 208387 69723 208390
rect 71630 208388 71636 208390
rect 71700 208450 71706 208452
rect 190310 208450 190316 208452
rect 71700 208390 190316 208450
rect 71700 208388 71706 208390
rect 190310 208388 190316 208390
rect 190380 208450 190386 208452
rect 200757 208450 200823 208453
rect 190380 208448 200823 208450
rect 190380 208392 200762 208448
rect 200818 208392 200823 208448
rect 190380 208390 200823 208392
rect 190380 208388 190386 208390
rect 200757 208387 200823 208390
rect 224902 207634 224908 207636
rect 219390 207574 224908 207634
rect 97206 207028 97212 207092
rect 97276 207090 97282 207092
rect 219390 207090 219450 207574
rect 224902 207572 224908 207574
rect 224972 207634 224978 207636
rect 263777 207634 263843 207637
rect 224972 207632 263843 207634
rect 224972 207576 263782 207632
rect 263838 207576 263843 207632
rect 224972 207574 263843 207576
rect 224972 207572 224978 207574
rect 263777 207571 263843 207574
rect 97276 207030 219450 207090
rect 224953 207090 225019 207093
rect 226006 207090 226012 207092
rect 224953 207088 226012 207090
rect 224953 207032 224958 207088
rect 225014 207032 226012 207088
rect 224953 207030 226012 207032
rect 97276 207028 97282 207030
rect 224953 207027 225019 207030
rect 226006 207028 226012 207030
rect 226076 207028 226082 207092
rect 80697 206410 80763 206413
rect 105629 206410 105695 206413
rect 80697 206408 105695 206410
rect 80697 206352 80702 206408
rect 80758 206352 105634 206408
rect 105690 206352 105695 206408
rect 80697 206350 105695 206352
rect 80697 206347 80763 206350
rect 105629 206347 105695 206350
rect 48221 206274 48287 206277
rect 207054 206274 207060 206276
rect 48221 206272 207060 206274
rect 48221 206216 48226 206272
rect 48282 206216 207060 206272
rect 48221 206214 207060 206216
rect 48221 206211 48287 206214
rect 207054 206212 207060 206214
rect 207124 206212 207130 206276
rect 213177 206274 213243 206277
rect 245694 206274 245700 206276
rect 213177 206272 245700 206274
rect 213177 206216 213182 206272
rect 213238 206216 245700 206272
rect 213177 206214 245700 206216
rect 213177 206211 213243 206214
rect 245694 206212 245700 206214
rect 245764 206212 245770 206276
rect 104985 205730 105051 205733
rect 105629 205730 105695 205733
rect 203190 205730 203196 205732
rect 104985 205728 203196 205730
rect 104985 205672 104990 205728
rect 105046 205672 105634 205728
rect 105690 205672 203196 205728
rect 104985 205670 203196 205672
rect 104985 205667 105051 205670
rect 105629 205667 105695 205670
rect 203190 205668 203196 205670
rect 203260 205668 203266 205732
rect 580257 205730 580323 205733
rect 583520 205730 584960 205820
rect 580257 205728 584960 205730
rect 580257 205672 580262 205728
rect 580318 205672 584960 205728
rect 580257 205670 584960 205672
rect 580257 205667 580323 205670
rect 583520 205580 584960 205670
rect 41321 204914 41387 204917
rect 204846 204914 204852 204916
rect 41321 204912 204852 204914
rect 41321 204856 41326 204912
rect 41382 204856 204852 204912
rect 41321 204854 204852 204856
rect 41321 204851 41387 204854
rect 204846 204852 204852 204854
rect 204916 204852 204922 204916
rect 68870 203492 68876 203556
rect 68940 203554 68946 203556
rect 82854 203554 82860 203556
rect 68940 203494 82860 203554
rect 68940 203492 68946 203494
rect 82854 203492 82860 203494
rect 82924 203492 82930 203556
rect 104801 203554 104867 203557
rect 214414 203554 214420 203556
rect 104801 203552 214420 203554
rect 104801 203496 104806 203552
rect 104862 203496 214420 203552
rect 104801 203494 214420 203496
rect 104801 203491 104867 203494
rect 214414 203492 214420 203494
rect 214484 203492 214490 203556
rect 203190 202812 203196 202876
rect 203260 202874 203266 202876
rect 258717 202874 258783 202877
rect 203260 202872 258783 202874
rect 203260 202816 258722 202872
rect 258778 202816 258783 202872
rect 203260 202814 258783 202816
rect 203260 202812 203266 202814
rect 258717 202811 258783 202814
rect 144821 202194 144887 202197
rect 196566 202194 196572 202196
rect 144821 202192 196572 202194
rect 144821 202136 144826 202192
rect 144882 202136 196572 202192
rect 144821 202134 196572 202136
rect 144821 202131 144887 202134
rect 196566 202132 196572 202134
rect 196636 202132 196642 202196
rect -960 201922 480 202012
rect 3325 201922 3391 201925
rect -960 201920 3391 201922
rect -960 201864 3330 201920
rect 3386 201864 3391 201920
rect -960 201862 3391 201864
rect -960 201772 480 201862
rect 3325 201859 3391 201862
rect 45369 199338 45435 199341
rect 205766 199338 205772 199340
rect 45369 199336 205772 199338
rect 45369 199280 45374 199336
rect 45430 199280 205772 199336
rect 45369 199278 205772 199280
rect 45369 199275 45435 199278
rect 205766 199276 205772 199278
rect 205836 199276 205842 199340
rect 105486 196692 105492 196756
rect 105556 196754 105562 196756
rect 232078 196754 232084 196756
rect 105556 196694 232084 196754
rect 105556 196692 105562 196694
rect 232078 196692 232084 196694
rect 232148 196692 232154 196756
rect 5441 196618 5507 196621
rect 194542 196618 194548 196620
rect 5441 196616 194548 196618
rect 5441 196560 5446 196616
rect 5502 196560 194548 196616
rect 5441 196558 194548 196560
rect 5441 196555 5507 196558
rect 194542 196556 194548 196558
rect 194612 196556 194618 196620
rect 204846 193972 204852 194036
rect 204916 194034 204922 194036
rect 251214 194034 251220 194036
rect 204916 193974 251220 194034
rect 204916 193972 204922 193974
rect 251214 193972 251220 193974
rect 251284 193972 251290 194036
rect 149697 193898 149763 193901
rect 208526 193898 208532 193900
rect 149697 193896 208532 193898
rect 149697 193840 149702 193896
rect 149758 193840 208532 193896
rect 149697 193838 208532 193840
rect 149697 193835 149763 193838
rect 208526 193836 208532 193838
rect 208596 193836 208602 193900
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 3509 188866 3575 188869
rect -960 188864 3575 188866
rect -960 188808 3514 188864
rect 3570 188808 3575 188864
rect -960 188806 3575 188808
rect -960 188716 480 188806
rect 3509 188803 3575 188806
rect 201350 186900 201356 186964
rect 201420 186962 201426 186964
rect 240910 186962 240916 186964
rect 201420 186902 240916 186962
rect 201420 186900 201426 186902
rect 240910 186900 240916 186902
rect 240980 186900 240986 186964
rect 65374 184180 65380 184244
rect 65444 184242 65450 184244
rect 229686 184242 229692 184244
rect 65444 184182 229692 184242
rect 65444 184180 65450 184182
rect 229686 184180 229692 184182
rect 229756 184180 229762 184244
rect 193857 181386 193923 181389
rect 247718 181386 247724 181388
rect 193857 181384 247724 181386
rect 193857 181328 193862 181384
rect 193918 181328 247724 181384
rect 193857 181326 247724 181328
rect 193857 181323 193923 181326
rect 247718 181324 247724 181326
rect 247788 181324 247794 181388
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect 180149 178666 180215 178669
rect 218646 178666 218652 178668
rect 180149 178664 218652 178666
rect 180149 178608 180154 178664
rect 180210 178608 218652 178664
rect 180149 178606 218652 178608
rect 180149 178603 180215 178606
rect 218646 178604 218652 178606
rect 218716 178604 218722 178668
rect 87822 177244 87828 177308
rect 87892 177306 87898 177308
rect 213177 177306 213243 177309
rect 87892 177304 213243 177306
rect 87892 177248 213182 177304
rect 213238 177248 213243 177304
rect 87892 177246 213243 177248
rect 87892 177244 87898 177246
rect 213177 177243 213243 177246
rect 87597 176762 87663 176765
rect 87822 176762 87828 176764
rect 87597 176760 87828 176762
rect 87597 176704 87602 176760
rect 87658 176704 87828 176760
rect 87597 176702 87828 176704
rect 87597 176699 87663 176702
rect 87822 176700 87828 176702
rect 87892 176700 87898 176764
rect -960 175796 480 176036
rect 52085 175402 52151 175405
rect 197997 175402 198063 175405
rect 52085 175400 198063 175402
rect 52085 175344 52090 175400
rect 52146 175344 198002 175400
rect 198058 175344 198063 175400
rect 52085 175342 198063 175344
rect 52085 175339 52151 175342
rect 197997 175339 198063 175342
rect 88977 174042 89043 174045
rect 214557 174042 214623 174045
rect 88977 174040 214623 174042
rect 88977 173984 88982 174040
rect 89038 173984 214562 174040
rect 214618 173984 214623 174040
rect 88977 173982 214623 173984
rect 88977 173979 89043 173982
rect 214557 173979 214623 173982
rect 206369 173906 206435 173909
rect 207054 173906 207060 173908
rect 206369 173904 207060 173906
rect 206369 173848 206374 173904
rect 206430 173848 207060 173904
rect 206369 173846 207060 173848
rect 206369 173843 206435 173846
rect 207054 173844 207060 173846
rect 207124 173844 207130 173908
rect 224861 173226 224927 173229
rect 239254 173226 239260 173228
rect 224861 173224 239260 173226
rect 224861 173168 224866 173224
rect 224922 173168 239260 173224
rect 224861 173166 239260 173168
rect 224861 173163 224927 173166
rect 239254 173164 239260 173166
rect 239324 173164 239330 173228
rect 222193 172410 222259 172413
rect 222929 172410 222995 172413
rect 222193 172408 222995 172410
rect 222193 172352 222198 172408
rect 222254 172352 222934 172408
rect 222990 172352 222995 172408
rect 222193 172350 222995 172352
rect 222193 172347 222259 172350
rect 222929 172347 222995 172350
rect 205449 171730 205515 171733
rect 241646 171730 241652 171732
rect 205449 171728 241652 171730
rect 205449 171672 205454 171728
rect 205510 171672 241652 171728
rect 205449 171670 241652 171672
rect 205449 171667 205515 171670
rect 241646 171668 241652 171670
rect 241716 171668 241722 171732
rect 92473 171186 92539 171189
rect 222193 171186 222259 171189
rect 92473 171184 222259 171186
rect 92473 171128 92478 171184
rect 92534 171128 222198 171184
rect 222254 171128 222259 171184
rect 92473 171126 222259 171128
rect 92473 171123 92539 171126
rect 222193 171123 222259 171126
rect 61837 169826 61903 169829
rect 205633 169826 205699 169829
rect 61837 169824 205699 169826
rect 61837 169768 61842 169824
rect 61898 169768 205638 169824
rect 205694 169768 205699 169824
rect 61837 169766 205699 169768
rect 61837 169763 61903 169766
rect 205633 169763 205699 169766
rect 82077 168466 82143 168469
rect 201493 168466 201559 168469
rect 202137 168466 202203 168469
rect 82077 168464 202203 168466
rect 82077 168408 82082 168464
rect 82138 168408 201498 168464
rect 201554 168408 202142 168464
rect 202198 168408 202203 168464
rect 82077 168406 202203 168408
rect 82077 168403 82143 168406
rect 201493 168403 201559 168406
rect 202137 168403 202203 168406
rect 117957 167242 118023 167245
rect 223573 167242 223639 167245
rect 224217 167242 224283 167245
rect 117957 167240 224283 167242
rect 117957 167184 117962 167240
rect 118018 167184 223578 167240
rect 223634 167184 224222 167240
rect 224278 167184 224283 167240
rect 117957 167182 224283 167184
rect 117957 167179 118023 167182
rect 223573 167179 223639 167182
rect 224217 167179 224283 167182
rect 86953 167106 87019 167109
rect 215477 167106 215543 167109
rect 216029 167106 216095 167109
rect 86953 167104 216095 167106
rect 86953 167048 86958 167104
rect 87014 167048 215482 167104
rect 215538 167048 216034 167104
rect 216090 167048 216095 167104
rect 86953 167046 216095 167048
rect 86953 167043 87019 167046
rect 215477 167043 215543 167046
rect 216029 167043 216095 167046
rect 97257 166290 97323 166293
rect 97809 166290 97875 166293
rect 252553 166292 252619 166293
rect 252502 166290 252508 166292
rect 97257 166288 252508 166290
rect 252572 166290 252619 166292
rect 252572 166288 252700 166290
rect 97257 166232 97262 166288
rect 97318 166232 97814 166288
rect 97870 166232 252508 166288
rect 252614 166232 252700 166288
rect 97257 166230 252508 166232
rect 97257 166227 97323 166230
rect 97809 166227 97875 166230
rect 252502 166228 252508 166230
rect 252572 166230 252700 166232
rect 252572 166228 252619 166230
rect 252553 166227 252619 166228
rect 582741 165882 582807 165885
rect 583520 165882 584960 165972
rect 582741 165880 584960 165882
rect 582741 165824 582746 165880
rect 582802 165824 584960 165880
rect 582741 165822 584960 165824
rect 582741 165819 582807 165822
rect 151169 165746 151235 165749
rect 238753 165746 238819 165749
rect 151169 165744 238819 165746
rect 151169 165688 151174 165744
rect 151230 165688 238758 165744
rect 238814 165688 238819 165744
rect 583520 165732 584960 165822
rect 151169 165686 238819 165688
rect 151169 165683 151235 165686
rect 238753 165683 238819 165686
rect 196617 164930 196683 164933
rect 190410 164928 196683 164930
rect 190410 164872 196622 164928
rect 196678 164872 196683 164928
rect 190410 164870 196683 164872
rect 69606 164324 69612 164388
rect 69676 164386 69682 164388
rect 187550 164386 187556 164388
rect 69676 164326 187556 164386
rect 69676 164324 69682 164326
rect 187550 164324 187556 164326
rect 187620 164386 187626 164388
rect 190410 164386 190470 164870
rect 196617 164867 196683 164870
rect 187620 164326 190470 164386
rect 187620 164324 187626 164326
rect 227662 164188 227668 164252
rect 227732 164250 227738 164252
rect 227805 164250 227871 164253
rect 227732 164248 227871 164250
rect 227732 164192 227810 164248
rect 227866 164192 227871 164248
rect 227732 164190 227871 164192
rect 227732 164188 227738 164190
rect 227805 164187 227871 164190
rect -960 162890 480 162980
rect 3509 162890 3575 162893
rect -960 162888 3575 162890
rect -960 162832 3514 162888
rect 3570 162832 3575 162888
rect -960 162830 3575 162832
rect -960 162740 480 162830
rect 3509 162827 3575 162830
rect 102777 162890 102843 162893
rect 227662 162890 227668 162892
rect 102777 162888 227668 162890
rect 102777 162832 102782 162888
rect 102838 162832 227668 162888
rect 102777 162830 227668 162832
rect 102777 162827 102843 162830
rect 227662 162828 227668 162830
rect 227732 162828 227738 162892
rect 222285 162754 222351 162757
rect 222837 162754 222903 162757
rect 222285 162752 222903 162754
rect 222285 162696 222290 162752
rect 222346 162696 222842 162752
rect 222898 162696 222903 162752
rect 222285 162694 222903 162696
rect 222285 162691 222351 162694
rect 222837 162691 222903 162694
rect 229185 162754 229251 162757
rect 229737 162754 229803 162757
rect 229185 162752 229803 162754
rect 229185 162696 229190 162752
rect 229246 162696 229742 162752
rect 229798 162696 229803 162752
rect 229185 162694 229803 162696
rect 229185 162691 229251 162694
rect 229737 162691 229803 162694
rect 153837 161802 153903 161805
rect 153837 161800 229110 161802
rect 153837 161744 153842 161800
rect 153898 161744 229110 161800
rect 153837 161742 229110 161744
rect 153837 161739 153903 161742
rect 72417 161666 72483 161669
rect 184473 161666 184539 161669
rect 72417 161664 184539 161666
rect 72417 161608 72422 161664
rect 72478 161608 184478 161664
rect 184534 161608 184539 161664
rect 72417 161606 184539 161608
rect 72417 161603 72483 161606
rect 184473 161603 184539 161606
rect 92657 161530 92723 161533
rect 222285 161530 222351 161533
rect 92657 161528 222351 161530
rect 92657 161472 92662 161528
rect 92718 161472 222290 161528
rect 222346 161472 222351 161528
rect 92657 161470 222351 161472
rect 229050 161530 229110 161742
rect 229185 161530 229251 161533
rect 229050 161528 229251 161530
rect 229050 161472 229190 161528
rect 229246 161472 229251 161528
rect 229050 161470 229251 161472
rect 92657 161467 92723 161470
rect 222285 161467 222351 161470
rect 229185 161467 229251 161470
rect 60549 160850 60615 160853
rect 193397 160850 193463 160853
rect 60549 160848 193463 160850
rect 60549 160792 60554 160848
rect 60610 160792 193402 160848
rect 193458 160792 193463 160848
rect 60549 160790 193463 160792
rect 60549 160787 60615 160790
rect 193397 160787 193463 160790
rect 188981 160714 189047 160717
rect 212390 160714 212396 160716
rect 188981 160712 212396 160714
rect 188981 160656 188986 160712
rect 189042 160656 212396 160712
rect 188981 160654 212396 160656
rect 188981 160651 189047 160654
rect 212390 160652 212396 160654
rect 212460 160714 212466 160716
rect 340137 160714 340203 160717
rect 212460 160712 340203 160714
rect 212460 160656 340142 160712
rect 340198 160656 340203 160712
rect 212460 160654 340203 160656
rect 212460 160652 212466 160654
rect 340137 160651 340203 160654
rect 145649 160170 145715 160173
rect 231945 160170 232011 160173
rect 232589 160170 232655 160173
rect 145649 160168 232655 160170
rect 145649 160112 145654 160168
rect 145710 160112 231950 160168
rect 232006 160112 232594 160168
rect 232650 160112 232655 160168
rect 145649 160110 232655 160112
rect 145649 160107 145715 160110
rect 231945 160107 232011 160110
rect 232589 160107 232655 160110
rect 73337 159354 73403 159357
rect 103421 159354 103487 159357
rect 188429 159354 188495 159357
rect 73337 159352 188495 159354
rect 73337 159296 73342 159352
rect 73398 159296 103426 159352
rect 103482 159296 188434 159352
rect 188490 159296 188495 159352
rect 73337 159294 188495 159296
rect 73337 159291 73403 159294
rect 103421 159291 103487 159294
rect 188429 159291 188495 159294
rect 196065 159354 196131 159357
rect 196893 159354 196959 159357
rect 231853 159354 231919 159357
rect 196065 159352 231919 159354
rect 196065 159296 196070 159352
rect 196126 159296 196898 159352
rect 196954 159296 231858 159352
rect 231914 159296 231919 159352
rect 196065 159294 231919 159296
rect 196065 159291 196131 159294
rect 196893 159291 196959 159294
rect 231853 159291 231919 159294
rect 173249 158810 173315 158813
rect 266445 158810 266511 158813
rect 173249 158808 266511 158810
rect 173249 158752 173254 158808
rect 173310 158752 266450 158808
rect 266506 158752 266511 158808
rect 173249 158750 266511 158752
rect 173249 158747 173315 158750
rect 266445 158747 266511 158750
rect 54937 157450 55003 157453
rect 142981 157450 143047 157453
rect 54937 157448 143047 157450
rect 54937 157392 54942 157448
rect 54998 157392 142986 157448
rect 143042 157392 143047 157448
rect 54937 157390 143047 157392
rect 54937 157387 55003 157390
rect 142981 157387 143047 157390
rect 154205 157450 154271 157453
rect 216673 157450 216739 157453
rect 217409 157450 217475 157453
rect 154205 157448 217475 157450
rect 154205 157392 154210 157448
rect 154266 157392 216678 157448
rect 216734 157392 217414 157448
rect 217470 157392 217475 157448
rect 154205 157390 217475 157392
rect 154205 157387 154271 157390
rect 216673 157387 216739 157390
rect 217409 157387 217475 157390
rect 86769 156634 86835 156637
rect 89846 156634 89852 156636
rect 86769 156632 89852 156634
rect 86769 156576 86774 156632
rect 86830 156576 89852 156632
rect 86769 156574 89852 156576
rect 86769 156571 86835 156574
rect 89846 156572 89852 156574
rect 89916 156572 89922 156636
rect 103421 156634 103487 156637
rect 189717 156634 189783 156637
rect 103421 156632 189783 156634
rect 103421 156576 103426 156632
rect 103482 156576 189722 156632
rect 189778 156576 189783 156632
rect 103421 156574 189783 156576
rect 103421 156571 103487 156574
rect 189717 156571 189783 156574
rect 205081 156226 205147 156229
rect 205541 156226 205607 156229
rect 222929 156226 222995 156229
rect 205081 156224 222995 156226
rect 205081 156168 205086 156224
rect 205142 156168 205546 156224
rect 205602 156168 222934 156224
rect 222990 156168 222995 156224
rect 205081 156166 222995 156168
rect 205081 156163 205147 156166
rect 205541 156163 205607 156166
rect 222929 156163 222995 156166
rect 187049 156090 187115 156093
rect 231853 156090 231919 156093
rect 232497 156090 232563 156093
rect 187049 156088 232563 156090
rect 187049 156032 187054 156088
rect 187110 156032 231858 156088
rect 231914 156032 232502 156088
rect 232558 156032 232563 156088
rect 187049 156030 232563 156032
rect 187049 156027 187115 156030
rect 231853 156027 231919 156030
rect 232497 156027 232563 156030
rect 60641 155274 60707 155277
rect 213678 155274 213684 155276
rect 60641 155272 213684 155274
rect 60641 155216 60646 155272
rect 60702 155216 213684 155272
rect 60641 155214 213684 155216
rect 60641 155211 60707 155214
rect 213678 155212 213684 155214
rect 213748 155212 213754 155276
rect 198089 154730 198155 154733
rect 198641 154730 198707 154733
rect 226374 154730 226380 154732
rect 198089 154728 226380 154730
rect 198089 154672 198094 154728
rect 198150 154672 198646 154728
rect 198702 154672 226380 154728
rect 198089 154670 226380 154672
rect 198089 154667 198155 154670
rect 198641 154667 198707 154670
rect 226374 154668 226380 154670
rect 226444 154668 226450 154732
rect 108481 154594 108547 154597
rect 228214 154594 228220 154596
rect 108481 154592 228220 154594
rect 108481 154536 108486 154592
rect 108542 154536 228220 154592
rect 108481 154534 228220 154536
rect 108481 154531 108547 154534
rect 228214 154532 228220 154534
rect 228284 154532 228290 154596
rect 77293 153778 77359 153781
rect 113173 153778 113239 153781
rect 188061 153778 188127 153781
rect 77293 153776 188127 153778
rect 77293 153720 77298 153776
rect 77354 153720 113178 153776
rect 113234 153720 188066 153776
rect 188122 153720 188127 153776
rect 77293 153718 188127 153720
rect 77293 153715 77359 153718
rect 113173 153715 113239 153718
rect 188061 153715 188127 153718
rect 116669 153234 116735 153237
rect 234613 153234 234679 153237
rect 116669 153232 234679 153234
rect 116669 153176 116674 153232
rect 116730 153176 234618 153232
rect 234674 153176 234679 153232
rect 116669 153174 234679 153176
rect 116669 153171 116735 153174
rect 234613 153171 234679 153174
rect 50705 153098 50771 153101
rect 50838 153098 50844 153100
rect 50705 153096 50844 153098
rect 50705 153040 50710 153096
rect 50766 153040 50844 153096
rect 50705 153038 50844 153040
rect 50705 153035 50771 153038
rect 50838 153036 50844 153038
rect 50908 153036 50914 153100
rect 582557 152690 582623 152693
rect 583520 152690 584960 152780
rect 582557 152688 584960 152690
rect 582557 152632 582562 152688
rect 582618 152632 584960 152688
rect 582557 152630 584960 152632
rect 582557 152627 582623 152630
rect 583520 152540 584960 152630
rect 148409 152418 148475 152421
rect 215937 152418 216003 152421
rect 229093 152418 229159 152421
rect 148409 152416 229159 152418
rect 148409 152360 148414 152416
rect 148470 152360 215942 152416
rect 215998 152360 229098 152416
rect 229154 152360 229159 152416
rect 148409 152358 229159 152360
rect 148409 152355 148475 152358
rect 215937 152355 216003 152358
rect 229093 152355 229159 152358
rect 50705 151874 50771 151877
rect 189717 151874 189783 151877
rect 50705 151872 189783 151874
rect 50705 151816 50710 151872
rect 50766 151816 189722 151872
rect 189778 151816 189783 151872
rect 50705 151814 189783 151816
rect 50705 151811 50771 151814
rect 189717 151811 189783 151814
rect 50797 150786 50863 150789
rect 188337 150786 188403 150789
rect 50797 150784 188403 150786
rect 50797 150728 50802 150784
rect 50858 150728 188342 150784
rect 188398 150728 188403 150784
rect 50797 150726 188403 150728
rect 50797 150723 50863 150726
rect 188337 150723 188403 150726
rect 229277 150650 229343 150653
rect 122790 150648 229343 150650
rect 122790 150592 229282 150648
rect 229338 150592 229343 150648
rect 122790 150590 229343 150592
rect 115197 150514 115263 150517
rect 115749 150514 115815 150517
rect 122790 150514 122850 150590
rect 229277 150587 229343 150590
rect 115197 150512 122850 150514
rect 115197 150456 115202 150512
rect 115258 150456 115754 150512
rect 115810 150456 122850 150512
rect 115197 150454 122850 150456
rect 187141 150514 187207 150517
rect 259453 150514 259519 150517
rect 187141 150512 259519 150514
rect 187141 150456 187146 150512
rect 187202 150456 259458 150512
rect 259514 150456 259519 150512
rect 187141 150454 259519 150456
rect 115197 150451 115263 150454
rect 115749 150451 115815 150454
rect 187141 150451 187207 150454
rect 259453 150451 259519 150454
rect 208393 150378 208459 150381
rect 271873 150378 271939 150381
rect 208393 150376 271939 150378
rect 208393 150320 208398 150376
rect 208454 150320 271878 150376
rect 271934 150320 271939 150376
rect 208393 150318 271939 150320
rect 208393 150315 208459 150318
rect 271873 150315 271939 150318
rect -960 149834 480 149924
rect 3141 149834 3207 149837
rect -960 149832 3207 149834
rect -960 149776 3146 149832
rect 3202 149776 3207 149832
rect -960 149774 3207 149776
rect -960 149684 480 149774
rect 3141 149771 3207 149774
rect 53649 149698 53715 149701
rect 169109 149698 169175 149701
rect 53649 149696 169175 149698
rect 53649 149640 53654 149696
rect 53710 149640 169114 149696
rect 169170 149640 169175 149696
rect 53649 149638 169175 149640
rect 53649 149635 53715 149638
rect 169109 149635 169175 149638
rect 184197 149698 184263 149701
rect 198089 149698 198155 149701
rect 184197 149696 198155 149698
rect 184197 149640 184202 149696
rect 184258 149640 198094 149696
rect 198150 149640 198155 149696
rect 184197 149638 198155 149640
rect 184197 149635 184263 149638
rect 198089 149635 198155 149638
rect 53557 149154 53623 149157
rect 127709 149154 127775 149157
rect 53557 149152 127775 149154
rect 53557 149096 53562 149152
rect 53618 149096 127714 149152
rect 127770 149096 127775 149152
rect 53557 149094 127775 149096
rect 53557 149091 53623 149094
rect 127709 149091 127775 149094
rect 169293 149154 169359 149157
rect 233233 149154 233299 149157
rect 169293 149152 233299 149154
rect 169293 149096 169298 149152
rect 169354 149096 233238 149152
rect 233294 149096 233299 149152
rect 169293 149094 233299 149096
rect 169293 149091 169359 149094
rect 233233 149091 233299 149094
rect 189901 148610 189967 148613
rect 197905 148610 197971 148613
rect 189901 148608 197971 148610
rect 189901 148552 189906 148608
rect 189962 148552 197910 148608
rect 197966 148552 197971 148608
rect 189901 148550 197971 148552
rect 189901 148547 189967 148550
rect 197905 148547 197971 148550
rect 191557 148474 191623 148477
rect 210233 148474 210299 148477
rect 191557 148472 210299 148474
rect 191557 148416 191562 148472
rect 191618 148416 210238 148472
rect 210294 148416 210299 148472
rect 191557 148414 210299 148416
rect 191557 148411 191623 148414
rect 210233 148411 210299 148414
rect 213678 148412 213684 148476
rect 213748 148474 213754 148476
rect 222377 148474 222443 148477
rect 213748 148472 222443 148474
rect 213748 148416 222382 148472
rect 222438 148416 222443 148472
rect 213748 148414 222443 148416
rect 213748 148412 213754 148414
rect 222377 148411 222443 148414
rect 50889 148338 50955 148341
rect 186957 148338 187023 148341
rect 50889 148336 187023 148338
rect 50889 148280 50894 148336
rect 50950 148280 186962 148336
rect 187018 148280 187023 148336
rect 50889 148278 187023 148280
rect 50889 148275 50955 148278
rect 186957 148275 187023 148278
rect 191649 148338 191715 148341
rect 242934 148338 242940 148340
rect 191649 148336 242940 148338
rect 191649 148280 191654 148336
rect 191710 148280 242940 148336
rect 191649 148278 242940 148280
rect 191649 148275 191715 148278
rect 242934 148276 242940 148278
rect 243004 148338 243010 148340
rect 268377 148338 268443 148341
rect 243004 148336 268443 148338
rect 243004 148280 268382 148336
rect 268438 148280 268443 148336
rect 243004 148278 268443 148280
rect 243004 148276 243010 148278
rect 268377 148275 268443 148278
rect 66662 147868 66668 147932
rect 66732 147930 66738 147932
rect 67541 147930 67607 147933
rect 66732 147928 67607 147930
rect 66732 147872 67546 147928
rect 67602 147872 67607 147928
rect 66732 147870 67607 147872
rect 66732 147868 66738 147870
rect 67541 147867 67607 147870
rect 65977 147794 66043 147797
rect 178677 147794 178743 147797
rect 65977 147792 178743 147794
rect 65977 147736 65982 147792
rect 66038 147736 178682 147792
rect 178738 147736 178743 147792
rect 65977 147734 178743 147736
rect 65977 147731 66043 147734
rect 178677 147731 178743 147734
rect 184289 147250 184355 147253
rect 196709 147250 196775 147253
rect 184289 147248 196775 147250
rect 184289 147192 184294 147248
rect 184350 147192 196714 147248
rect 196770 147192 196775 147248
rect 184289 147190 196775 147192
rect 184289 147187 184355 147190
rect 196709 147187 196775 147190
rect 96521 147114 96587 147117
rect 175825 147114 175891 147117
rect 96521 147112 175891 147114
rect 96521 147056 96526 147112
rect 96582 147056 175830 147112
rect 175886 147056 175891 147112
rect 96521 147054 175891 147056
rect 96521 147051 96587 147054
rect 175825 147051 175891 147054
rect 192702 147052 192708 147116
rect 192772 147114 192778 147116
rect 244406 147114 244412 147116
rect 192772 147054 244412 147114
rect 192772 147052 192778 147054
rect 244406 147052 244412 147054
rect 244476 147052 244482 147116
rect 81985 146978 82051 146981
rect 116577 146978 116643 146981
rect 210049 146978 210115 146981
rect 81985 146976 210115 146978
rect 81985 146920 81990 146976
rect 82046 146920 116582 146976
rect 116638 146920 210054 146976
rect 210110 146920 210115 146976
rect 81985 146918 210115 146920
rect 81985 146915 82051 146918
rect 116577 146915 116643 146918
rect 210049 146915 210115 146918
rect 188061 145890 188127 145893
rect 204437 145890 204503 145893
rect 188061 145888 204503 145890
rect 188061 145832 188066 145888
rect 188122 145832 204442 145888
rect 204498 145832 204503 145888
rect 188061 145830 204503 145832
rect 188061 145827 188127 145830
rect 204437 145827 204503 145830
rect 184473 145754 184539 145757
rect 196525 145754 196591 145757
rect 184473 145752 196591 145754
rect 184473 145696 184478 145752
rect 184534 145696 196530 145752
rect 196586 145696 196591 145752
rect 184473 145694 196591 145696
rect 184473 145691 184539 145694
rect 196525 145691 196591 145694
rect 201401 145754 201467 145757
rect 219382 145754 219388 145756
rect 201401 145752 219388 145754
rect 201401 145696 201406 145752
rect 201462 145696 219388 145752
rect 201401 145694 219388 145696
rect 201401 145691 201467 145694
rect 219382 145692 219388 145694
rect 219452 145692 219458 145756
rect 85481 145618 85547 145621
rect 100702 145618 100708 145620
rect 85481 145616 100708 145618
rect 85481 145560 85486 145616
rect 85542 145560 100708 145616
rect 85481 145558 100708 145560
rect 85481 145555 85547 145558
rect 100702 145556 100708 145558
rect 100772 145556 100778 145620
rect 178769 145618 178835 145621
rect 188889 145618 188955 145621
rect 282913 145618 282979 145621
rect 178769 145616 282979 145618
rect 178769 145560 178774 145616
rect 178830 145560 188894 145616
rect 188950 145560 282918 145616
rect 282974 145560 282979 145616
rect 178769 145558 282979 145560
rect 178769 145555 178835 145558
rect 188889 145555 188955 145558
rect 282913 145555 282979 145558
rect 63125 144938 63191 144941
rect 161565 144938 161631 144941
rect 162117 144938 162183 144941
rect 63125 144936 162183 144938
rect 63125 144880 63130 144936
rect 63186 144880 161570 144936
rect 161626 144880 162122 144936
rect 162178 144880 162183 144936
rect 63125 144878 162183 144880
rect 63125 144875 63191 144878
rect 161565 144875 161631 144878
rect 162117 144875 162183 144878
rect 65742 144740 65748 144804
rect 65812 144802 65818 144804
rect 65885 144802 65951 144805
rect 65812 144800 65951 144802
rect 65812 144744 65890 144800
rect 65946 144744 65951 144800
rect 65812 144742 65951 144744
rect 65812 144740 65818 144742
rect 65885 144739 65951 144742
rect 182173 144802 182239 144805
rect 183461 144802 183527 144805
rect 182173 144800 183527 144802
rect 182173 144744 182178 144800
rect 182234 144744 183466 144800
rect 183522 144744 183527 144800
rect 182173 144742 183527 144744
rect 182173 144739 182239 144742
rect 183461 144739 183527 144742
rect 188429 144258 188495 144261
rect 200205 144258 200271 144261
rect 188429 144256 200271 144258
rect 188429 144200 188434 144256
rect 188490 144200 200210 144256
rect 200266 144200 200271 144256
rect 188429 144198 200271 144200
rect 188429 144195 188495 144198
rect 200205 144195 200271 144198
rect 93025 144122 93091 144125
rect 117957 144122 118023 144125
rect 93025 144120 118023 144122
rect 93025 144064 93030 144120
rect 93086 144064 117962 144120
rect 118018 144064 118023 144120
rect 93025 144062 118023 144064
rect 93025 144059 93091 144062
rect 117957 144059 118023 144062
rect 118601 144122 118667 144125
rect 184054 144122 184060 144124
rect 118601 144120 184060 144122
rect 118601 144064 118606 144120
rect 118662 144064 184060 144120
rect 118601 144062 184060 144064
rect 118601 144059 118667 144062
rect 184054 144060 184060 144062
rect 184124 144060 184130 144124
rect 193121 144122 193187 144125
rect 205633 144122 205699 144125
rect 193121 144120 205699 144122
rect 193121 144064 193126 144120
rect 193182 144064 205638 144120
rect 205694 144064 205699 144120
rect 193121 144062 205699 144064
rect 193121 144059 193187 144062
rect 205633 144059 205699 144062
rect 94957 143986 95023 143989
rect 84150 143984 95023 143986
rect 84150 143928 94962 143984
rect 95018 143928 95023 143984
rect 84150 143926 95023 143928
rect 65885 143714 65951 143717
rect 84150 143714 84210 143926
rect 94957 143923 95023 143926
rect 65885 143712 84210 143714
rect 65885 143656 65890 143712
rect 65946 143656 84210 143712
rect 65885 143654 84210 143656
rect 84561 143714 84627 143717
rect 88742 143714 88748 143716
rect 84561 143712 88748 143714
rect 84561 143656 84566 143712
rect 84622 143656 88748 143712
rect 84561 143654 88748 143656
rect 65885 143651 65951 143654
rect 84561 143651 84627 143654
rect 88742 143652 88748 143654
rect 88812 143714 88818 143716
rect 89161 143714 89227 143717
rect 198825 143716 198891 143717
rect 88812 143712 89227 143714
rect 88812 143656 89166 143712
rect 89222 143656 89227 143712
rect 88812 143654 89227 143656
rect 88812 143652 88818 143654
rect 89161 143651 89227 143654
rect 198774 143652 198780 143716
rect 198844 143714 198891 143716
rect 198844 143712 198936 143714
rect 198886 143656 198936 143712
rect 198844 143654 198936 143656
rect 198844 143652 198891 143654
rect 198825 143651 198891 143652
rect 59077 143578 59143 143581
rect 160737 143578 160803 143581
rect 59077 143576 160803 143578
rect 59077 143520 59082 143576
rect 59138 143520 160742 143576
rect 160798 143520 160803 143576
rect 59077 143518 160803 143520
rect 59077 143515 59143 143518
rect 160737 143515 160803 143518
rect 183461 143578 183527 143581
rect 201309 143578 201375 143581
rect 183461 143576 201375 143578
rect 183461 143520 183466 143576
rect 183522 143520 201314 143576
rect 201370 143520 201375 143576
rect 183461 143518 201375 143520
rect 183461 143515 183527 143518
rect 201309 143515 201375 143518
rect 204897 143578 204963 143581
rect 205541 143578 205607 143581
rect 249149 143578 249215 143581
rect 204897 143576 249215 143578
rect 204897 143520 204902 143576
rect 204958 143520 205546 143576
rect 205602 143520 249154 143576
rect 249210 143520 249215 143576
rect 204897 143518 249215 143520
rect 204897 143515 204963 143518
rect 205541 143515 205607 143518
rect 249149 143515 249215 143518
rect 194685 143442 194751 143445
rect 195237 143442 195303 143445
rect 194685 143440 195303 143442
rect 194685 143384 194690 143440
rect 194746 143384 195242 143440
rect 195298 143384 195303 143440
rect 194685 143382 195303 143384
rect 194685 143379 194751 143382
rect 195237 143379 195303 143382
rect 197997 143442 198063 143445
rect 198917 143442 198983 143445
rect 197997 143440 198983 143442
rect 197997 143384 198002 143440
rect 198058 143384 198922 143440
rect 198978 143384 198983 143440
rect 197997 143382 198983 143384
rect 197997 143379 198063 143382
rect 198917 143379 198983 143382
rect 89161 142762 89227 142765
rect 213453 142762 213519 142765
rect 89161 142760 213519 142762
rect 89161 142704 89166 142760
rect 89222 142704 213458 142760
rect 213514 142704 213519 142760
rect 89161 142702 213519 142704
rect 89161 142699 89227 142702
rect 213453 142699 213519 142702
rect 219525 142762 219591 142765
rect 220997 142762 221063 142765
rect 582833 142762 582899 142765
rect 219525 142760 582899 142762
rect 219525 142704 219530 142760
rect 219586 142704 221002 142760
rect 221058 142704 582838 142760
rect 582894 142704 582899 142760
rect 219525 142702 582899 142704
rect 219525 142699 219591 142702
rect 220997 142699 221063 142702
rect 582833 142699 582899 142702
rect 189073 142354 189139 142357
rect 196566 142354 196572 142356
rect 189073 142352 196572 142354
rect 189073 142296 189078 142352
rect 189134 142296 196572 142352
rect 189073 142294 196572 142296
rect 189073 142291 189139 142294
rect 196566 142292 196572 142294
rect 196636 142354 196642 142356
rect 197077 142354 197143 142357
rect 196636 142352 197143 142354
rect 196636 142296 197082 142352
rect 197138 142296 197143 142352
rect 196636 142294 197143 142296
rect 196636 142292 196642 142294
rect 197077 142291 197143 142294
rect 63309 142218 63375 142221
rect 90950 142218 90956 142220
rect 63309 142216 90956 142218
rect 63309 142160 63314 142216
rect 63370 142160 90956 142216
rect 63309 142158 90956 142160
rect 63309 142155 63375 142158
rect 90950 142156 90956 142158
rect 91020 142156 91026 142220
rect 105077 142218 105143 142221
rect 194685 142218 194751 142221
rect 105077 142216 194751 142218
rect 105077 142160 105082 142216
rect 105138 142160 194690 142216
rect 194746 142160 194751 142216
rect 105077 142158 194751 142160
rect 105077 142155 105143 142158
rect 194685 142155 194751 142158
rect 195973 142218 196039 142221
rect 196893 142218 196959 142221
rect 197118 142218 197124 142220
rect 195973 142216 197124 142218
rect 195973 142160 195978 142216
rect 196034 142160 196898 142216
rect 196954 142160 197124 142216
rect 195973 142158 197124 142160
rect 195973 142155 196039 142158
rect 196893 142155 196959 142158
rect 197118 142156 197124 142158
rect 197188 142156 197194 142220
rect 200614 142156 200620 142220
rect 200684 142218 200690 142220
rect 201401 142218 201467 142221
rect 200684 142216 201467 142218
rect 200684 142160 201406 142216
rect 201462 142160 201467 142216
rect 200684 142158 201467 142160
rect 200684 142156 200690 142158
rect 201401 142155 201467 142158
rect 213453 142218 213519 142221
rect 257337 142218 257403 142221
rect 213453 142216 257403 142218
rect 213453 142160 213458 142216
rect 213514 142160 257342 142216
rect 257398 142160 257403 142216
rect 213453 142158 257403 142160
rect 213453 142155 213519 142158
rect 257337 142155 257403 142158
rect 222929 142082 222995 142085
rect 224350 142082 224356 142084
rect 222929 142080 224356 142082
rect 222929 142024 222934 142080
rect 222990 142024 224356 142080
rect 222929 142022 224356 142024
rect 222929 142019 222995 142022
rect 224350 142020 224356 142022
rect 224420 142020 224426 142084
rect 74257 141538 74323 141541
rect 173801 141538 173867 141541
rect 74257 141536 173867 141538
rect 74257 141480 74262 141536
rect 74318 141480 173806 141536
rect 173862 141480 173867 141536
rect 74257 141478 173867 141480
rect 74257 141475 74323 141478
rect 173801 141475 173867 141478
rect 70301 141404 70367 141405
rect 70301 141402 70348 141404
rect 70256 141400 70348 141402
rect 70256 141344 70306 141400
rect 70256 141342 70348 141344
rect 70301 141340 70348 141342
rect 70412 141340 70418 141404
rect 81341 141402 81407 141405
rect 204989 141402 205055 141405
rect 205449 141402 205515 141405
rect 81341 141400 205515 141402
rect 81341 141344 81346 141400
rect 81402 141344 204994 141400
rect 205050 141344 205454 141400
rect 205510 141344 205515 141400
rect 81341 141342 205515 141344
rect 70301 141339 70367 141340
rect 81341 141339 81407 141342
rect 204989 141339 205055 141342
rect 205449 141339 205515 141342
rect 218789 141402 218855 141405
rect 225321 141402 225387 141405
rect 218789 141400 225387 141402
rect 218789 141344 218794 141400
rect 218850 141344 225326 141400
rect 225382 141344 225387 141400
rect 218789 141342 225387 141344
rect 218789 141339 218855 141342
rect 225321 141339 225387 141342
rect 198641 141130 198707 141133
rect 198774 141130 198780 141132
rect 198641 141128 198780 141130
rect 198641 141072 198646 141128
rect 198702 141072 198780 141128
rect 198641 141070 198780 141072
rect 198641 141067 198707 141070
rect 198774 141068 198780 141070
rect 198844 141130 198850 141132
rect 214741 141130 214807 141133
rect 198844 141128 214807 141130
rect 198844 141072 214746 141128
rect 214802 141072 214807 141128
rect 198844 141070 214807 141072
rect 198844 141068 198850 141070
rect 214741 141067 214807 141070
rect 205081 140994 205147 140997
rect 238017 140994 238083 140997
rect 205081 140992 238083 140994
rect 205081 140936 205086 140992
rect 205142 140936 238022 140992
rect 238078 140936 238083 140992
rect 205081 140934 238083 140936
rect 205081 140931 205147 140934
rect 238017 140931 238083 140934
rect 73061 140860 73127 140861
rect 73061 140856 73108 140860
rect 73172 140858 73178 140860
rect 89621 140858 89687 140861
rect 218881 140858 218947 140861
rect 73061 140800 73066 140856
rect 73061 140796 73108 140800
rect 73172 140798 73218 140858
rect 89621 140856 218947 140858
rect 89621 140800 89626 140856
rect 89682 140800 218886 140856
rect 218942 140800 218947 140856
rect 89621 140798 218947 140800
rect 73172 140796 73178 140798
rect 73061 140795 73127 140796
rect 89621 140795 89687 140798
rect 218881 140795 218947 140798
rect 203517 140450 203583 140453
rect 195930 140448 203583 140450
rect 195930 140392 203522 140448
rect 203578 140392 203583 140448
rect 195930 140390 203583 140392
rect 76649 140178 76715 140181
rect 195930 140178 195990 140390
rect 203517 140387 203583 140390
rect 76649 140176 195990 140178
rect 76649 140120 76654 140176
rect 76710 140120 195990 140176
rect 76649 140118 195990 140120
rect 76649 140115 76715 140118
rect 231945 140042 232011 140045
rect 229050 140040 232011 140042
rect 229050 139984 231950 140040
rect 232006 139984 232011 140040
rect 229050 139982 232011 139984
rect 229050 139906 229110 139982
rect 231945 139979 232011 139982
rect 84469 139634 84535 139637
rect 87597 139634 87663 139637
rect 84469 139632 87663 139634
rect 84469 139576 84474 139632
rect 84530 139576 87602 139632
rect 87658 139576 87663 139632
rect 84469 139574 87663 139576
rect 84469 139571 84535 139574
rect 87597 139571 87663 139574
rect 193254 139572 193260 139636
rect 193324 139634 193330 139636
rect 193397 139634 193463 139637
rect 193324 139632 193463 139634
rect 193324 139576 193402 139632
rect 193458 139576 193463 139632
rect 193324 139574 193463 139576
rect 193324 139572 193330 139574
rect 193397 139571 193463 139574
rect 62021 139498 62087 139501
rect 102869 139498 102935 139501
rect 62021 139496 102935 139498
rect 62021 139440 62026 139496
rect 62082 139440 102874 139496
rect 102930 139440 102935 139496
rect 62021 139438 102935 139440
rect 62021 139435 62087 139438
rect 102869 139435 102935 139438
rect 187693 139498 187759 139501
rect 188981 139498 189047 139501
rect 193630 139498 193690 139876
rect 224940 139846 229110 139906
rect 187693 139496 193690 139498
rect 187693 139440 187698 139496
rect 187754 139440 188986 139496
rect 189042 139440 193690 139496
rect 187693 139438 193690 139440
rect 187693 139435 187759 139438
rect 188981 139435 189047 139438
rect 580349 139362 580415 139365
rect 583520 139362 584960 139452
rect 580349 139360 584960 139362
rect 580349 139304 580354 139360
rect 580410 139304 584960 139360
rect 580349 139302 584960 139304
rect 580349 139299 580415 139302
rect 583520 139212 584960 139302
rect 227662 139090 227668 139092
rect 64597 138818 64663 138821
rect 76557 138818 76623 138821
rect 64597 138816 76623 138818
rect 64597 138760 64602 138816
rect 64658 138760 76562 138816
rect 76618 138760 76623 138816
rect 64597 138758 76623 138760
rect 64597 138755 64663 138758
rect 76557 138755 76623 138758
rect 75821 138682 75887 138685
rect 167821 138682 167887 138685
rect 75821 138680 167887 138682
rect 75821 138624 75826 138680
rect 75882 138624 167826 138680
rect 167882 138624 167887 138680
rect 75821 138622 167887 138624
rect 75821 138619 75887 138622
rect 167821 138619 167887 138622
rect 189717 138546 189783 138549
rect 193630 138546 193690 139060
rect 224940 139030 227668 139090
rect 227662 139028 227668 139030
rect 227732 139028 227738 139092
rect 229185 138682 229251 138685
rect 582557 138682 582623 138685
rect 189717 138544 193690 138546
rect 189717 138488 189722 138544
rect 189778 138488 193690 138544
rect 189717 138486 193690 138488
rect 224910 138680 582623 138682
rect 224910 138624 229190 138680
rect 229246 138624 582562 138680
rect 582618 138624 582623 138680
rect 224910 138622 582623 138624
rect 189717 138483 189783 138486
rect 95141 138274 95207 138277
rect 95417 138274 95483 138277
rect 95141 138272 95483 138274
rect 95141 138216 95146 138272
rect 95202 138216 95422 138272
rect 95478 138216 95483 138272
rect 95141 138214 95483 138216
rect 95141 138211 95207 138214
rect 95417 138211 95483 138214
rect 191557 138274 191623 138277
rect 191557 138272 193660 138274
rect 191557 138216 191562 138272
rect 191618 138216 193660 138272
rect 224910 138244 224970 138622
rect 229185 138619 229251 138622
rect 582557 138619 582623 138622
rect 191557 138214 193660 138216
rect 191557 138211 191623 138214
rect 69422 138076 69428 138140
rect 69492 138138 69498 138140
rect 104157 138138 104223 138141
rect 69492 138136 104223 138138
rect 69492 138080 104162 138136
rect 104218 138080 104223 138136
rect 69492 138078 104223 138080
rect 69492 138076 69498 138078
rect 104157 138075 104223 138078
rect 69289 138002 69355 138005
rect 70342 138002 70348 138004
rect 69289 138000 70348 138002
rect 69289 137944 69294 138000
rect 69350 137944 70348 138000
rect 69289 137942 70348 137944
rect 69289 137939 69355 137942
rect 70342 137940 70348 137942
rect 70412 137940 70418 138004
rect 75545 138002 75611 138005
rect 82077 138002 82143 138005
rect 75545 138000 82143 138002
rect 75545 137944 75550 138000
rect 75606 137944 82082 138000
rect 82138 137944 82143 138000
rect 75545 137942 82143 137944
rect 75545 137939 75611 137942
rect 82077 137939 82143 137942
rect 72325 137866 72391 137869
rect 75177 137866 75243 137869
rect 72325 137864 75243 137866
rect 72325 137808 72330 137864
rect 72386 137808 75182 137864
rect 75238 137808 75243 137864
rect 72325 137806 75243 137808
rect 72325 137803 72391 137806
rect 75177 137803 75243 137806
rect 192845 137458 192911 137461
rect 192845 137456 193660 137458
rect 192845 137400 192850 137456
rect 192906 137400 193660 137456
rect 192845 137398 193660 137400
rect 192845 137395 192911 137398
rect 71681 137322 71747 137325
rect 86309 137322 86375 137325
rect 71681 137320 86375 137322
rect 71681 137264 71686 137320
rect 71742 137264 86314 137320
rect 86370 137264 86375 137320
rect 71681 137262 86375 137264
rect 71681 137259 71747 137262
rect 86309 137259 86375 137262
rect 70853 137186 70919 137189
rect 72417 137186 72483 137189
rect 226333 137186 226399 137189
rect 70853 137184 72483 137186
rect 70853 137128 70858 137184
rect 70914 137128 72422 137184
rect 72478 137128 72483 137184
rect 70853 137126 72483 137128
rect 224940 137184 226399 137186
rect 224940 137128 226338 137184
rect 226394 137128 226399 137184
rect 224940 137126 226399 137128
rect 70853 137123 70919 137126
rect 72417 137123 72483 137126
rect 226333 137123 226399 137126
rect -960 136778 480 136868
rect 68134 136852 68140 136916
rect 68204 136914 68210 136916
rect 94814 136914 94820 136916
rect 68204 136854 94820 136914
rect 68204 136852 68210 136854
rect 94814 136852 94820 136854
rect 94884 136852 94890 136916
rect 3509 136778 3575 136781
rect -960 136776 3575 136778
rect -960 136720 3514 136776
rect 3570 136720 3575 136776
rect -960 136718 3575 136720
rect -960 136628 480 136718
rect 3509 136715 3575 136718
rect 85481 136778 85547 136781
rect 88977 136778 89043 136781
rect 85481 136776 89043 136778
rect 85481 136720 85486 136776
rect 85542 136720 88982 136776
rect 89038 136720 89043 136776
rect 85481 136718 89043 136720
rect 85481 136715 85547 136718
rect 88977 136715 89043 136718
rect 224350 136580 224356 136644
rect 224420 136580 224426 136644
rect 226926 136580 226932 136644
rect 226996 136642 227002 136644
rect 227846 136642 227852 136644
rect 226996 136582 227852 136642
rect 226996 136580 227002 136582
rect 227846 136580 227852 136582
rect 227916 136580 227922 136644
rect 191557 136370 191623 136373
rect 191557 136368 193660 136370
rect 191557 136312 191562 136368
rect 191618 136312 193660 136368
rect 224358 136340 224418 136580
rect 191557 136310 193660 136312
rect 191557 136307 191623 136310
rect 54477 136098 54543 136101
rect 91093 136098 91159 136101
rect 91277 136098 91343 136101
rect 54477 136096 91343 136098
rect 54477 136040 54482 136096
rect 54538 136040 91098 136096
rect 91154 136040 91282 136096
rect 91338 136040 91343 136096
rect 54477 136038 91343 136040
rect 54477 136035 54543 136038
rect 91093 136035 91159 136038
rect 91277 136035 91343 136038
rect 74993 135962 75059 135965
rect 182173 135962 182239 135965
rect 74993 135960 182239 135962
rect 74993 135904 74998 135960
rect 75054 135904 182178 135960
rect 182234 135904 182239 135960
rect 74993 135902 182239 135904
rect 74993 135899 75059 135902
rect 182173 135899 182239 135902
rect 231945 135962 232011 135965
rect 341517 135962 341583 135965
rect 231945 135960 341583 135962
rect 231945 135904 231950 135960
rect 232006 135904 341522 135960
rect 341578 135904 341583 135960
rect 231945 135902 341583 135904
rect 231945 135899 232011 135902
rect 341517 135899 341583 135902
rect 191557 135554 191623 135557
rect 225321 135554 225387 135557
rect 191557 135552 193660 135554
rect 191557 135496 191562 135552
rect 191618 135496 193660 135552
rect 191557 135494 193660 135496
rect 224940 135552 225387 135554
rect 224940 135496 225326 135552
rect 225382 135496 225387 135552
rect 224940 135494 225387 135496
rect 191557 135491 191623 135494
rect 225321 135491 225387 135494
rect 90950 135220 90956 135284
rect 91020 135282 91026 135284
rect 95734 135282 95740 135284
rect 91020 135222 95740 135282
rect 91020 135220 91026 135222
rect 95734 135220 95740 135222
rect 95804 135220 95810 135284
rect 94129 135146 94195 135149
rect 187693 135146 187759 135149
rect 94129 135144 187759 135146
rect 94129 135088 94134 135144
rect 94190 135088 187698 135144
rect 187754 135088 187759 135144
rect 94129 135086 187759 135088
rect 94129 135083 94195 135086
rect 187693 135083 187759 135086
rect 69565 135010 69631 135013
rect 69430 135008 69631 135010
rect 69430 134952 69570 135008
rect 69626 134952 69631 135008
rect 69430 134950 69631 134952
rect 69430 134436 69490 134950
rect 69565 134947 69631 134950
rect 193029 134738 193095 134741
rect 226517 134738 226583 134741
rect 226701 134738 226767 134741
rect 193029 134736 193660 134738
rect 193029 134680 193034 134736
rect 193090 134680 193660 134736
rect 193029 134678 193660 134680
rect 224940 134736 226767 134738
rect 224940 134680 226522 134736
rect 226578 134680 226706 134736
rect 226762 134680 226767 134736
rect 224940 134678 226767 134680
rect 193029 134675 193095 134678
rect 226517 134675 226583 134678
rect 226701 134675 226767 134678
rect 96705 133922 96771 133925
rect 94668 133920 96771 133922
rect 94668 133864 96710 133920
rect 96766 133864 96771 133920
rect 94668 133862 96771 133864
rect 96705 133859 96771 133862
rect 189809 133922 189875 133925
rect 189809 133920 193660 133922
rect 189809 133864 189814 133920
rect 189870 133864 193660 133920
rect 189809 133862 193660 133864
rect 189809 133859 189875 133862
rect 94814 133724 94820 133788
rect 94884 133786 94890 133788
rect 190361 133786 190427 133789
rect 94884 133784 190427 133786
rect 94884 133728 190366 133784
rect 190422 133728 190427 133784
rect 94884 133726 190427 133728
rect 94884 133724 94890 133726
rect 190361 133723 190427 133726
rect 67725 133650 67791 133653
rect 226701 133650 226767 133653
rect 67725 133648 68908 133650
rect 67725 133592 67730 133648
rect 67786 133592 68908 133648
rect 67725 133590 68908 133592
rect 224940 133648 226767 133650
rect 224940 133592 226706 133648
rect 226762 133592 226767 133648
rect 224940 133590 226767 133592
rect 67725 133587 67791 133590
rect 226701 133587 226767 133590
rect 68829 133378 68895 133381
rect 68829 133376 68938 133378
rect 68829 133320 68834 133376
rect 68890 133320 68938 133376
rect 68829 133315 68938 133320
rect 68878 132804 68938 133315
rect 96705 133106 96771 133109
rect 94668 133104 96771 133106
rect 94668 133048 96710 133104
rect 96766 133048 96771 133104
rect 94668 133046 96771 133048
rect 96705 133043 96771 133046
rect 227069 132834 227135 132837
rect 224940 132832 227135 132834
rect 190361 132562 190427 132565
rect 193630 132562 193690 132804
rect 224940 132776 227074 132832
rect 227130 132776 227135 132832
rect 224940 132774 227135 132776
rect 227069 132771 227135 132774
rect 190361 132560 193690 132562
rect 190361 132504 190366 132560
rect 190422 132504 193690 132560
rect 190361 132502 193690 132504
rect 190361 132499 190427 132502
rect 66253 132018 66319 132021
rect 66253 132016 68908 132018
rect 66253 131960 66258 132016
rect 66314 131960 68908 132016
rect 66253 131958 68908 131960
rect 66253 131955 66319 131958
rect 94638 131746 94698 132260
rect 191649 132018 191715 132021
rect 226701 132018 226767 132021
rect 191649 132016 193660 132018
rect 191649 131960 191654 132016
rect 191710 131960 193660 132016
rect 191649 131958 193660 131960
rect 224940 132016 226767 132018
rect 224940 131960 226706 132016
rect 226762 131960 226767 132016
rect 224940 131958 226767 131960
rect 191649 131955 191715 131958
rect 226701 131955 226767 131958
rect 94638 131686 103530 131746
rect 96613 131474 96679 131477
rect 94668 131472 96679 131474
rect 94668 131416 96618 131472
rect 96674 131416 96679 131472
rect 94668 131414 96679 131416
rect 96613 131411 96679 131414
rect 66345 131202 66411 131205
rect 103470 131202 103530 131686
rect 153837 131202 153903 131205
rect 66345 131200 68908 131202
rect 66345 131144 66350 131200
rect 66406 131144 68908 131200
rect 66345 131142 68908 131144
rect 103470 131200 153903 131202
rect 103470 131144 153842 131200
rect 153898 131144 153903 131200
rect 103470 131142 153903 131144
rect 66345 131139 66411 131142
rect 153837 131139 153903 131142
rect 187550 131140 187556 131204
rect 187620 131202 187626 131204
rect 187620 131142 193660 131202
rect 187620 131140 187626 131142
rect 69422 131004 69428 131068
rect 69492 131004 69498 131068
rect 69430 130628 69490 131004
rect 97901 130930 97967 130933
rect 226701 130930 226767 130933
rect 94668 130928 97967 130930
rect 94668 130872 97906 130928
rect 97962 130872 97967 130928
rect 94668 130870 97967 130872
rect 224940 130928 226767 130930
rect 224940 130872 226706 130928
rect 226762 130872 226767 130928
rect 224940 130870 226767 130872
rect 97901 130867 97967 130870
rect 226701 130867 226767 130870
rect 96613 130114 96679 130117
rect 226374 130114 226380 130116
rect 94668 130112 96679 130114
rect 94668 130056 96618 130112
rect 96674 130056 96679 130112
rect 94668 130054 96679 130056
rect 96613 130051 96679 130054
rect 67265 129842 67331 129845
rect 190361 129842 190427 129845
rect 193630 129842 193690 130084
rect 224940 130054 226380 130114
rect 226374 130052 226380 130054
rect 226444 130052 226450 130116
rect 67265 129840 68908 129842
rect 67265 129784 67270 129840
rect 67326 129784 68908 129840
rect 67265 129782 68908 129784
rect 190361 129840 193690 129842
rect 190361 129784 190366 129840
rect 190422 129784 193690 129840
rect 190361 129782 193690 129784
rect 67265 129779 67331 129782
rect 190361 129779 190427 129782
rect 97533 129298 97599 129301
rect 191649 129300 191715 129301
rect 191598 129298 191604 129300
rect 94668 129296 97599 129298
rect 94668 129240 97538 129296
rect 97594 129240 97599 129296
rect 94668 129238 97599 129240
rect 191522 129238 191604 129298
rect 191668 129298 191715 129300
rect 226701 129298 226767 129301
rect 191668 129296 193660 129298
rect 191710 129240 193660 129296
rect 97533 129235 97599 129238
rect 191598 129236 191604 129238
rect 191668 129238 193660 129240
rect 224940 129296 226767 129298
rect 224940 129240 226706 129296
rect 226762 129240 226767 129296
rect 224940 129238 226767 129240
rect 191668 129236 191715 129238
rect 191649 129235 191715 129236
rect 226701 129235 226767 129238
rect 67725 129026 67791 129029
rect 67725 129024 68908 129026
rect 67725 128968 67730 129024
rect 67786 128968 68908 129024
rect 67725 128966 68908 128968
rect 67725 128963 67791 128966
rect 96705 128482 96771 128485
rect 94668 128480 96771 128482
rect 94668 128424 96710 128480
rect 96766 128424 96771 128480
rect 94668 128422 96771 128424
rect 96705 128419 96771 128422
rect 193121 128482 193187 128485
rect 226701 128482 226767 128485
rect 193121 128480 193660 128482
rect 193121 128424 193126 128480
rect 193182 128424 193660 128480
rect 193121 128422 193660 128424
rect 224940 128480 226767 128482
rect 224940 128424 226706 128480
rect 226762 128424 226767 128480
rect 224940 128422 226767 128424
rect 193121 128419 193187 128422
rect 226701 128419 226767 128422
rect 67817 128210 67883 128213
rect 67817 128208 68908 128210
rect 67817 128152 67822 128208
rect 67878 128152 68908 128208
rect 67817 128150 68908 128152
rect 67817 128147 67883 128150
rect 66805 127666 66871 127669
rect 95509 127666 95575 127669
rect 66805 127664 68908 127666
rect 66805 127608 66810 127664
rect 66866 127608 68908 127664
rect 66805 127606 68908 127608
rect 94668 127664 95575 127666
rect 94668 127608 95514 127664
rect 95570 127608 95575 127664
rect 94668 127606 95575 127608
rect 66805 127603 66871 127606
rect 95509 127603 95575 127606
rect 192477 127666 192543 127669
rect 192937 127666 193003 127669
rect 192477 127664 193660 127666
rect 192477 127608 192482 127664
rect 192538 127608 192942 127664
rect 192998 127608 193660 127664
rect 192477 127606 193660 127608
rect 192477 127603 192543 127606
rect 192937 127603 193003 127606
rect 226609 127394 226675 127397
rect 224940 127392 226675 127394
rect 224940 127336 226614 127392
rect 226670 127336 226675 127392
rect 224940 127334 226675 127336
rect 226609 127331 226675 127334
rect 97901 127122 97967 127125
rect 94668 127120 97967 127122
rect 94668 127064 97906 127120
rect 97962 127064 97967 127120
rect 94668 127062 97967 127064
rect 97901 127059 97967 127062
rect 68134 126788 68140 126852
rect 68204 126850 68210 126852
rect 68204 126790 68908 126850
rect 68204 126788 68210 126790
rect 191649 126578 191715 126581
rect 226333 126578 226399 126581
rect 191649 126576 193660 126578
rect 191649 126520 191654 126576
rect 191710 126520 193660 126576
rect 191649 126518 193660 126520
rect 224940 126576 226399 126578
rect 224940 126520 226338 126576
rect 226394 126520 226399 126576
rect 224940 126518 226399 126520
rect 191649 126515 191715 126518
rect 226333 126515 226399 126518
rect 97165 126306 97231 126309
rect 94668 126304 97231 126306
rect 94668 126248 97170 126304
rect 97226 126248 97231 126304
rect 94668 126246 97231 126248
rect 97165 126243 97231 126246
rect 66805 126034 66871 126037
rect 580257 126034 580323 126037
rect 583520 126034 584960 126124
rect 66805 126032 68908 126034
rect 66805 125976 66810 126032
rect 66866 125976 68908 126032
rect 66805 125974 68908 125976
rect 580257 126032 584960 126034
rect 580257 125976 580262 126032
rect 580318 125976 584960 126032
rect 580257 125974 584960 125976
rect 66805 125971 66871 125974
rect 580257 125971 580323 125974
rect 583520 125884 584960 125974
rect 193254 125700 193260 125764
rect 193324 125762 193330 125764
rect 226701 125762 226767 125765
rect 193324 125732 193844 125762
rect 224940 125760 226767 125762
rect 193324 125702 193874 125732
rect 224940 125704 226706 125760
rect 226762 125704 226767 125760
rect 224940 125702 226767 125704
rect 193324 125700 193330 125702
rect 193814 125628 193874 125702
rect 226701 125699 226767 125702
rect 69238 125564 69244 125628
rect 69308 125564 69314 125628
rect 193806 125564 193812 125628
rect 193876 125564 193882 125628
rect 69246 125188 69306 125564
rect 94638 124949 94698 125460
rect 94589 124944 94698 124949
rect 94589 124888 94594 124944
rect 94650 124888 94698 124944
rect 94589 124886 94698 124888
rect 94589 124883 94655 124886
rect 97441 124674 97507 124677
rect 94668 124672 97507 124674
rect 94668 124616 97446 124672
rect 97502 124616 97507 124672
rect 94668 124614 97507 124616
rect 97441 124611 97507 124614
rect 66805 124402 66871 124405
rect 66805 124400 68908 124402
rect 66805 124344 66810 124400
rect 66866 124344 68908 124400
rect 66805 124342 68908 124344
rect 66805 124339 66871 124342
rect 97390 124204 97396 124268
rect 97460 124266 97466 124268
rect 104985 124266 105051 124269
rect 97460 124264 105051 124266
rect 97460 124208 104990 124264
rect 105046 124208 105051 124264
rect 97460 124206 105051 124208
rect 97460 124204 97466 124206
rect 104985 124203 105051 124206
rect 184289 124266 184355 124269
rect 192334 124266 192340 124268
rect 184289 124264 192340 124266
rect 184289 124208 184294 124264
rect 184350 124208 192340 124264
rect 184289 124206 192340 124208
rect 184289 124203 184355 124206
rect 192334 124204 192340 124206
rect 192404 124266 192410 124268
rect 193630 124266 193690 124916
rect 226701 124674 226767 124677
rect 224940 124672 226767 124674
rect 224940 124616 226706 124672
rect 226762 124616 226767 124672
rect 224940 124614 226767 124616
rect 226701 124611 226767 124614
rect 192404 124206 193690 124266
rect 192404 124204 192410 124206
rect 95417 124130 95483 124133
rect 94668 124128 95483 124130
rect 94668 124072 95422 124128
rect 95478 124072 95483 124128
rect 94668 124070 95483 124072
rect 95417 124067 95483 124070
rect 66897 123858 66963 123861
rect 191649 123858 191715 123861
rect 225137 123858 225203 123861
rect 66897 123856 68908 123858
rect -960 123572 480 123812
rect 66897 123800 66902 123856
rect 66958 123800 68908 123856
rect 66897 123798 68908 123800
rect 191649 123856 193660 123858
rect 191649 123800 191654 123856
rect 191710 123800 193660 123856
rect 191649 123798 193660 123800
rect 224940 123856 225203 123858
rect 224940 123800 225142 123856
rect 225198 123800 225203 123856
rect 224940 123798 225203 123800
rect 66897 123795 66963 123798
rect 191649 123795 191715 123798
rect 225137 123795 225203 123798
rect 97349 123314 97415 123317
rect 94668 123312 97415 123314
rect 94668 123256 97354 123312
rect 97410 123256 97415 123312
rect 94668 123254 97415 123256
rect 97349 123251 97415 123254
rect 66621 123042 66687 123045
rect 190637 123042 190703 123045
rect 226701 123042 226767 123045
rect 66621 123040 68908 123042
rect 66621 122984 66626 123040
rect 66682 122984 68908 123040
rect 66621 122982 68908 122984
rect 190637 123040 193660 123042
rect 190637 122984 190642 123040
rect 190698 122984 193660 123040
rect 190637 122982 193660 122984
rect 224940 123040 226767 123042
rect 224940 122984 226706 123040
rect 226762 122984 226767 123040
rect 224940 122982 226767 122984
rect 66621 122979 66687 122982
rect 190637 122979 190703 122982
rect 226701 122979 226767 122982
rect 97257 122498 97323 122501
rect 94668 122496 97323 122498
rect 94668 122440 97262 122496
rect 97318 122440 97323 122496
rect 94668 122438 97323 122440
rect 97257 122435 97323 122438
rect 66805 122226 66871 122229
rect 191649 122226 191715 122229
rect 226333 122226 226399 122229
rect 66805 122224 68908 122226
rect 66805 122168 66810 122224
rect 66866 122168 68908 122224
rect 66805 122166 68908 122168
rect 191649 122224 193660 122226
rect 191649 122168 191654 122224
rect 191710 122168 193660 122224
rect 191649 122166 193660 122168
rect 224940 122224 226399 122226
rect 224940 122168 226338 122224
rect 226394 122168 226399 122224
rect 224940 122166 226399 122168
rect 66805 122163 66871 122166
rect 191649 122163 191715 122166
rect 226333 122163 226399 122166
rect 97901 121682 97967 121685
rect 94668 121680 97967 121682
rect 94668 121624 97906 121680
rect 97962 121624 97967 121680
rect 94668 121622 97967 121624
rect 97901 121619 97967 121622
rect 66805 121410 66871 121413
rect 191557 121410 191623 121413
rect 66805 121408 68908 121410
rect 66805 121352 66810 121408
rect 66866 121352 68908 121408
rect 66805 121350 68908 121352
rect 191557 121408 193660 121410
rect 191557 121352 191562 121408
rect 191618 121352 193660 121408
rect 191557 121350 193660 121352
rect 66805 121347 66871 121350
rect 191557 121347 191623 121350
rect 226926 121138 226932 121140
rect 224940 121078 226932 121138
rect 226926 121076 226932 121078
rect 226996 121076 227002 121140
rect 97165 120866 97231 120869
rect 94668 120864 97231 120866
rect 94668 120808 97170 120864
rect 97226 120808 97231 120864
rect 94668 120806 97231 120808
rect 97165 120803 97231 120806
rect 39941 120730 40007 120733
rect 66897 120730 66963 120733
rect 39941 120728 66963 120730
rect 39941 120672 39946 120728
rect 40002 120672 66902 120728
rect 66958 120672 66963 120728
rect 39941 120670 66963 120672
rect 39941 120667 40007 120670
rect 66897 120667 66963 120670
rect 66621 120594 66687 120597
rect 66621 120592 68908 120594
rect 66621 120536 66626 120592
rect 66682 120536 68908 120592
rect 66621 120534 68908 120536
rect 66621 120531 66687 120534
rect 95325 120322 95391 120325
rect 96061 120322 96127 120325
rect 94668 120320 96127 120322
rect 94668 120264 95330 120320
rect 95386 120264 96066 120320
rect 96122 120264 96127 120320
rect 94668 120262 96127 120264
rect 95325 120259 95391 120262
rect 96061 120259 96127 120262
rect 191097 120322 191163 120325
rect 192702 120322 192708 120324
rect 191097 120320 192708 120322
rect 191097 120264 191102 120320
rect 191158 120264 192708 120320
rect 191097 120262 192708 120264
rect 191097 120259 191163 120262
rect 192702 120260 192708 120262
rect 192772 120322 192778 120324
rect 226701 120322 226767 120325
rect 192772 120262 193660 120322
rect 224940 120320 226767 120322
rect 224940 120264 226706 120320
rect 226762 120264 226767 120320
rect 224940 120262 226767 120264
rect 192772 120260 192778 120262
rect 226701 120259 226767 120262
rect 190361 120186 190427 120189
rect 191557 120186 191623 120189
rect 190361 120184 191623 120186
rect 190361 120128 190366 120184
rect 190422 120128 191562 120184
rect 191618 120128 191623 120184
rect 190361 120126 191623 120128
rect 190361 120123 190427 120126
rect 191557 120123 191623 120126
rect 66805 120050 66871 120053
rect 66805 120048 68908 120050
rect 66805 119992 66810 120048
rect 66866 119992 68908 120048
rect 66805 119990 68908 119992
rect 66805 119987 66871 119990
rect 191649 119506 191715 119509
rect 226517 119506 226583 119509
rect 191649 119504 193660 119506
rect 66897 119234 66963 119237
rect 66897 119232 68908 119234
rect 66897 119176 66902 119232
rect 66958 119176 68908 119232
rect 66897 119174 68908 119176
rect 66897 119171 66963 119174
rect 94638 118962 94698 119476
rect 191649 119448 191654 119504
rect 191710 119448 193660 119504
rect 191649 119446 193660 119448
rect 224940 119504 226583 119506
rect 224940 119448 226522 119504
rect 226578 119448 226583 119504
rect 224940 119446 226583 119448
rect 191649 119443 191715 119446
rect 226517 119443 226583 119446
rect 131757 118962 131823 118965
rect 94638 118960 131823 118962
rect 94638 118904 131762 118960
rect 131818 118904 131823 118960
rect 94638 118902 131823 118904
rect 131757 118899 131823 118902
rect 97809 118690 97875 118693
rect 191097 118690 191163 118693
rect 94668 118688 97875 118690
rect 94668 118632 97814 118688
rect 97870 118632 97875 118688
rect 94668 118630 97875 118632
rect 97809 118627 97875 118630
rect 103470 118688 191163 118690
rect 103470 118632 191102 118688
rect 191158 118632 191163 118688
rect 103470 118630 191163 118632
rect 95734 118492 95740 118556
rect 95804 118554 95810 118556
rect 103470 118554 103530 118630
rect 191097 118627 191163 118630
rect 192150 118628 192156 118692
rect 192220 118690 192226 118692
rect 192220 118630 193660 118690
rect 192220 118628 192226 118630
rect 95804 118494 103530 118554
rect 95804 118492 95810 118494
rect 65977 118418 66043 118421
rect 226609 118418 226675 118421
rect 65977 118416 68908 118418
rect 65977 118360 65982 118416
rect 66038 118360 68908 118416
rect 65977 118358 68908 118360
rect 224940 118416 226675 118418
rect 224940 118360 226614 118416
rect 226670 118360 226675 118416
rect 224940 118358 226675 118360
rect 65977 118355 66043 118358
rect 226609 118355 226675 118358
rect 225045 118146 225111 118149
rect 224910 118144 225111 118146
rect 224910 118088 225050 118144
rect 225106 118088 225111 118144
rect 224910 118086 225111 118088
rect 180149 118010 180215 118013
rect 180149 118008 180810 118010
rect 180149 117952 180154 118008
rect 180210 117952 180810 118008
rect 180149 117950 180810 117952
rect 180149 117947 180215 117950
rect 97901 117874 97967 117877
rect 94668 117872 97967 117874
rect 94668 117816 97906 117872
rect 97962 117816 97967 117872
rect 94668 117814 97967 117816
rect 97901 117811 97967 117814
rect 66253 117602 66319 117605
rect 66253 117600 68908 117602
rect 66253 117544 66258 117600
rect 66314 117544 68908 117600
rect 66253 117542 68908 117544
rect 66253 117539 66319 117542
rect 180750 117330 180810 117950
rect 224910 117602 224970 118086
rect 225045 118083 225111 118086
rect 226333 117602 226399 117605
rect 224910 117600 226399 117602
rect 224910 117572 226338 117600
rect 188981 117466 189047 117469
rect 191189 117466 191255 117469
rect 193630 117466 193690 117572
rect 224940 117544 226338 117572
rect 226394 117544 226399 117600
rect 224940 117542 226399 117544
rect 226333 117539 226399 117542
rect 188981 117464 193690 117466
rect 188981 117408 188986 117464
rect 189042 117408 191194 117464
rect 191250 117408 193690 117464
rect 188981 117406 193690 117408
rect 188981 117403 189047 117406
rect 191189 117403 191255 117406
rect 192150 117330 192156 117332
rect 180750 117270 192156 117330
rect 192150 117268 192156 117270
rect 192220 117330 192226 117332
rect 192702 117330 192708 117332
rect 192220 117270 192708 117330
rect 192220 117268 192226 117270
rect 192702 117268 192708 117270
rect 192772 117268 192778 117332
rect 162117 117194 162183 117197
rect 190361 117194 190427 117197
rect 162117 117192 190427 117194
rect 162117 117136 162122 117192
rect 162178 117136 190366 117192
rect 190422 117136 190427 117192
rect 162117 117134 190427 117136
rect 162117 117131 162183 117134
rect 190361 117131 190427 117134
rect 66897 117058 66963 117061
rect 97901 117058 97967 117061
rect 66897 117056 68908 117058
rect 66897 117000 66902 117056
rect 66958 117000 68908 117056
rect 66897 116998 68908 117000
rect 94668 117056 97967 117058
rect 94668 117000 97906 117056
rect 97962 117000 97967 117056
rect 94668 116998 97967 117000
rect 66897 116995 66963 116998
rect 97901 116995 97967 116998
rect 190637 116786 190703 116789
rect 225137 116786 225203 116789
rect 190637 116784 193660 116786
rect 190637 116728 190642 116784
rect 190698 116728 193660 116784
rect 190637 116726 193660 116728
rect 224940 116784 225203 116786
rect 224940 116728 225142 116784
rect 225198 116728 225203 116784
rect 224940 116726 225203 116728
rect 190637 116723 190703 116726
rect 225137 116723 225203 116726
rect 97809 116514 97875 116517
rect 94668 116512 97875 116514
rect 94668 116456 97814 116512
rect 97870 116456 97875 116512
rect 94668 116454 97875 116456
rect 97809 116451 97875 116454
rect 66253 116242 66319 116245
rect 66253 116240 68908 116242
rect 66253 116184 66258 116240
rect 66314 116184 68908 116240
rect 66253 116182 68908 116184
rect 66253 116179 66319 116182
rect 191649 115970 191715 115973
rect 226701 115970 226767 115973
rect 191649 115968 193660 115970
rect 191649 115912 191654 115968
rect 191710 115912 193660 115968
rect 191649 115910 193660 115912
rect 224940 115968 226767 115970
rect 224940 115912 226706 115968
rect 226762 115912 226767 115968
rect 224940 115910 226767 115912
rect 191649 115907 191715 115910
rect 226701 115907 226767 115910
rect 97901 115698 97967 115701
rect 94668 115696 97967 115698
rect 94668 115640 97906 115696
rect 97962 115640 97967 115696
rect 94668 115638 97967 115640
rect 97901 115635 97967 115638
rect 66805 115426 66871 115429
rect 66805 115424 68908 115426
rect 66805 115368 66810 115424
rect 66866 115368 68908 115424
rect 66805 115366 68908 115368
rect 66805 115363 66871 115366
rect 97809 114882 97875 114885
rect 94668 114880 97875 114882
rect 94668 114824 97814 114880
rect 97870 114824 97875 114880
rect 94668 114822 97875 114824
rect 97809 114819 97875 114822
rect 65885 114610 65951 114613
rect 172329 114610 172395 114613
rect 193630 114610 193690 115124
rect 226517 114882 226583 114885
rect 224940 114880 226583 114882
rect 224940 114824 226522 114880
rect 226578 114824 226583 114880
rect 224940 114822 226583 114824
rect 226517 114819 226583 114822
rect 65885 114608 68908 114610
rect 65885 114552 65890 114608
rect 65946 114552 68908 114608
rect 65885 114550 68908 114552
rect 172329 114608 193690 114610
rect 172329 114552 172334 114608
rect 172390 114552 193690 114608
rect 172329 114550 193690 114552
rect 65885 114547 65951 114550
rect 172329 114547 172395 114550
rect 224350 114412 224356 114476
rect 224420 114412 224426 114476
rect 97257 114066 97323 114069
rect 94668 114064 97323 114066
rect 94668 114008 97262 114064
rect 97318 114008 97323 114064
rect 224358 114066 224418 114412
rect 227345 114066 227411 114069
rect 224358 114064 227411 114066
rect 224358 114036 227350 114064
rect 94668 114006 97323 114008
rect 97257 114003 97323 114006
rect 66805 113794 66871 113797
rect 66805 113792 68908 113794
rect 66805 113736 66810 113792
rect 66866 113736 68908 113792
rect 66805 113734 68908 113736
rect 66805 113731 66871 113734
rect 97533 113522 97599 113525
rect 94668 113520 97599 113522
rect 94668 113464 97538 113520
rect 97594 113464 97599 113520
rect 94668 113462 97599 113464
rect 97533 113459 97599 113462
rect 190361 113522 190427 113525
rect 193630 113522 193690 114036
rect 224388 114008 227350 114036
rect 227406 114008 227411 114064
rect 224388 114006 227411 114008
rect 227345 114003 227411 114006
rect 190361 113520 193690 113522
rect 190361 113464 190366 113520
rect 190422 113464 193690 113520
rect 190361 113462 193690 113464
rect 190361 113459 190427 113462
rect 66897 113250 66963 113253
rect 191005 113250 191071 113253
rect 227805 113250 227871 113253
rect 66897 113248 68908 113250
rect 66897 113192 66902 113248
rect 66958 113192 68908 113248
rect 66897 113190 68908 113192
rect 191005 113248 193660 113250
rect 191005 113192 191010 113248
rect 191066 113192 193660 113248
rect 191005 113190 193660 113192
rect 224940 113248 227871 113250
rect 224940 113192 227810 113248
rect 227866 113192 227871 113248
rect 224940 113190 227871 113192
rect 66897 113187 66963 113190
rect 191005 113187 191071 113190
rect 227805 113187 227871 113190
rect 237966 113114 237972 113116
rect 229050 113054 237972 113114
rect 229050 112842 229110 113054
rect 237966 113052 237972 113054
rect 238036 113052 238042 113116
rect 224910 112782 229110 112842
rect 582833 112842 582899 112845
rect 583520 112842 584960 112932
rect 582833 112840 584960 112842
rect 582833 112784 582838 112840
rect 582894 112784 584960 112840
rect 582833 112782 584960 112784
rect 97809 112706 97875 112709
rect 94668 112704 97875 112706
rect 94668 112648 97814 112704
rect 97870 112648 97875 112704
rect 94668 112646 97875 112648
rect 97809 112643 97875 112646
rect 67633 112434 67699 112437
rect 191741 112434 191807 112437
rect 67633 112432 68908 112434
rect 67633 112376 67638 112432
rect 67694 112376 68908 112432
rect 67633 112374 68908 112376
rect 191741 112432 193660 112434
rect 191741 112376 191746 112432
rect 191802 112376 193660 112432
rect 191741 112374 193660 112376
rect 67633 112371 67699 112374
rect 191741 112371 191807 112374
rect 224910 112132 224970 112782
rect 582833 112779 582899 112782
rect 583520 112692 584960 112782
rect 97901 111890 97967 111893
rect 94668 111888 97967 111890
rect 94668 111832 97906 111888
rect 97962 111832 97967 111888
rect 94668 111830 97967 111832
rect 97901 111827 97967 111830
rect 237966 111828 237972 111892
rect 238036 111890 238042 111892
rect 238109 111890 238175 111893
rect 238036 111888 238175 111890
rect 238036 111832 238114 111888
rect 238170 111832 238175 111888
rect 238036 111830 238175 111832
rect 238036 111828 238042 111830
rect 238109 111827 238175 111830
rect 240685 111892 240751 111893
rect 240685 111888 240732 111892
rect 240796 111890 240802 111892
rect 240685 111832 240690 111888
rect 240685 111828 240732 111832
rect 240796 111830 240842 111890
rect 240796 111828 240802 111830
rect 240685 111827 240751 111828
rect 66161 111618 66227 111621
rect 66161 111616 68908 111618
rect 66161 111560 66166 111616
rect 66222 111560 68908 111616
rect 66161 111558 68908 111560
rect 66161 111555 66227 111558
rect 225321 111346 225387 111349
rect 224940 111344 225387 111346
rect 96797 111074 96863 111077
rect 94668 111072 96863 111074
rect 94668 111016 96802 111072
rect 96858 111016 96863 111072
rect 94668 111014 96863 111016
rect 96797 111011 96863 111014
rect 66621 110802 66687 110805
rect 190361 110802 190427 110805
rect 193630 110802 193690 111316
rect 224940 111288 225326 111344
rect 225382 111288 225387 111344
rect 224940 111286 225387 111288
rect 225321 111283 225387 111286
rect 66621 110800 68908 110802
rect -960 110666 480 110756
rect 66621 110744 66626 110800
rect 66682 110744 68908 110800
rect 66621 110742 68908 110744
rect 190361 110800 193690 110802
rect 190361 110744 190366 110800
rect 190422 110744 193690 110800
rect 190361 110742 193690 110744
rect 66621 110739 66687 110742
rect 190361 110739 190427 110742
rect 3141 110666 3207 110669
rect -960 110664 3207 110666
rect -960 110608 3146 110664
rect 3202 110608 3207 110664
rect -960 110606 3207 110608
rect -960 110516 480 110606
rect 3141 110603 3207 110606
rect 191741 110530 191807 110533
rect 226517 110530 226583 110533
rect 191741 110528 193660 110530
rect 191741 110472 191746 110528
rect 191802 110472 193660 110528
rect 191741 110470 193660 110472
rect 224940 110528 226583 110530
rect 224940 110472 226522 110528
rect 226578 110472 226583 110528
rect 224940 110470 226583 110472
rect 191741 110467 191807 110470
rect 226517 110467 226583 110470
rect 66805 110258 66871 110261
rect 97441 110258 97507 110261
rect 66805 110256 68908 110258
rect 66805 110200 66810 110256
rect 66866 110200 68908 110256
rect 66805 110198 68908 110200
rect 94668 110256 97507 110258
rect 94668 110200 97446 110256
rect 97502 110200 97507 110256
rect 94668 110198 97507 110200
rect 66805 110195 66871 110198
rect 97441 110195 97507 110198
rect 97165 109714 97231 109717
rect 94668 109712 97231 109714
rect 94668 109656 97170 109712
rect 97226 109656 97231 109712
rect 94668 109654 97231 109656
rect 97165 109651 97231 109654
rect 191557 109714 191623 109717
rect 227805 109714 227871 109717
rect 191557 109712 193660 109714
rect 191557 109656 191562 109712
rect 191618 109656 193660 109712
rect 191557 109654 193660 109656
rect 224940 109712 227871 109714
rect 224940 109656 227810 109712
rect 227866 109656 227871 109712
rect 224940 109654 227871 109656
rect 191557 109651 191623 109654
rect 227805 109651 227871 109654
rect 66478 109380 66484 109444
rect 66548 109442 66554 109444
rect 66548 109382 68908 109442
rect 66548 109380 66554 109382
rect 182081 109170 182147 109173
rect 186814 109170 186820 109172
rect 182081 109168 186820 109170
rect 182081 109112 182086 109168
rect 182142 109112 186820 109168
rect 182081 109110 186820 109112
rect 182081 109107 182147 109110
rect 186814 109108 186820 109110
rect 186884 109108 186890 109172
rect 159449 109034 159515 109037
rect 160001 109034 160067 109037
rect 190361 109034 190427 109037
rect 159449 109032 190427 109034
rect 159449 108976 159454 109032
rect 159510 108976 160006 109032
rect 160062 108976 190366 109032
rect 190422 108976 190427 109032
rect 159449 108974 190427 108976
rect 159449 108971 159515 108974
rect 160001 108971 160067 108974
rect 190361 108971 190427 108974
rect 97942 108898 97948 108900
rect 94668 108838 97948 108898
rect 97942 108836 97948 108838
rect 98012 108836 98018 108900
rect 66805 108626 66871 108629
rect 66805 108624 68908 108626
rect 66805 108568 66810 108624
rect 66866 108568 68908 108624
rect 66805 108566 68908 108568
rect 66805 108563 66871 108566
rect 186129 108218 186195 108221
rect 193630 108218 193690 108868
rect 226609 108626 226675 108629
rect 224940 108624 226675 108626
rect 224940 108568 226614 108624
rect 226670 108568 226675 108624
rect 224940 108566 226675 108568
rect 226609 108563 226675 108566
rect 186129 108216 193690 108218
rect 186129 108160 186134 108216
rect 186190 108160 193690 108216
rect 186129 108158 193690 108160
rect 186129 108155 186195 108158
rect 97901 108082 97967 108085
rect 94668 108080 97967 108082
rect 94668 108024 97906 108080
rect 97962 108024 97967 108080
rect 94668 108022 97967 108024
rect 97901 108019 97967 108022
rect 66897 107810 66963 107813
rect 191741 107810 191807 107813
rect 226701 107810 226767 107813
rect 66897 107808 68908 107810
rect 66897 107752 66902 107808
rect 66958 107752 68908 107808
rect 66897 107750 68908 107752
rect 191741 107808 193660 107810
rect 191741 107752 191746 107808
rect 191802 107752 193660 107808
rect 191741 107750 193660 107752
rect 224940 107808 226767 107810
rect 224940 107752 226706 107808
rect 226762 107752 226767 107808
rect 224940 107750 226767 107752
rect 66897 107747 66963 107750
rect 191741 107747 191807 107750
rect 226701 107747 226767 107750
rect 97533 107266 97599 107269
rect 94668 107264 97599 107266
rect 94668 107208 97538 107264
rect 97594 107208 97599 107264
rect 94668 107206 97599 107208
rect 97533 107203 97599 107206
rect 66805 106994 66871 106997
rect 191557 106994 191623 106997
rect 226701 106994 226767 106997
rect 66805 106992 68908 106994
rect 66805 106936 66810 106992
rect 66866 106936 68908 106992
rect 66805 106934 68908 106936
rect 191557 106992 193660 106994
rect 191557 106936 191562 106992
rect 191618 106936 193660 106992
rect 191557 106934 193660 106936
rect 224940 106992 226767 106994
rect 224940 106936 226706 106992
rect 226762 106936 226767 106992
rect 224940 106934 226767 106936
rect 66805 106931 66871 106934
rect 191557 106931 191623 106934
rect 226701 106931 226767 106934
rect 97901 106722 97967 106725
rect 94668 106720 97967 106722
rect 94668 106664 97906 106720
rect 97962 106664 97967 106720
rect 94668 106662 97967 106664
rect 97901 106659 97967 106662
rect 66897 106450 66963 106453
rect 66897 106448 68908 106450
rect 66897 106392 66902 106448
rect 66958 106392 68908 106448
rect 66897 106390 68908 106392
rect 66897 106387 66963 106390
rect 191741 106178 191807 106181
rect 191741 106176 193660 106178
rect 191741 106120 191746 106176
rect 191802 106120 193660 106176
rect 191741 106118 193660 106120
rect 191741 106115 191807 106118
rect 97901 105906 97967 105909
rect 226333 105906 226399 105909
rect 94668 105904 97967 105906
rect 94668 105848 97906 105904
rect 97962 105848 97967 105904
rect 94668 105846 97967 105848
rect 224940 105904 226399 105906
rect 224940 105848 226338 105904
rect 226394 105848 226399 105904
rect 224940 105846 226399 105848
rect 97901 105843 97967 105846
rect 226333 105843 226399 105846
rect 66529 105634 66595 105637
rect 66529 105632 68908 105634
rect 66529 105576 66534 105632
rect 66590 105576 68908 105632
rect 66529 105574 68908 105576
rect 66529 105571 66595 105574
rect 97533 105090 97599 105093
rect 94668 105088 97599 105090
rect 94668 105032 97538 105088
rect 97594 105032 97599 105088
rect 94668 105030 97599 105032
rect 97533 105027 97599 105030
rect 190453 105090 190519 105093
rect 226609 105090 226675 105093
rect 190453 105088 193660 105090
rect 190453 105032 190458 105088
rect 190514 105032 193660 105088
rect 190453 105030 193660 105032
rect 224940 105088 226675 105090
rect 224940 105032 226614 105088
rect 226670 105032 226675 105088
rect 224940 105030 226675 105032
rect 190453 105027 190519 105030
rect 226609 105027 226675 105030
rect 66253 104818 66319 104821
rect 66253 104816 68908 104818
rect 66253 104760 66258 104816
rect 66314 104760 68908 104816
rect 66253 104758 68908 104760
rect 66253 104755 66319 104758
rect 97901 104274 97967 104277
rect 94668 104272 97967 104274
rect 94668 104216 97906 104272
rect 97962 104216 97967 104272
rect 94668 104214 97967 104216
rect 97901 104211 97967 104214
rect 191649 104274 191715 104277
rect 226517 104274 226583 104277
rect 191649 104272 193660 104274
rect 191649 104216 191654 104272
rect 191710 104216 193660 104272
rect 191649 104214 193660 104216
rect 224940 104272 226583 104274
rect 224940 104216 226522 104272
rect 226578 104216 226583 104272
rect 224940 104214 226583 104216
rect 191649 104211 191715 104214
rect 226517 104211 226583 104214
rect 66662 103940 66668 104004
rect 66732 104002 66738 104004
rect 66732 103942 68908 104002
rect 66732 103940 66738 103942
rect 97717 103458 97783 103461
rect 94668 103456 97783 103458
rect 94668 103400 97722 103456
rect 97778 103400 97783 103456
rect 94668 103398 97783 103400
rect 97717 103395 97783 103398
rect 191005 103458 191071 103461
rect 226609 103458 226675 103461
rect 191005 103456 193660 103458
rect 191005 103400 191010 103456
rect 191066 103400 193660 103456
rect 191005 103398 193660 103400
rect 224940 103456 226675 103458
rect 224940 103400 226614 103456
rect 226670 103400 226675 103456
rect 224940 103398 226675 103400
rect 191005 103395 191071 103398
rect 226609 103395 226675 103398
rect 66069 103186 66135 103189
rect 66069 103184 68908 103186
rect 66069 103128 66074 103184
rect 66130 103128 68908 103184
rect 66069 103126 68908 103128
rect 66069 103123 66135 103126
rect 97901 102914 97967 102917
rect 94668 102912 97967 102914
rect 94668 102856 97906 102912
rect 97962 102856 97967 102912
rect 94668 102854 97967 102856
rect 97901 102851 97967 102854
rect 226241 102778 226307 102781
rect 249057 102778 249123 102781
rect 226241 102776 249123 102778
rect 226241 102720 226246 102776
rect 226302 102720 249062 102776
rect 249118 102720 249123 102776
rect 226241 102718 249123 102720
rect 226241 102715 226307 102718
rect 249057 102715 249123 102718
rect 66529 102642 66595 102645
rect 66529 102640 68908 102642
rect 66529 102584 66534 102640
rect 66590 102584 68908 102640
rect 66529 102582 68908 102584
rect 66529 102579 66595 102582
rect 100109 102234 100175 102237
rect 193630 102234 193690 102612
rect 225229 102370 225295 102373
rect 227897 102370 227963 102373
rect 224940 102368 227963 102370
rect 224940 102312 225234 102368
rect 225290 102312 227902 102368
rect 227958 102312 227963 102368
rect 224940 102310 227963 102312
rect 225229 102307 225295 102310
rect 227897 102307 227963 102310
rect 100109 102232 193690 102234
rect 100109 102176 100114 102232
rect 100170 102176 193690 102232
rect 100109 102174 193690 102176
rect 100109 102171 100175 102174
rect 97625 102098 97691 102101
rect 94668 102096 97691 102098
rect 94668 102040 97630 102096
rect 97686 102040 97691 102096
rect 94668 102038 97691 102040
rect 97625 102035 97691 102038
rect 66805 101826 66871 101829
rect 66805 101824 68908 101826
rect 66805 101768 66810 101824
rect 66866 101768 68908 101824
rect 66805 101766 68908 101768
rect 66805 101763 66871 101766
rect 190637 101554 190703 101557
rect 226701 101554 226767 101557
rect 190637 101552 193660 101554
rect 190637 101496 190642 101552
rect 190698 101496 193660 101552
rect 190637 101494 193660 101496
rect 224940 101552 226767 101554
rect 224940 101496 226706 101552
rect 226762 101496 226767 101552
rect 224940 101494 226767 101496
rect 190637 101491 190703 101494
rect 226701 101491 226767 101494
rect 97901 101282 97967 101285
rect 94668 101280 97967 101282
rect 94668 101224 97906 101280
rect 97962 101224 97967 101280
rect 94668 101222 97967 101224
rect 97901 101219 97967 101222
rect 66437 101010 66503 101013
rect 66437 101008 68908 101010
rect 66437 100952 66442 101008
rect 66498 100952 68908 101008
rect 66437 100950 68908 100952
rect 66437 100947 66503 100950
rect 191649 100738 191715 100741
rect 193397 100738 193463 100741
rect 226241 100738 226307 100741
rect 191649 100736 193660 100738
rect 191649 100680 191654 100736
rect 191710 100680 193402 100736
rect 193458 100680 193660 100736
rect 191649 100678 193660 100680
rect 224940 100736 226307 100738
rect 224940 100680 226246 100736
rect 226302 100680 226307 100736
rect 224940 100678 226307 100680
rect 191649 100675 191715 100678
rect 193397 100675 193463 100678
rect 226241 100675 226307 100678
rect 97809 100466 97875 100469
rect 94668 100464 97875 100466
rect 94668 100408 97814 100464
rect 97870 100408 97875 100464
rect 94668 100406 97875 100408
rect 97809 100403 97875 100406
rect 69430 99924 69490 100164
rect 69422 99860 69428 99924
rect 69492 99860 69498 99924
rect 190637 99922 190703 99925
rect 190637 99920 193660 99922
rect 190637 99864 190642 99920
rect 190698 99864 193660 99920
rect 190637 99862 193660 99864
rect 190637 99859 190703 99862
rect 66805 99650 66871 99653
rect 97901 99650 97967 99653
rect 227529 99650 227595 99653
rect 66805 99648 68908 99650
rect 66805 99592 66810 99648
rect 66866 99592 68908 99648
rect 66805 99590 68908 99592
rect 94668 99648 97967 99650
rect 94668 99592 97906 99648
rect 97962 99592 97967 99648
rect 94668 99590 97967 99592
rect 224940 99648 227595 99650
rect 224940 99592 227534 99648
rect 227590 99592 227595 99648
rect 224940 99590 227595 99592
rect 66805 99587 66871 99590
rect 97901 99587 97967 99590
rect 227529 99587 227595 99590
rect 582373 99514 582439 99517
rect 583520 99514 584960 99604
rect 582373 99512 584960 99514
rect 582373 99456 582378 99512
rect 582434 99456 584960 99512
rect 582373 99454 584960 99456
rect 582373 99451 582439 99454
rect 583520 99364 584960 99454
rect 97533 99106 97599 99109
rect 94668 99104 97599 99106
rect 94668 99048 97538 99104
rect 97594 99048 97599 99104
rect 94668 99046 97599 99048
rect 97533 99043 97599 99046
rect 66621 98834 66687 98837
rect 190821 98834 190887 98837
rect 66621 98832 68908 98834
rect 66621 98776 66626 98832
rect 66682 98776 68908 98832
rect 66621 98774 68908 98776
rect 190821 98832 193660 98834
rect 190821 98776 190826 98832
rect 190882 98776 193660 98832
rect 190821 98774 193660 98776
rect 66621 98771 66687 98774
rect 190821 98771 190887 98774
rect 97809 98290 97875 98293
rect 94668 98288 97875 98290
rect 94668 98232 97814 98288
rect 97870 98232 97875 98288
rect 94668 98230 97875 98232
rect 224910 98290 224970 98804
rect 225086 98290 225092 98292
rect 224910 98230 225092 98290
rect 97809 98227 97875 98230
rect 225086 98228 225092 98230
rect 225156 98228 225162 98292
rect 67173 98018 67239 98021
rect 191741 98018 191807 98021
rect 225137 98018 225203 98021
rect 226149 98018 226215 98021
rect 67173 98016 68908 98018
rect 67173 97960 67178 98016
rect 67234 97960 68908 98016
rect 67173 97958 68908 97960
rect 191741 98016 193660 98018
rect 191741 97960 191746 98016
rect 191802 97960 193660 98016
rect 191741 97958 193660 97960
rect 224940 98016 226215 98018
rect 224940 97960 225142 98016
rect 225198 97960 226154 98016
rect 226210 97960 226215 98016
rect 224940 97958 226215 97960
rect 67173 97955 67239 97958
rect 191741 97955 191807 97958
rect 225137 97955 225203 97958
rect 226149 97955 226215 97958
rect -960 97610 480 97700
rect 3049 97610 3115 97613
rect -960 97608 3115 97610
rect -960 97552 3054 97608
rect 3110 97552 3115 97608
rect -960 97550 3115 97552
rect -960 97460 480 97550
rect 3049 97547 3115 97550
rect 97901 97474 97967 97477
rect 94668 97472 97967 97474
rect 94668 97416 97906 97472
rect 97962 97416 97967 97472
rect 94668 97414 97967 97416
rect 97901 97411 97967 97414
rect 67357 97202 67423 97205
rect 226374 97202 226380 97204
rect 67357 97200 68908 97202
rect 67357 97144 67362 97200
rect 67418 97144 68908 97200
rect 67357 97142 68908 97144
rect 67357 97139 67423 97142
rect 96613 96658 96679 96661
rect 94668 96656 96679 96658
rect 94668 96600 96618 96656
rect 96674 96600 96679 96656
rect 94668 96598 96679 96600
rect 96613 96595 96679 96598
rect 184790 96596 184796 96660
rect 184860 96658 184866 96660
rect 193630 96658 193690 97172
rect 224940 97142 226380 97202
rect 226374 97140 226380 97142
rect 226444 97202 226450 97204
rect 226609 97202 226675 97205
rect 226444 97200 226675 97202
rect 226444 97144 226614 97200
rect 226670 97144 226675 97200
rect 226444 97142 226675 97144
rect 226444 97140 226450 97142
rect 226609 97139 226675 97142
rect 184860 96598 193690 96658
rect 184860 96596 184866 96598
rect 66621 96386 66687 96389
rect 191557 96386 191623 96389
rect 66621 96384 68908 96386
rect 66621 96328 66626 96384
rect 66682 96328 68908 96384
rect 66621 96326 68908 96328
rect 191557 96384 193660 96386
rect 191557 96328 191562 96384
rect 191618 96328 193660 96384
rect 191557 96326 193660 96328
rect 66621 96323 66687 96326
rect 191557 96323 191623 96326
rect 99005 96114 99071 96117
rect 226425 96114 226491 96117
rect 94668 96112 99071 96114
rect 94668 96056 99010 96112
rect 99066 96056 99071 96112
rect 94668 96054 99071 96056
rect 224940 96112 226491 96114
rect 224940 96056 226430 96112
rect 226486 96056 226491 96112
rect 224940 96054 226491 96056
rect 99005 96051 99071 96054
rect 226425 96051 226491 96054
rect 55029 95842 55095 95845
rect 66846 95842 66852 95844
rect 55029 95840 66852 95842
rect 55029 95784 55034 95840
rect 55090 95784 66852 95840
rect 55029 95782 66852 95784
rect 55029 95779 55095 95782
rect 66846 95780 66852 95782
rect 66916 95780 66922 95844
rect 67449 95842 67515 95845
rect 67449 95840 68908 95842
rect 67449 95784 67454 95840
rect 67510 95784 68908 95840
rect 67449 95782 68908 95784
rect 67449 95779 67515 95782
rect 97901 95298 97967 95301
rect 226609 95300 226675 95301
rect 94668 95296 97967 95298
rect 94668 95240 97906 95296
rect 97962 95240 97967 95296
rect 94668 95238 97967 95240
rect 97901 95235 97967 95238
rect 188838 95236 188844 95300
rect 188908 95298 188914 95300
rect 226558 95298 226564 95300
rect 188908 95238 193660 95298
rect 224940 95238 226564 95298
rect 226628 95296 226675 95300
rect 226670 95240 226675 95296
rect 188908 95236 188914 95238
rect 226558 95236 226564 95238
rect 226628 95236 226675 95240
rect 226609 95235 226675 95236
rect 66846 94964 66852 95028
rect 66916 95026 66922 95028
rect 66916 94966 68908 95026
rect 66916 94964 66922 94966
rect 97809 94482 97875 94485
rect 94668 94480 97875 94482
rect 94668 94424 97814 94480
rect 97870 94424 97875 94480
rect 94668 94422 97875 94424
rect 97809 94419 97875 94422
rect 191649 94482 191715 94485
rect 226701 94482 226767 94485
rect 191649 94480 193660 94482
rect 191649 94424 191654 94480
rect 191710 94424 193660 94480
rect 224388 94480 226767 94482
rect 224388 94452 226706 94480
rect 191649 94422 193660 94424
rect 224358 94424 226706 94452
rect 226762 94424 226767 94480
rect 224358 94422 226767 94424
rect 191649 94419 191715 94422
rect 224358 94348 224418 94422
rect 226701 94419 226767 94422
rect 224350 94284 224356 94348
rect 224420 94284 224426 94348
rect 67541 94210 67607 94213
rect 67541 94208 68908 94210
rect 67541 94152 67546 94208
rect 67602 94152 68908 94208
rect 67541 94150 68908 94152
rect 67541 94147 67607 94150
rect 226977 93666 227043 93669
rect 224940 93664 227043 93666
rect 67817 93394 67883 93397
rect 67817 93392 68908 93394
rect 67817 93336 67822 93392
rect 67878 93336 68908 93392
rect 67817 93334 68908 93336
rect 67817 93331 67883 93334
rect 94638 93122 94698 93636
rect 94638 93062 103530 93122
rect 97206 92850 97212 92852
rect 94668 92790 97212 92850
rect 97206 92788 97212 92790
rect 97276 92788 97282 92852
rect 72969 92716 73035 92717
rect 72918 92652 72924 92716
rect 72988 92714 73035 92716
rect 93255 92714 93321 92717
rect 93710 92714 93716 92716
rect 72988 92712 73080 92714
rect 73030 92656 73080 92712
rect 72988 92654 73080 92656
rect 93255 92712 93716 92714
rect 93255 92656 93260 92712
rect 93316 92656 93716 92712
rect 93255 92654 93716 92656
rect 72988 92652 73035 92654
rect 72969 92651 73035 92652
rect 93255 92651 93321 92654
rect 93710 92652 93716 92654
rect 93780 92652 93786 92716
rect 103470 92578 103530 93062
rect 194182 92986 194242 93636
rect 224940 93608 226982 93664
rect 227038 93608 227043 93664
rect 224940 93606 227043 93608
rect 226977 93603 227043 93606
rect 215334 93332 215340 93396
rect 215404 93394 215410 93396
rect 216121 93394 216187 93397
rect 215404 93392 216187 93394
rect 215404 93336 216126 93392
rect 216182 93336 216187 93392
rect 215404 93334 216187 93336
rect 215404 93332 215410 93334
rect 216121 93331 216187 93334
rect 224493 93394 224559 93397
rect 224902 93394 224908 93396
rect 224493 93392 224908 93394
rect 224493 93336 224498 93392
rect 224554 93336 224908 93392
rect 224493 93334 224908 93336
rect 224493 93331 224559 93334
rect 224902 93332 224908 93334
rect 224972 93332 224978 93396
rect 229737 93122 229803 93125
rect 200070 93120 229803 93122
rect 200070 93064 229742 93120
rect 229798 93064 229803 93120
rect 200070 93062 229803 93064
rect 200070 92986 200130 93062
rect 201401 92988 201467 92989
rect 201350 92986 201356 92988
rect 194182 92926 200130 92986
rect 201310 92926 201356 92986
rect 201420 92984 201467 92988
rect 201462 92928 201467 92984
rect 201350 92924 201356 92926
rect 201420 92924 201467 92928
rect 201401 92923 201467 92924
rect 193857 92850 193923 92853
rect 193990 92850 193996 92852
rect 193857 92848 193996 92850
rect 193857 92792 193862 92848
rect 193918 92792 193996 92848
rect 193857 92790 193996 92792
rect 193857 92787 193923 92790
rect 193990 92788 193996 92790
rect 194060 92788 194066 92852
rect 195513 92850 195579 92853
rect 195830 92850 195836 92852
rect 195513 92848 195836 92850
rect 195513 92792 195518 92848
rect 195574 92792 195836 92848
rect 195513 92790 195836 92792
rect 195513 92787 195579 92790
rect 195830 92788 195836 92790
rect 195900 92788 195906 92852
rect 200481 92850 200547 92853
rect 201585 92852 201651 92853
rect 200614 92850 200620 92852
rect 200481 92848 200620 92850
rect 200481 92792 200486 92848
rect 200542 92792 200620 92848
rect 200481 92790 200620 92792
rect 200481 92787 200547 92790
rect 200614 92788 200620 92790
rect 200684 92788 200690 92852
rect 201534 92850 201540 92852
rect 201494 92790 201540 92850
rect 201604 92848 201651 92852
rect 201646 92792 201651 92848
rect 201534 92788 201540 92790
rect 201604 92788 201651 92792
rect 201585 92787 201651 92788
rect 204670 92717 204730 93062
rect 229737 93059 229803 93062
rect 207105 92852 207171 92853
rect 208761 92852 208827 92853
rect 207054 92850 207060 92852
rect 207014 92790 207060 92850
rect 207124 92848 207171 92852
rect 208710 92850 208716 92852
rect 207166 92792 207171 92848
rect 207054 92788 207060 92790
rect 207124 92788 207171 92792
rect 208670 92790 208716 92850
rect 208780 92848 208827 92852
rect 208822 92792 208827 92848
rect 208710 92788 208716 92790
rect 208780 92788 208827 92792
rect 209814 92788 209820 92852
rect 209884 92850 209890 92852
rect 210049 92850 210115 92853
rect 209884 92848 210115 92850
rect 209884 92792 210054 92848
rect 210110 92792 210115 92848
rect 209884 92790 210115 92792
rect 209884 92788 209890 92790
rect 207105 92787 207171 92788
rect 208761 92787 208827 92788
rect 210049 92787 210115 92790
rect 213637 92852 213703 92853
rect 213637 92848 213684 92852
rect 213748 92850 213754 92852
rect 213637 92792 213642 92848
rect 213637 92788 213684 92792
rect 213748 92790 213794 92850
rect 213748 92788 213754 92790
rect 213637 92787 213703 92788
rect 204621 92712 204730 92717
rect 204621 92656 204626 92712
rect 204682 92656 204730 92712
rect 204621 92654 204730 92656
rect 204621 92651 204687 92654
rect 204846 92652 204852 92716
rect 204916 92714 204922 92716
rect 205081 92714 205147 92717
rect 204916 92712 205147 92714
rect 204916 92656 205086 92712
rect 205142 92656 205147 92712
rect 204916 92654 205147 92656
rect 204916 92652 204922 92654
rect 205081 92651 205147 92654
rect 125593 92578 125659 92581
rect 103470 92576 125659 92578
rect 103470 92520 125598 92576
rect 125654 92520 125659 92576
rect 103470 92518 125659 92520
rect 125593 92515 125659 92518
rect 64597 92442 64663 92445
rect 76281 92442 76347 92445
rect 64597 92440 76347 92442
rect 64597 92384 64602 92440
rect 64658 92384 76286 92440
rect 76342 92384 76347 92440
rect 64597 92382 76347 92384
rect 64597 92379 64663 92382
rect 76281 92379 76347 92382
rect 91001 92442 91067 92445
rect 91686 92442 91692 92444
rect 91001 92440 91692 92442
rect 91001 92384 91006 92440
rect 91062 92384 91692 92440
rect 91001 92382 91692 92384
rect 91001 92379 91067 92382
rect 91686 92380 91692 92382
rect 91756 92380 91762 92444
rect 92381 92442 92447 92445
rect 94773 92442 94839 92445
rect 92381 92440 94839 92442
rect 92381 92384 92386 92440
rect 92442 92384 94778 92440
rect 94834 92384 94839 92440
rect 92381 92382 94839 92384
rect 92381 92379 92447 92382
rect 94773 92379 94839 92382
rect 99005 92442 99071 92445
rect 166165 92442 166231 92445
rect 99005 92440 166231 92442
rect 99005 92384 99010 92440
rect 99066 92384 166170 92440
rect 166226 92384 166231 92440
rect 99005 92382 166231 92384
rect 99005 92379 99071 92382
rect 166165 92379 166231 92382
rect 176561 92442 176627 92445
rect 196525 92442 196591 92445
rect 176561 92440 196591 92442
rect 176561 92384 176566 92440
rect 176622 92384 196530 92440
rect 196586 92384 196591 92440
rect 176561 92382 196591 92384
rect 176561 92379 176627 92382
rect 196525 92379 196591 92382
rect 203190 92380 203196 92444
rect 203260 92442 203266 92444
rect 204161 92442 204227 92445
rect 203260 92440 204227 92442
rect 203260 92384 204166 92440
rect 204222 92384 204227 92440
rect 203260 92382 204227 92384
rect 203260 92380 203266 92382
rect 204161 92379 204227 92382
rect 223573 92442 223639 92445
rect 226558 92442 226564 92444
rect 223573 92440 226564 92442
rect 223573 92384 223578 92440
rect 223634 92384 226564 92440
rect 223573 92382 226564 92384
rect 223573 92379 223639 92382
rect 226558 92380 226564 92382
rect 226628 92380 226634 92444
rect 91829 92306 91895 92309
rect 98729 92306 98795 92309
rect 91829 92304 98795 92306
rect 91829 92248 91834 92304
rect 91890 92248 98734 92304
rect 98790 92248 98795 92304
rect 91829 92246 98795 92248
rect 91829 92243 91895 92246
rect 98729 92243 98795 92246
rect 186814 92244 186820 92308
rect 186884 92306 186890 92308
rect 193029 92306 193095 92309
rect 186884 92304 193095 92306
rect 186884 92248 193034 92304
rect 193090 92248 193095 92304
rect 186884 92246 193095 92248
rect 186884 92244 186890 92246
rect 193029 92243 193095 92246
rect 203517 92306 203583 92309
rect 241329 92306 241395 92309
rect 203517 92304 241395 92306
rect 203517 92248 203522 92304
rect 203578 92248 241334 92304
rect 241390 92248 241395 92304
rect 203517 92246 241395 92248
rect 203517 92243 203583 92246
rect 241329 92243 241395 92246
rect 79501 92170 79567 92173
rect 97390 92170 97396 92172
rect 79501 92168 97396 92170
rect 79501 92112 79506 92168
rect 79562 92112 97396 92168
rect 79501 92110 97396 92112
rect 79501 92107 79567 92110
rect 97390 92108 97396 92110
rect 97460 92108 97466 92172
rect 191833 92170 191899 92173
rect 224350 92170 224356 92172
rect 191833 92168 224356 92170
rect 191833 92112 191838 92168
rect 191894 92112 224356 92168
rect 191833 92110 224356 92112
rect 191833 92107 191899 92110
rect 224350 92108 224356 92110
rect 224420 92108 224426 92172
rect 197997 92034 198063 92037
rect 249793 92034 249859 92037
rect 197997 92032 249859 92034
rect 197997 91976 198002 92032
rect 198058 91976 249798 92032
rect 249854 91976 249859 92032
rect 197997 91974 249859 91976
rect 197997 91971 198063 91974
rect 249793 91971 249859 91974
rect 190310 91836 190316 91900
rect 190380 91898 190386 91900
rect 200757 91898 200823 91901
rect 190380 91896 200823 91898
rect 190380 91840 200762 91896
rect 200818 91840 200823 91896
rect 190380 91838 200823 91840
rect 190380 91836 190386 91838
rect 200757 91835 200823 91838
rect 41229 91762 41295 91765
rect 68001 91762 68067 91765
rect 41229 91760 68067 91762
rect 41229 91704 41234 91760
rect 41290 91704 68006 91760
rect 68062 91704 68067 91760
rect 41229 91702 68067 91704
rect 41229 91699 41295 91702
rect 68001 91699 68067 91702
rect 70301 91218 70367 91221
rect 71037 91218 71103 91221
rect 70301 91216 71103 91218
rect 70301 91160 70306 91216
rect 70362 91160 71042 91216
rect 71098 91160 71103 91216
rect 70301 91158 71103 91160
rect 70301 91155 70367 91158
rect 71037 91155 71103 91158
rect 192334 91156 192340 91220
rect 192404 91218 192410 91220
rect 193029 91218 193095 91221
rect 192404 91216 193095 91218
rect 192404 91160 193034 91216
rect 193090 91160 193095 91216
rect 192404 91158 193095 91160
rect 192404 91156 192410 91158
rect 193029 91155 193095 91158
rect 68001 91082 68067 91085
rect 71129 91082 71195 91085
rect 68001 91080 71195 91082
rect 68001 91024 68006 91080
rect 68062 91024 71134 91080
rect 71190 91024 71195 91080
rect 68001 91022 71195 91024
rect 68001 91019 68067 91022
rect 71129 91019 71195 91022
rect 71630 91020 71636 91084
rect 71700 91082 71706 91084
rect 74809 91082 74875 91085
rect 100753 91084 100819 91085
rect 100702 91082 100708 91084
rect 71700 91080 74875 91082
rect 71700 91024 74814 91080
rect 74870 91024 74875 91080
rect 71700 91022 74875 91024
rect 100662 91022 100708 91082
rect 100772 91080 100819 91084
rect 100814 91024 100819 91080
rect 71700 91020 71706 91022
rect 74809 91019 74875 91022
rect 100702 91020 100708 91022
rect 100772 91020 100819 91024
rect 100753 91019 100819 91020
rect 223757 91082 223823 91085
rect 224861 91082 224927 91085
rect 254577 91082 254643 91085
rect 223757 91080 254643 91082
rect 223757 91024 223762 91080
rect 223818 91024 224866 91080
rect 224922 91024 254582 91080
rect 254638 91024 254643 91080
rect 223757 91022 254643 91024
rect 223757 91019 223823 91022
rect 224861 91019 224927 91022
rect 254577 91019 254643 91022
rect 52361 90946 52427 90949
rect 74257 90946 74323 90949
rect 52361 90944 74323 90946
rect 52361 90888 52366 90944
rect 52422 90888 74262 90944
rect 74318 90888 74323 90944
rect 52361 90886 74323 90888
rect 52361 90883 52427 90886
rect 74257 90883 74323 90886
rect 78949 90946 79015 90949
rect 109125 90946 109191 90949
rect 205081 90946 205147 90949
rect 78949 90944 205147 90946
rect 78949 90888 78954 90944
rect 79010 90888 109130 90944
rect 109186 90888 205086 90944
rect 205142 90888 205147 90944
rect 78949 90886 205147 90888
rect 78949 90883 79015 90886
rect 109125 90883 109191 90886
rect 205081 90883 205147 90886
rect 108389 90402 108455 90405
rect 203609 90402 203675 90405
rect 108389 90400 203675 90402
rect 108389 90344 108394 90400
rect 108450 90344 203614 90400
rect 203670 90344 203675 90400
rect 108389 90342 203675 90344
rect 108389 90339 108455 90342
rect 203609 90339 203675 90342
rect 219893 90402 219959 90405
rect 230473 90402 230539 90405
rect 580257 90402 580323 90405
rect 219893 90400 580323 90402
rect 219893 90344 219898 90400
rect 219954 90344 230478 90400
rect 230534 90344 580262 90400
rect 580318 90344 580323 90400
rect 219893 90342 580323 90344
rect 219893 90339 219959 90342
rect 230473 90339 230539 90342
rect 580257 90339 580323 90342
rect 207381 90266 207447 90269
rect 208301 90266 208367 90269
rect 207381 90264 208367 90266
rect 207381 90208 207386 90264
rect 207442 90208 208306 90264
rect 208362 90208 208367 90264
rect 207381 90206 208367 90208
rect 207381 90203 207447 90206
rect 208301 90203 208367 90206
rect 78029 89858 78095 89861
rect 204437 89858 204503 89861
rect 78029 89856 204503 89858
rect 78029 89800 78034 89856
rect 78090 89800 204442 89856
rect 204498 89800 204503 89856
rect 78029 89798 204503 89800
rect 78029 89795 78138 89798
rect 204437 89795 204503 89798
rect 56501 89722 56567 89725
rect 78078 89722 78138 89795
rect 56501 89720 78138 89722
rect 56501 89664 56506 89720
rect 56562 89664 78138 89720
rect 56501 89662 78138 89664
rect 198365 89722 198431 89725
rect 269205 89722 269271 89725
rect 582373 89722 582439 89725
rect 198365 89720 582439 89722
rect 198365 89664 198370 89720
rect 198426 89664 269210 89720
rect 269266 89664 582378 89720
rect 582434 89664 582439 89720
rect 198365 89662 582439 89664
rect 56501 89659 56567 89662
rect 198365 89659 198431 89662
rect 269205 89659 269271 89662
rect 582373 89659 582439 89662
rect 91277 89586 91343 89589
rect 186221 89586 186287 89589
rect 220077 89586 220143 89589
rect 91277 89584 220143 89586
rect 91277 89528 91282 89584
rect 91338 89528 186226 89584
rect 186282 89528 220082 89584
rect 220138 89528 220143 89584
rect 91277 89526 220143 89528
rect 91277 89523 91343 89526
rect 186221 89523 186287 89526
rect 220077 89523 220143 89526
rect 82077 89450 82143 89453
rect 111793 89450 111859 89453
rect 82077 89448 111859 89450
rect 82077 89392 82082 89448
rect 82138 89392 111798 89448
rect 111854 89392 111859 89448
rect 82077 89390 111859 89392
rect 82077 89387 82143 89390
rect 111793 89387 111859 89390
rect 82997 89314 83063 89317
rect 210325 89314 210391 89317
rect 82997 89312 210391 89314
rect 82997 89256 83002 89312
rect 83058 89256 210330 89312
rect 210386 89256 210391 89312
rect 82997 89254 210391 89256
rect 82997 89251 83063 89254
rect 210325 89251 210391 89254
rect 68870 88164 68876 88228
rect 68940 88226 68946 88228
rect 82261 88226 82327 88229
rect 68940 88224 82327 88226
rect 68940 88168 82266 88224
rect 82322 88168 82327 88224
rect 68940 88166 82327 88168
rect 68940 88164 68946 88166
rect 82261 88163 82327 88166
rect 89253 88226 89319 88229
rect 122097 88226 122163 88229
rect 122649 88226 122715 88229
rect 221917 88226 221983 88229
rect 89253 88224 118802 88226
rect 89253 88168 89258 88224
rect 89314 88168 118802 88224
rect 89253 88166 118802 88168
rect 89253 88163 89319 88166
rect 84101 88090 84167 88093
rect 113265 88090 113331 88093
rect 84101 88088 113331 88090
rect 84101 88032 84106 88088
rect 84162 88032 113270 88088
rect 113326 88032 113331 88088
rect 84101 88030 113331 88032
rect 118742 88090 118802 88166
rect 122097 88224 221983 88226
rect 122097 88168 122102 88224
rect 122158 88168 122654 88224
rect 122710 88168 221922 88224
rect 221978 88168 221983 88224
rect 122097 88166 221983 88168
rect 122097 88163 122163 88166
rect 122649 88163 122715 88166
rect 221917 88163 221983 88166
rect 120165 88090 120231 88093
rect 217685 88090 217751 88093
rect 118742 88088 217751 88090
rect 118742 88032 120170 88088
rect 120226 88032 217690 88088
rect 217746 88032 217751 88088
rect 118742 88030 217751 88032
rect 84101 88027 84167 88030
rect 113265 88027 113331 88030
rect 120165 88027 120231 88030
rect 217685 88027 217751 88030
rect 69657 87546 69723 87549
rect 97349 87546 97415 87549
rect 69657 87544 97415 87546
rect 69657 87488 69662 87544
rect 69718 87488 97354 87544
rect 97410 87488 97415 87544
rect 69657 87486 97415 87488
rect 69657 87483 69723 87486
rect 97349 87483 97415 87486
rect 193806 87484 193812 87548
rect 193876 87546 193882 87548
rect 298093 87546 298159 87549
rect 193876 87544 298159 87546
rect 193876 87488 298098 87544
rect 298154 87488 298159 87544
rect 193876 87486 298159 87488
rect 193876 87484 193882 87486
rect 298093 87483 298159 87486
rect 86125 86866 86191 86869
rect 103605 86866 103671 86869
rect 104709 86866 104775 86869
rect 86125 86864 104775 86866
rect 86125 86808 86130 86864
rect 86186 86808 103610 86864
rect 103666 86808 104714 86864
rect 104770 86808 104775 86864
rect 86125 86806 104775 86808
rect 86125 86803 86191 86806
rect 103605 86803 103671 86806
rect 104709 86803 104775 86806
rect 208393 86866 208459 86869
rect 285765 86866 285831 86869
rect 208393 86864 285831 86866
rect 208393 86808 208398 86864
rect 208454 86808 285770 86864
rect 285826 86808 285831 86864
rect 208393 86806 285831 86808
rect 208393 86803 208459 86806
rect 285765 86803 285831 86806
rect 89805 86730 89871 86733
rect 119337 86730 119403 86733
rect 218237 86730 218303 86733
rect 89805 86728 218303 86730
rect 89805 86672 89810 86728
rect 89866 86672 119342 86728
rect 119398 86672 218242 86728
rect 218298 86672 218303 86728
rect 89805 86670 218303 86672
rect 89805 86667 89871 86670
rect 119337 86667 119403 86670
rect 218237 86667 218303 86670
rect 57237 86594 57303 86597
rect 94681 86594 94747 86597
rect 57237 86592 94747 86594
rect 57237 86536 57242 86592
rect 57298 86536 94686 86592
rect 94742 86536 94747 86592
rect 57237 86534 94747 86536
rect 57237 86531 57303 86534
rect 94681 86531 94747 86534
rect 104709 86594 104775 86597
rect 214005 86594 214071 86597
rect 104709 86592 214071 86594
rect 104709 86536 104714 86592
rect 104770 86536 214010 86592
rect 214066 86536 214071 86592
rect 104709 86534 214071 86536
rect 104709 86531 104775 86534
rect 214005 86531 214071 86534
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect 78397 85506 78463 85509
rect 110413 85506 110479 85509
rect 204989 85506 205055 85509
rect 78397 85504 205055 85506
rect 78397 85448 78402 85504
rect 78458 85448 110418 85504
rect 110474 85448 204994 85504
rect 205050 85448 205055 85504
rect 78397 85446 205055 85448
rect 78397 85443 78463 85446
rect 110413 85443 110479 85446
rect 204989 85443 205055 85446
rect 87229 85370 87295 85373
rect 122833 85370 122899 85373
rect 124029 85370 124095 85373
rect 87229 85368 124095 85370
rect 87229 85312 87234 85368
rect 87290 85312 122838 85368
rect 122894 85312 124034 85368
rect 124090 85312 124095 85368
rect 87229 85310 124095 85312
rect 87229 85307 87295 85310
rect 122833 85307 122899 85310
rect 124029 85307 124095 85310
rect 184289 85370 184355 85373
rect 226374 85370 226380 85372
rect 184289 85368 226380 85370
rect 184289 85312 184294 85368
rect 184350 85312 226380 85368
rect 184289 85310 226380 85312
rect 184289 85307 184355 85310
rect 226374 85308 226380 85310
rect 226444 85308 226450 85372
rect -960 84690 480 84780
rect 3417 84690 3483 84693
rect -960 84688 3483 84690
rect -960 84632 3422 84688
rect 3478 84632 3483 84688
rect -960 84630 3483 84632
rect -960 84540 480 84630
rect 3417 84627 3483 84630
rect 66478 84084 66484 84148
rect 66548 84146 66554 84148
rect 156597 84146 156663 84149
rect 66548 84144 156663 84146
rect 66548 84088 156602 84144
rect 156658 84088 156663 84144
rect 66548 84086 156663 84088
rect 66548 84084 66554 84086
rect 156597 84083 156663 84086
rect 160829 84146 160895 84149
rect 225045 84146 225111 84149
rect 160829 84144 225111 84146
rect 160829 84088 160834 84144
rect 160890 84088 225050 84144
rect 225106 84088 225111 84144
rect 160829 84086 225111 84088
rect 160829 84083 160895 84086
rect 225045 84083 225111 84086
rect 192845 83466 192911 83469
rect 335353 83466 335419 83469
rect 192845 83464 335419 83466
rect 192845 83408 192850 83464
rect 192906 83408 335358 83464
rect 335414 83408 335419 83464
rect 192845 83406 335419 83408
rect 192845 83403 192911 83406
rect 335353 83403 335419 83406
rect 65977 82786 66043 82789
rect 189073 82786 189139 82789
rect 65977 82784 189139 82786
rect 65977 82728 65982 82784
rect 66038 82728 189078 82784
rect 189134 82728 189139 82784
rect 65977 82726 189139 82728
rect 65977 82723 66043 82726
rect 189073 82723 189139 82726
rect 184197 82650 184263 82653
rect 231945 82650 232011 82653
rect 184197 82648 232011 82650
rect 184197 82592 184202 82648
rect 184258 82592 231950 82648
rect 232006 82592 232011 82648
rect 184197 82590 232011 82592
rect 184197 82587 184263 82590
rect 231945 82587 232011 82590
rect 88241 82106 88307 82109
rect 182817 82106 182883 82109
rect 88241 82104 182883 82106
rect 88241 82048 88246 82104
rect 88302 82048 182822 82104
rect 182878 82048 182883 82104
rect 88241 82046 182883 82048
rect 88241 82043 88307 82046
rect 182817 82043 182883 82046
rect 189073 81562 189139 81565
rect 189717 81562 189783 81565
rect 189073 81560 189783 81562
rect 189073 81504 189078 81560
rect 189134 81504 189722 81560
rect 189778 81504 189783 81560
rect 189073 81502 189783 81504
rect 189073 81499 189139 81502
rect 189717 81499 189783 81502
rect 82813 81426 82879 81429
rect 180701 81426 180767 81429
rect 209865 81426 209931 81429
rect 211061 81426 211127 81429
rect 82813 81424 211127 81426
rect 82813 81368 82818 81424
rect 82874 81368 180706 81424
rect 180762 81368 209870 81424
rect 209926 81368 211066 81424
rect 211122 81368 211127 81424
rect 82813 81366 211127 81368
rect 82813 81363 82879 81366
rect 180701 81363 180767 81366
rect 209865 81363 209931 81366
rect 211061 81363 211127 81366
rect 212533 81426 212599 81429
rect 246297 81426 246363 81429
rect 212533 81424 246363 81426
rect 212533 81368 212538 81424
rect 212594 81368 246302 81424
rect 246358 81368 246363 81424
rect 212533 81366 246363 81368
rect 212533 81363 212599 81366
rect 246297 81363 246363 81366
rect 212533 80202 212599 80205
rect 213177 80202 213243 80205
rect 212533 80200 213243 80202
rect 212533 80144 212538 80200
rect 212594 80144 213182 80200
rect 213238 80144 213243 80200
rect 212533 80142 213243 80144
rect 212533 80139 212599 80142
rect 213177 80139 213243 80142
rect 69606 80004 69612 80068
rect 69676 80066 69682 80068
rect 98821 80066 98887 80069
rect 69676 80064 98887 80066
rect 69676 80008 98826 80064
rect 98882 80008 98887 80064
rect 69676 80006 98887 80008
rect 69676 80004 69682 80006
rect 98821 80003 98887 80006
rect 99281 80066 99347 80069
rect 224902 80066 224908 80068
rect 99281 80064 224908 80066
rect 99281 80008 99286 80064
rect 99342 80008 224908 80064
rect 99281 80006 224908 80008
rect 99281 80003 99347 80006
rect 224902 80004 224908 80006
rect 224972 80004 224978 80068
rect 187141 78570 187207 78573
rect 233233 78570 233299 78573
rect 187141 78568 233299 78570
rect 187141 78512 187146 78568
rect 187202 78512 233238 78568
rect 233294 78512 233299 78568
rect 187141 78510 233299 78512
rect 187141 78507 187207 78510
rect 233233 78507 233299 78510
rect 62021 77890 62087 77893
rect 185577 77890 185643 77893
rect 62021 77888 185643 77890
rect 62021 77832 62026 77888
rect 62082 77832 185582 77888
rect 185638 77832 185643 77888
rect 62021 77830 185643 77832
rect 62021 77827 62087 77830
rect 185577 77827 185643 77830
rect 209957 77210 210023 77213
rect 250437 77210 250503 77213
rect 209957 77208 250503 77210
rect 209957 77152 209962 77208
rect 210018 77152 250442 77208
rect 250498 77152 250503 77208
rect 209957 77150 250503 77152
rect 209957 77147 210023 77150
rect 250437 77147 250503 77150
rect 71681 76530 71747 76533
rect 174537 76530 174603 76533
rect 71681 76528 174603 76530
rect 71681 76472 71686 76528
rect 71742 76472 174542 76528
rect 174598 76472 174603 76528
rect 71681 76470 174603 76472
rect 71681 76467 71747 76470
rect 174537 76467 174603 76470
rect 101489 75850 101555 75853
rect 229185 75850 229251 75853
rect 101489 75848 229251 75850
rect 101489 75792 101494 75848
rect 101550 75792 229190 75848
rect 229246 75792 229251 75848
rect 101489 75790 229251 75792
rect 101489 75787 101555 75790
rect 229185 75787 229251 75790
rect 66161 74490 66227 74493
rect 184749 74490 184815 74493
rect 264237 74490 264303 74493
rect 66161 74488 264303 74490
rect 66161 74432 66166 74488
rect 66222 74432 184754 74488
rect 184810 74432 264242 74488
rect 264298 74432 264303 74488
rect 66161 74430 264303 74432
rect 66161 74427 66227 74430
rect 184749 74427 184815 74430
rect 264237 74427 264303 74430
rect 192702 73748 192708 73812
rect 192772 73810 192778 73812
rect 280153 73810 280219 73813
rect 192772 73808 280219 73810
rect 192772 73752 280158 73808
rect 280214 73752 280219 73808
rect 192772 73750 280219 73752
rect 192772 73748 192778 73750
rect 280153 73747 280219 73750
rect 263593 73266 263659 73269
rect 264237 73266 264303 73269
rect 263593 73264 264303 73266
rect 263593 73208 263598 73264
rect 263654 73208 264242 73264
rect 264298 73208 264303 73264
rect 263593 73206 264303 73208
rect 263593 73203 263659 73206
rect 264237 73203 264303 73206
rect 57881 73130 57947 73133
rect 188337 73130 188403 73133
rect 57881 73128 188403 73130
rect 57881 73072 57886 73128
rect 57942 73072 188342 73128
rect 188398 73072 188403 73128
rect 57881 73070 188403 73072
rect 57881 73067 57947 73070
rect 188337 73067 188403 73070
rect 97257 72994 97323 72997
rect 224217 72994 224283 72997
rect 97257 72992 224283 72994
rect 97257 72936 97262 72992
rect 97318 72936 224222 72992
rect 224278 72936 224283 72992
rect 97257 72934 224283 72936
rect 97257 72931 97323 72934
rect 224217 72931 224283 72934
rect 580257 72994 580323 72997
rect 583520 72994 584960 73084
rect 580257 72992 584960 72994
rect 580257 72936 580262 72992
rect 580318 72936 584960 72992
rect 580257 72934 584960 72936
rect 580257 72931 580323 72934
rect 583520 72844 584960 72934
rect 57237 71906 57303 71909
rect 57881 71906 57947 71909
rect 57237 71904 57947 71906
rect 57237 71848 57242 71904
rect 57298 71848 57886 71904
rect 57942 71848 57947 71904
rect 57237 71846 57947 71848
rect 57237 71843 57303 71846
rect 57881 71843 57947 71846
rect 71037 71770 71103 71773
rect 194685 71770 194751 71773
rect 71037 71768 194751 71770
rect -960 71634 480 71724
rect 71037 71712 71042 71768
rect 71098 71712 194690 71768
rect 194746 71712 194751 71768
rect 71037 71710 194751 71712
rect 71037 71707 71103 71710
rect 194685 71707 194751 71710
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 194685 70410 194751 70413
rect 195237 70410 195303 70413
rect 194685 70408 195303 70410
rect 194685 70352 194690 70408
rect 194746 70352 195242 70408
rect 195298 70352 195303 70408
rect 194685 70350 195303 70352
rect 194685 70347 194751 70350
rect 195237 70347 195303 70350
rect 69749 70274 69815 70277
rect 194593 70274 194659 70277
rect 69749 70272 194659 70274
rect 69749 70216 69754 70272
rect 69810 70216 194598 70272
rect 194654 70216 194659 70272
rect 69749 70214 194659 70216
rect 69749 70211 69815 70214
rect 194593 70211 194659 70214
rect 194593 69866 194659 69869
rect 195329 69866 195395 69869
rect 194593 69864 195395 69866
rect 194593 69808 194598 69864
rect 194654 69808 195334 69864
rect 195390 69808 195395 69864
rect 194593 69806 195395 69808
rect 194593 69803 194659 69806
rect 195329 69803 195395 69806
rect 99281 66874 99347 66877
rect 235993 66874 236059 66877
rect 99281 66872 236059 66874
rect 99281 66816 99286 66872
rect 99342 66816 235998 66872
rect 236054 66816 236059 66872
rect 99281 66814 236059 66816
rect 99281 66811 99347 66814
rect 235993 66811 236059 66814
rect 195329 64154 195395 64157
rect 345013 64154 345079 64157
rect 195329 64152 345079 64154
rect 195329 64096 195334 64152
rect 195390 64096 345018 64152
rect 345074 64096 345079 64152
rect 195329 64094 345079 64096
rect 195329 64091 195395 64094
rect 345013 64091 345079 64094
rect 83457 62794 83523 62797
rect 233366 62794 233372 62796
rect 83457 62792 233372 62794
rect 83457 62736 83462 62792
rect 83518 62736 233372 62792
rect 83457 62734 233372 62736
rect 83457 62731 83523 62734
rect 233366 62732 233372 62734
rect 233436 62732 233442 62796
rect 90357 61434 90423 61437
rect 230422 61434 230428 61436
rect 90357 61432 230428 61434
rect 90357 61376 90362 61432
rect 90418 61376 230428 61432
rect 90357 61374 230428 61376
rect 90357 61371 90423 61374
rect 230422 61372 230428 61374
rect 230492 61372 230498 61436
rect 67817 60618 67883 60621
rect 204621 60618 204687 60621
rect 67817 60616 204687 60618
rect 67817 60560 67822 60616
rect 67878 60560 204626 60616
rect 204682 60560 204687 60616
rect 67817 60558 204687 60560
rect 67817 60555 67883 60558
rect 204621 60555 204687 60558
rect 204621 60210 204687 60213
rect 204989 60210 205055 60213
rect 204621 60208 205055 60210
rect 204621 60152 204626 60208
rect 204682 60152 204994 60208
rect 205050 60152 205055 60208
rect 204621 60150 205055 60152
rect 204621 60147 204687 60150
rect 204989 60147 205055 60150
rect 582649 59666 582715 59669
rect 583520 59666 584960 59756
rect 582649 59664 584960 59666
rect 582649 59608 582654 59664
rect 582710 59608 584960 59664
rect 582649 59606 584960 59608
rect 582649 59603 582715 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3509 58578 3575 58581
rect -960 58576 3575 58578
rect -960 58520 3514 58576
rect 3570 58520 3575 58576
rect -960 58518 3575 58520
rect -960 58428 480 58518
rect 3509 58515 3575 58518
rect 196566 58516 196572 58580
rect 196636 58578 196642 58580
rect 262213 58578 262279 58581
rect 196636 58576 262279 58578
rect 196636 58520 262218 58576
rect 262274 58520 262279 58576
rect 196636 58518 262279 58520
rect 196636 58516 196642 58518
rect 262213 58515 262279 58518
rect 95141 55858 95207 55861
rect 234654 55858 234660 55860
rect 95141 55856 234660 55858
rect 95141 55800 95146 55856
rect 95202 55800 234660 55856
rect 95141 55798 234660 55800
rect 95141 55795 95207 55798
rect 234654 55796 234660 55798
rect 234724 55796 234730 55860
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 582833 33146 582899 33149
rect 583520 33146 584960 33236
rect 582833 33144 584960 33146
rect 582833 33088 582838 33144
rect 582894 33088 584960 33144
rect 582833 33086 584960 33088
rect 582833 33083 582899 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 2865 32466 2931 32469
rect -960 32464 2931 32466
rect -960 32408 2870 32464
rect 2926 32408 2931 32464
rect -960 32406 2931 32408
rect -960 32316 480 32406
rect 2865 32403 2931 32406
rect 197118 24108 197124 24172
rect 197188 24170 197194 24172
rect 303613 24170 303679 24173
rect 197188 24168 303679 24170
rect 197188 24112 303618 24168
rect 303674 24112 303679 24168
rect 197188 24110 303679 24112
rect 197188 24108 197194 24110
rect 303613 24107 303679 24110
rect 582557 19818 582623 19821
rect 583520 19818 584960 19908
rect 582557 19816 584960 19818
rect 582557 19760 582562 19816
rect 582618 19760 584960 19816
rect 582557 19758 584960 19760
rect 582557 19755 582623 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 85481 17234 85547 17237
rect 233182 17234 233188 17236
rect 85481 17232 233188 17234
rect 85481 17176 85486 17232
rect 85542 17176 233188 17232
rect 85481 17174 233188 17176
rect 85481 17171 85547 17174
rect 233182 17172 233188 17174
rect 233252 17172 233258 17236
rect 79317 15874 79383 15877
rect 232262 15874 232268 15876
rect 79317 15872 232268 15874
rect 79317 15816 79322 15872
rect 79378 15816 232268 15872
rect 79317 15814 232268 15816
rect 79317 15811 79383 15814
rect 232262 15812 232268 15814
rect 232332 15812 232338 15876
rect 70117 14514 70183 14517
rect 230790 14514 230796 14516
rect 70117 14512 230796 14514
rect 70117 14456 70122 14512
rect 70178 14456 230796 14512
rect 70117 14454 230796 14456
rect 70117 14451 70183 14454
rect 230790 14452 230796 14454
rect 230860 14452 230866 14516
rect 64781 10298 64847 10301
rect 178534 10298 178540 10300
rect 64781 10296 178540 10298
rect 64781 10240 64786 10296
rect 64842 10240 178540 10296
rect 64781 10238 178540 10240
rect 64781 10235 64847 10238
rect 178534 10236 178540 10238
rect 178604 10236 178610 10300
rect 82077 8938 82143 8941
rect 160686 8938 160692 8940
rect 82077 8936 160692 8938
rect 82077 8880 82082 8936
rect 82138 8880 160692 8936
rect 82077 8878 160692 8880
rect 82077 8875 82143 8878
rect 160686 8876 160692 8878
rect 160756 8876 160762 8940
rect 582741 6626 582807 6629
rect 583520 6626 584960 6716
rect 582741 6624 584960 6626
rect -960 6490 480 6580
rect 582741 6568 582746 6624
rect 582802 6568 584960 6624
rect 582741 6566 584960 6568
rect 582741 6563 582807 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 19425 4858 19491 4861
rect 168966 4858 168972 4860
rect 19425 4856 168972 4858
rect 19425 4800 19430 4856
rect 19486 4800 168972 4856
rect 19425 4798 168972 4800
rect 19425 4795 19491 4798
rect 168966 4796 168972 4798
rect 169036 4796 169042 4860
rect 63217 4042 63283 4045
rect 65374 4042 65380 4044
rect 63217 4040 65380 4042
rect 63217 3984 63222 4040
rect 63278 3984 65380 4040
rect 63217 3982 65380 3984
rect 63217 3979 63283 3982
rect 65374 3980 65380 3982
rect 65444 3980 65450 4044
rect 73797 3498 73863 3501
rect 105486 3498 105492 3500
rect 73797 3496 105492 3498
rect 73797 3440 73802 3496
rect 73858 3440 105492 3496
rect 73797 3438 105492 3440
rect 73797 3435 73863 3438
rect 105486 3436 105492 3438
rect 105556 3436 105562 3500
rect 109309 3498 109375 3501
rect 148317 3498 148383 3501
rect 109309 3496 148383 3498
rect 109309 3440 109314 3496
rect 109370 3440 148322 3496
rect 148378 3440 148383 3496
rect 109309 3438 148383 3440
rect 109309 3435 109375 3438
rect 148317 3435 148383 3438
rect 8753 3362 8819 3365
rect 35157 3362 35223 3365
rect 8753 3360 35223 3362
rect 8753 3304 8758 3360
rect 8814 3304 35162 3360
rect 35218 3304 35223 3360
rect 8753 3302 35223 3304
rect 8753 3299 8819 3302
rect 35157 3299 35223 3302
rect 101029 3362 101095 3365
rect 152457 3362 152523 3365
rect 101029 3360 152523 3362
rect 101029 3304 101034 3360
rect 101090 3304 152462 3360
rect 152518 3304 152523 3360
rect 101029 3302 152523 3304
rect 101029 3299 101095 3302
rect 152457 3299 152523 3302
rect 214557 3362 214623 3365
rect 246389 3362 246455 3365
rect 214557 3360 246455 3362
rect 214557 3304 214562 3360
rect 214618 3304 246394 3360
rect 246450 3304 246455 3360
rect 214557 3302 246455 3304
rect 214557 3299 214623 3302
rect 246389 3299 246455 3302
<< via3 >>
rect 268332 702476 268396 702540
rect 260052 699756 260116 699820
rect 74580 621556 74644 621620
rect 125732 590684 125796 590748
rect 76052 584836 76116 584900
rect 74580 582388 74644 582452
rect 75684 580892 75748 580956
rect 70532 580756 70596 580820
rect 79732 580816 79796 580820
rect 79732 580760 79782 580816
rect 79782 580760 79796 580816
rect 79732 580756 79796 580760
rect 83964 580756 84028 580820
rect 88380 580756 88444 580820
rect 91508 580756 91572 580820
rect 104940 571372 105004 571436
rect 94084 567020 94148 567084
rect 110644 559404 110708 559468
rect 100708 549340 100772 549404
rect 69060 548252 69124 548316
rect 96660 547028 96724 547092
rect 67772 542404 67836 542468
rect 69428 542132 69492 542196
rect 96844 541588 96908 541652
rect 76052 539548 76116 539612
rect 111748 534652 111812 534716
rect 96844 531932 96908 531996
rect 79916 530708 79980 530772
rect 93900 530708 93964 530772
rect 96660 530572 96724 530636
rect 73476 524996 73540 525060
rect 91508 524996 91572 525060
rect 77156 523636 77220 523700
rect 102180 522276 102244 522340
rect 107700 479436 107764 479500
rect 100156 476716 100220 476780
rect 72372 473996 72436 474060
rect 81940 471820 82004 471884
rect 83964 471820 84028 471884
rect 106412 468556 106476 468620
rect 69612 468420 69676 468484
rect 88748 468420 88812 468484
rect 75684 462844 75748 462908
rect 93900 462844 93964 462908
rect 79732 456044 79796 456108
rect 80100 456044 80164 456108
rect 114324 450468 114388 450532
rect 67772 449924 67836 449988
rect 67772 442852 67836 442916
rect 70532 442852 70596 442916
rect 71452 441628 71516 441692
rect 115980 440268 116044 440332
rect 109540 439452 109604 439516
rect 88380 438092 88444 438156
rect 78444 437472 78508 437476
rect 78444 437416 78458 437472
rect 78458 437416 78508 437472
rect 78444 437412 78508 437416
rect 71636 436324 71700 436388
rect 90220 436324 90284 436388
rect 72740 436188 72804 436252
rect 83412 436188 83476 436252
rect 95004 436188 95068 436252
rect 69060 436052 69124 436116
rect 78444 436052 78508 436116
rect 93900 436052 93964 436116
rect 103284 436112 103348 436116
rect 103284 436056 103334 436112
rect 103334 436056 103348 436112
rect 103284 436052 103348 436056
rect 105124 436052 105188 436116
rect 73660 435236 73724 435300
rect 92980 434556 93044 434620
rect 80652 434420 80716 434484
rect 74580 434284 74644 434348
rect 75868 434284 75932 434348
rect 94820 434344 94884 434348
rect 94820 434288 94834 434344
rect 94834 434288 94884 434344
rect 94820 434284 94884 434288
rect 96292 434344 96356 434348
rect 96292 434288 96342 434344
rect 96342 434288 96356 434344
rect 96292 434284 96356 434288
rect 108988 434284 109052 434348
rect 92612 434208 92676 434212
rect 92612 434152 92662 434208
rect 92662 434152 92676 434208
rect 92612 434148 92676 434152
rect 96844 434148 96908 434212
rect 96476 434012 96540 434076
rect 109540 434012 109604 434076
rect 112116 434012 112180 434076
rect 82676 433876 82740 433940
rect 97212 433876 97276 433940
rect 75684 433740 75748 433804
rect 86172 433740 86236 433804
rect 91324 433740 91388 433804
rect 98500 433740 98564 433804
rect 108436 433740 108500 433804
rect 69612 433604 69676 433668
rect 77340 433604 77404 433668
rect 78628 433604 78692 433668
rect 83596 433604 83660 433668
rect 84148 433604 84212 433668
rect 85252 433604 85316 433668
rect 85804 433604 85868 433668
rect 87092 433664 87156 433668
rect 87092 433608 87142 433664
rect 87142 433608 87156 433664
rect 87092 433604 87156 433608
rect 87460 433604 87524 433668
rect 89852 433604 89916 433668
rect 91508 433604 91572 433668
rect 98316 433604 98380 433668
rect 99972 433664 100036 433668
rect 99972 433608 99986 433664
rect 99986 433608 100036 433664
rect 99972 433604 100036 433608
rect 100892 433604 100956 433668
rect 102180 433604 102244 433668
rect 104204 433664 104268 433668
rect 104204 433608 104218 433664
rect 104218 433608 104268 433664
rect 104204 433604 104268 433608
rect 105124 433604 105188 433668
rect 106412 433604 106476 433668
rect 110644 433604 110708 433668
rect 111932 433664 111996 433668
rect 111932 433608 111946 433664
rect 111946 433608 111996 433664
rect 111932 433604 111996 433608
rect 112116 432788 112180 432852
rect 64644 425172 64708 425236
rect 66852 422180 66916 422244
rect 66852 420820 66916 420884
rect 114508 417828 114572 417892
rect 66116 415924 66180 415988
rect 66668 409668 66732 409732
rect 67772 409668 67836 409732
rect 114692 408580 114756 408644
rect 114324 399468 114388 399532
rect 68140 394572 68204 394636
rect 85252 390628 85316 390692
rect 103284 390900 103348 390964
rect 106228 390900 106292 390964
rect 72372 390416 72436 390420
rect 72372 390360 72386 390416
rect 72386 390360 72436 390416
rect 72372 390356 72436 390360
rect 73476 390356 73540 390420
rect 77156 390416 77220 390420
rect 77156 390360 77206 390416
rect 77206 390360 77220 390416
rect 77156 390356 77220 390360
rect 79916 390356 79980 390420
rect 81940 390416 82004 390420
rect 81940 390360 81990 390416
rect 81990 390360 82004 390416
rect 81940 390356 82004 390360
rect 107700 390552 107764 390556
rect 107700 390496 107750 390552
rect 107750 390496 107764 390552
rect 107700 390492 107764 390496
rect 111748 390416 111812 390420
rect 111748 390360 111762 390416
rect 111762 390360 111812 390416
rect 111748 390356 111812 390360
rect 108620 390220 108684 390284
rect 96292 389540 96356 389604
rect 71452 388996 71516 389060
rect 78812 389056 78876 389060
rect 78812 389000 78862 389056
rect 78862 389000 78876 389056
rect 78812 388996 78876 389000
rect 80100 389056 80164 389060
rect 80100 389000 80114 389056
rect 80114 389000 80164 389056
rect 80100 388996 80164 389000
rect 88748 388996 88812 389060
rect 100156 388996 100220 389060
rect 100708 389056 100772 389060
rect 100708 389000 100758 389056
rect 100758 389000 100772 389056
rect 100708 388996 100772 389000
rect 104940 388996 105004 389060
rect 125732 388996 125796 389060
rect 57100 388860 57164 388924
rect 78444 387908 78508 387972
rect 70900 387772 70964 387836
rect 91508 387772 91572 387836
rect 73476 387636 73540 387700
rect 73476 387500 73540 387564
rect 102180 386956 102244 387020
rect 72924 385732 72988 385796
rect 97212 385596 97276 385660
rect 78812 384236 78876 384300
rect 105124 384236 105188 384300
rect 108252 384236 108316 384300
rect 85804 383692 85868 383756
rect 68140 383556 68204 383620
rect 95004 382196 95068 382260
rect 95188 380972 95252 381036
rect 100708 380972 100772 381036
rect 78628 380156 78692 380220
rect 96844 380156 96908 380220
rect 87460 378660 87524 378724
rect 91324 375940 91388 376004
rect 91508 375940 91572 376004
rect 108988 375940 109052 376004
rect 106412 374580 106476 374644
rect 100892 373220 100956 373284
rect 83964 365604 84028 365668
rect 74580 364380 74644 364444
rect 104204 353908 104268 353972
rect 88012 351868 88076 351932
rect 82860 339492 82924 339556
rect 83596 339552 83660 339556
rect 83596 339496 83610 339552
rect 83610 339496 83660 339552
rect 83596 339492 83660 339496
rect 237972 335412 238036 335476
rect 98132 332556 98196 332620
rect 98500 332556 98564 332620
rect 92612 330380 92676 330444
rect 242020 329836 242084 329900
rect 111932 327660 111996 327724
rect 82860 326980 82924 327044
rect 99972 326300 100036 326364
rect 86172 323580 86236 323644
rect 86724 322900 86788 322964
rect 75684 321540 75748 321604
rect 90956 321404 91020 321468
rect 89852 320724 89916 320788
rect 210372 320180 210436 320244
rect 98316 319500 98380 319564
rect 115980 319364 116044 319428
rect 262260 319364 262324 319428
rect 94820 318820 94884 318884
rect 77340 318684 77404 318748
rect 87092 318276 87156 318340
rect 114692 318276 114756 318340
rect 258396 318276 258460 318340
rect 253060 318140 253124 318204
rect 260052 318004 260116 318068
rect 75868 317460 75932 317524
rect 98132 316644 98196 316708
rect 258396 314876 258460 314940
rect 66484 312156 66548 312220
rect 66668 312020 66732 312084
rect 201540 310796 201604 310860
rect 201540 308212 201604 308276
rect 254532 306988 254596 307052
rect 197308 306444 197372 306508
rect 80652 304132 80716 304196
rect 239260 303860 239324 303924
rect 83412 303588 83476 303652
rect 213684 303588 213748 303652
rect 219940 303588 220004 303652
rect 237972 303588 238036 303652
rect 240732 303648 240796 303652
rect 240732 303592 240746 303648
rect 240746 303592 240796 303648
rect 240732 303588 240796 303592
rect 242020 303588 242084 303652
rect 193444 302228 193508 302292
rect 193260 301820 193324 301884
rect 254164 301684 254228 301748
rect 224172 301276 224236 301340
rect 233188 301276 233252 301340
rect 234660 301276 234724 301340
rect 236500 301276 236564 301340
rect 238156 301276 238220 301340
rect 212396 301140 212460 301204
rect 215892 301004 215956 301068
rect 218652 301004 218716 301068
rect 194548 300868 194612 300932
rect 198780 300868 198844 300932
rect 204852 300868 204916 300932
rect 205772 300868 205836 300932
rect 207060 300928 207124 300932
rect 207060 300872 207110 300928
rect 207110 300872 207124 300928
rect 207060 300868 207124 300872
rect 214420 300868 214484 300932
rect 217180 300868 217244 300932
rect 219204 300868 219268 300932
rect 220860 300868 220924 300932
rect 222332 300928 222396 300932
rect 222332 300872 222382 300928
rect 222382 300872 222396 300928
rect 222332 300868 222396 300872
rect 224356 300868 224420 300932
rect 226012 300928 226076 300932
rect 226012 300872 226026 300928
rect 226026 300872 226076 300928
rect 226012 300868 226076 300872
rect 226564 300928 226628 300932
rect 226564 300872 226578 300928
rect 226578 300872 226628 300928
rect 226564 300868 226628 300872
rect 226748 300868 226812 300932
rect 229692 300868 229756 300932
rect 230428 300868 230492 300932
rect 230796 300868 230860 300932
rect 232084 300928 232148 300932
rect 232084 300872 232098 300928
rect 232098 300872 232148 300928
rect 232084 300868 232148 300872
rect 232268 300868 232332 300932
rect 233372 300928 233436 300932
rect 233372 300872 233386 300928
rect 233386 300872 233436 300928
rect 233372 300868 233436 300872
rect 234844 300868 234908 300932
rect 236684 300928 236748 300932
rect 236684 300872 236698 300928
rect 236698 300872 236748 300928
rect 236684 300868 236748 300872
rect 238708 300868 238772 300932
rect 240916 300868 240980 300932
rect 241652 300868 241716 300932
rect 242940 300868 243004 300932
rect 244412 300868 244476 300932
rect 245700 300868 245764 300932
rect 247724 300928 247788 300932
rect 247724 300872 247774 300928
rect 247774 300872 247788 300928
rect 247724 300868 247788 300872
rect 248460 300928 248524 300932
rect 248460 300872 248510 300928
rect 248510 300872 248524 300928
rect 248460 300868 248524 300872
rect 251220 300868 251284 300932
rect 252508 300928 252572 300932
rect 252508 300872 252522 300928
rect 252522 300872 252572 300928
rect 252508 300868 252572 300872
rect 86172 300732 86236 300796
rect 196572 300732 196636 300796
rect 208532 300732 208596 300796
rect 197308 300596 197372 300660
rect 210372 300596 210436 300660
rect 255452 300324 255516 300388
rect 256740 300188 256804 300252
rect 255268 299508 255332 299572
rect 256556 299372 256620 299436
rect 254532 298964 254596 299028
rect 193444 298828 193508 298892
rect 72740 298692 72804 298756
rect 255452 298692 255516 298756
rect 255268 298556 255332 298620
rect 254532 298148 254596 298212
rect 193260 296652 193324 296716
rect 193076 296516 193140 296580
rect 191604 295156 191668 295220
rect 94452 294612 94516 294676
rect 101260 294612 101324 294676
rect 256556 294476 256620 294540
rect 254164 294204 254228 294268
rect 92980 293312 93044 293316
rect 92980 293256 93030 293312
rect 93030 293256 93044 293312
rect 92980 293252 93044 293256
rect 83412 293116 83476 293180
rect 253612 292708 253676 292772
rect 70164 292572 70228 292636
rect 100708 291892 100772 291956
rect 256740 290668 256804 290732
rect 82676 289096 82740 289100
rect 82676 289040 82726 289096
rect 82726 289040 82740 289096
rect 82676 289036 82740 289040
rect 90220 288356 90284 288420
rect 97948 287268 98012 287332
rect 193996 286452 194060 286516
rect 71636 286044 71700 286108
rect 50844 285772 50908 285836
rect 69612 285636 69676 285700
rect 82676 285636 82740 285700
rect 88748 285636 88812 285700
rect 97948 284820 98012 284884
rect 72372 284140 72436 284204
rect 91324 284140 91388 284204
rect 95188 283732 95252 283796
rect 96476 283732 96540 283796
rect 68876 283596 68940 283660
rect 69980 283596 70044 283660
rect 84700 283596 84764 283660
rect 73108 283520 73172 283524
rect 73108 283464 73158 283520
rect 73158 283464 73172 283520
rect 73108 283460 73172 283464
rect 89852 283520 89916 283524
rect 89852 283464 89866 283520
rect 89866 283464 89916 283520
rect 89852 283460 89916 283464
rect 92612 283520 92676 283524
rect 92612 283464 92626 283520
rect 92626 283464 92676 283520
rect 92612 283460 92676 283464
rect 75684 283248 75748 283252
rect 75684 283192 75734 283248
rect 75734 283192 75748 283248
rect 75684 283188 75748 283192
rect 70348 282916 70412 282980
rect 83964 282916 84028 282980
rect 87828 282976 87892 282980
rect 87828 282920 87878 282976
rect 87878 282920 87892 282976
rect 87828 282916 87892 282920
rect 88748 282916 88812 282980
rect 98868 282916 98932 282980
rect 100708 282704 100772 282708
rect 100708 282648 100758 282704
rect 100758 282648 100772 282704
rect 100708 282644 100772 282648
rect 101260 278564 101324 278628
rect 66300 277612 66364 277676
rect 98868 277340 98932 277404
rect 66300 274756 66364 274820
rect 184060 274620 184124 274684
rect 114508 271084 114572 271148
rect 64644 269724 64708 269788
rect 108252 268500 108316 268564
rect 259500 267412 259564 267476
rect 110644 267004 110708 267068
rect 108252 266324 108316 266388
rect 268332 265372 268396 265436
rect 258396 265236 258460 265300
rect 65748 265160 65812 265164
rect 65748 265104 65762 265160
rect 65762 265104 65812 265160
rect 65748 265100 65812 265104
rect 110644 264964 110708 265028
rect 160692 263604 160756 263668
rect 108436 262788 108500 262852
rect 255452 261896 255516 261900
rect 255452 261840 255502 261896
rect 255502 261840 255516 261896
rect 255452 261836 255516 261840
rect 66116 261700 66180 261764
rect 108252 260748 108316 260812
rect 255268 260748 255332 260812
rect 256740 260476 256804 260540
rect 262260 259796 262324 259860
rect 64644 258708 64708 258772
rect 111012 258708 111076 258772
rect 263548 258572 263612 258636
rect 178540 258164 178604 258228
rect 262260 258164 262324 258228
rect 259500 257348 259564 257412
rect 267780 257212 267844 257276
rect 99972 256668 100036 256732
rect 98132 255308 98196 255372
rect 269068 255580 269132 255644
rect 258396 254764 258460 254828
rect 108252 254492 108316 254556
rect 266308 253948 266372 254012
rect 273300 253948 273364 254012
rect 66668 253812 66732 253876
rect 254716 253404 254780 253468
rect 188292 253132 188356 253196
rect 259684 248372 259748 248436
rect 61884 248296 61948 248300
rect 61884 248240 61934 248296
rect 61934 248240 61948 248296
rect 61884 248236 61948 248240
rect 193260 247556 193324 247620
rect 258396 247012 258460 247076
rect 168972 244292 169036 244356
rect 259684 244156 259748 244220
rect 252876 243612 252940 243676
rect 57100 242932 57164 242996
rect 57836 242932 57900 242996
rect 193260 242796 193324 242860
rect 99972 242524 100036 242588
rect 192892 242116 192956 242180
rect 70164 241708 70228 241772
rect 70900 241768 70964 241772
rect 70900 241712 70950 241768
rect 70950 241712 70964 241768
rect 70900 241708 70964 241712
rect 72372 241768 72436 241772
rect 72372 241712 72386 241768
rect 72386 241712 72436 241768
rect 72372 241708 72436 241712
rect 73476 241708 73540 241772
rect 83412 241768 83476 241772
rect 83412 241712 83426 241768
rect 83426 241712 83476 241768
rect 83412 241708 83476 241712
rect 84700 241708 84764 241772
rect 86172 241708 86236 241772
rect 86724 241768 86788 241772
rect 86724 241712 86738 241768
rect 86738 241712 86788 241768
rect 86724 241708 86788 241712
rect 88012 241768 88076 241772
rect 88012 241712 88062 241768
rect 88062 241712 88076 241768
rect 88012 241708 88076 241712
rect 69980 241632 70044 241636
rect 69980 241576 70030 241632
rect 70030 241576 70044 241632
rect 69980 241572 70044 241576
rect 72924 241572 72988 241636
rect 91324 241572 91388 241636
rect 57836 241300 57900 241364
rect 83964 241300 84028 241364
rect 104940 241436 105004 241500
rect 193076 241436 193140 241500
rect 111012 241300 111076 241364
rect 192892 240892 192956 240956
rect 258396 240756 258460 240820
rect 201540 240212 201604 240276
rect 84700 240076 84764 240140
rect 91508 240076 91572 240140
rect 95004 240076 95068 240140
rect 97764 240076 97828 240140
rect 215340 240136 215404 240140
rect 215340 240080 215390 240136
rect 215390 240080 215404 240136
rect 215340 240076 215404 240080
rect 72556 239940 72620 240004
rect 234844 240076 234908 240140
rect 236684 240076 236748 240140
rect 254716 240076 254780 240140
rect 215340 239804 215404 239868
rect 90956 239668 91020 239732
rect 256740 239532 256804 239596
rect 252508 239396 252572 239460
rect 238708 238716 238772 238780
rect 259684 238716 259748 238780
rect 93716 238172 93780 238236
rect 242020 238036 242084 238100
rect 262260 238036 262324 238100
rect 64644 237900 64708 237964
rect 198780 237220 198844 237284
rect 95188 236948 95252 237012
rect 210372 235860 210436 235924
rect 92612 235724 92676 235788
rect 269068 235860 269132 235924
rect 266308 235180 266372 235244
rect 125732 234500 125796 234564
rect 228220 234364 228284 234428
rect 267780 234364 267844 234428
rect 209820 233140 209884 233204
rect 195836 231100 195900 231164
rect 254532 231100 254596 231164
rect 68876 230556 68940 230620
rect 208716 227700 208780 227764
rect 223620 227020 223684 227084
rect 220860 226884 220924 226948
rect 224356 226476 224420 226540
rect 65932 226340 65996 226404
rect 259500 226204 259564 226268
rect 273300 226068 273364 226132
rect 201540 223484 201604 223548
rect 224172 222804 224236 222868
rect 108252 221580 108316 221644
rect 255452 221444 255516 221508
rect 263548 220764 263612 220828
rect 217180 220084 217244 220148
rect 226564 218588 226628 218652
rect 226748 217228 226812 217292
rect 61884 216744 61948 216748
rect 61884 216688 61934 216744
rect 61934 216688 61948 216744
rect 61884 216684 61948 216688
rect 215892 216004 215956 216068
rect 72924 215868 72988 215932
rect 238156 214508 238220 214572
rect 248460 213420 248524 213484
rect 184796 213284 184860 213348
rect 255268 213284 255332 213348
rect 236500 213148 236564 213212
rect 184796 212604 184860 212668
rect 188292 212468 188356 212532
rect 222332 211788 222396 211852
rect 188844 211108 188908 211172
rect 219940 210292 220004 210356
rect 71636 208388 71700 208452
rect 190316 208388 190380 208452
rect 97212 207028 97276 207092
rect 224908 207572 224972 207636
rect 226012 207028 226076 207092
rect 207060 206212 207124 206276
rect 245700 206212 245764 206276
rect 203196 205668 203260 205732
rect 204852 204852 204916 204916
rect 68876 203492 68940 203556
rect 82860 203492 82924 203556
rect 214420 203492 214484 203556
rect 203196 202812 203260 202876
rect 196572 202132 196636 202196
rect 205772 199276 205836 199340
rect 105492 196692 105556 196756
rect 232084 196692 232148 196756
rect 194548 196556 194612 196620
rect 204852 193972 204916 194036
rect 251220 193972 251284 194036
rect 208532 193836 208596 193900
rect 201356 186900 201420 186964
rect 240916 186900 240980 186964
rect 65380 184180 65444 184244
rect 229692 184180 229756 184244
rect 247724 181324 247788 181388
rect 218652 178604 218716 178668
rect 87828 177244 87892 177308
rect 87828 176700 87892 176764
rect 207060 173844 207124 173908
rect 239260 173164 239324 173228
rect 241652 171668 241716 171732
rect 252508 166288 252572 166292
rect 252508 166232 252558 166288
rect 252558 166232 252572 166288
rect 252508 166228 252572 166232
rect 69612 164324 69676 164388
rect 187556 164324 187620 164388
rect 227668 164188 227732 164252
rect 227668 162828 227732 162892
rect 212396 160652 212460 160716
rect 89852 156572 89916 156636
rect 213684 155212 213748 155276
rect 226380 154668 226444 154732
rect 228220 154532 228284 154596
rect 50844 153036 50908 153100
rect 213684 148412 213748 148476
rect 242940 148276 243004 148340
rect 66668 147868 66732 147932
rect 192708 147052 192772 147116
rect 244412 147052 244476 147116
rect 219388 145692 219452 145756
rect 100708 145556 100772 145620
rect 65748 144740 65812 144804
rect 184060 144060 184124 144124
rect 88748 143652 88812 143716
rect 198780 143712 198844 143716
rect 198780 143656 198830 143712
rect 198830 143656 198844 143712
rect 198780 143652 198844 143656
rect 196572 142292 196636 142356
rect 90956 142156 91020 142220
rect 197124 142156 197188 142220
rect 200620 142156 200684 142220
rect 224356 142020 224420 142084
rect 70348 141400 70412 141404
rect 70348 141344 70362 141400
rect 70362 141344 70412 141400
rect 70348 141340 70412 141344
rect 198780 141068 198844 141132
rect 73108 140856 73172 140860
rect 73108 140800 73122 140856
rect 73122 140800 73172 140856
rect 73108 140796 73172 140800
rect 193260 139572 193324 139636
rect 227668 139028 227732 139092
rect 69428 138076 69492 138140
rect 70348 137940 70412 138004
rect 68140 136852 68204 136916
rect 94820 136852 94884 136916
rect 224356 136580 224420 136644
rect 226932 136580 226996 136644
rect 227852 136580 227916 136644
rect 90956 135220 91020 135284
rect 95740 135220 95804 135284
rect 94820 133724 94884 133788
rect 187556 131140 187620 131204
rect 69428 131004 69492 131068
rect 226380 130052 226444 130116
rect 191604 129296 191668 129300
rect 191604 129240 191654 129296
rect 191654 129240 191668 129296
rect 191604 129236 191668 129240
rect 68140 126788 68204 126852
rect 193260 125700 193324 125764
rect 69244 125564 69308 125628
rect 193812 125564 193876 125628
rect 97396 124204 97460 124268
rect 192340 124204 192404 124268
rect 226932 121076 226996 121140
rect 192708 120260 192772 120324
rect 95740 118492 95804 118556
rect 192156 118628 192220 118692
rect 192156 117268 192220 117332
rect 192708 117268 192772 117332
rect 224356 114412 224420 114476
rect 237972 113052 238036 113116
rect 237972 111828 238036 111892
rect 240732 111888 240796 111892
rect 240732 111832 240746 111888
rect 240746 111832 240796 111888
rect 240732 111828 240796 111832
rect 66484 109380 66548 109444
rect 186820 109108 186884 109172
rect 97948 108836 98012 108900
rect 66668 103940 66732 104004
rect 69428 99860 69492 99924
rect 225092 98228 225156 98292
rect 184796 96596 184860 96660
rect 226380 97140 226444 97204
rect 66852 95780 66916 95844
rect 188844 95236 188908 95300
rect 226564 95296 226628 95300
rect 226564 95240 226614 95296
rect 226614 95240 226628 95296
rect 226564 95236 226628 95240
rect 66852 94964 66916 95028
rect 224356 94284 224420 94348
rect 97212 92788 97276 92852
rect 72924 92712 72988 92716
rect 72924 92656 72974 92712
rect 72974 92656 72988 92712
rect 72924 92652 72988 92656
rect 93716 92652 93780 92716
rect 215340 93332 215404 93396
rect 224908 93332 224972 93396
rect 201356 92984 201420 92988
rect 201356 92928 201406 92984
rect 201406 92928 201420 92984
rect 201356 92924 201420 92928
rect 193996 92788 194060 92852
rect 195836 92788 195900 92852
rect 200620 92788 200684 92852
rect 201540 92848 201604 92852
rect 201540 92792 201590 92848
rect 201590 92792 201604 92848
rect 201540 92788 201604 92792
rect 207060 92848 207124 92852
rect 207060 92792 207110 92848
rect 207110 92792 207124 92848
rect 207060 92788 207124 92792
rect 208716 92848 208780 92852
rect 208716 92792 208766 92848
rect 208766 92792 208780 92848
rect 208716 92788 208780 92792
rect 209820 92788 209884 92852
rect 213684 92848 213748 92852
rect 213684 92792 213698 92848
rect 213698 92792 213748 92848
rect 213684 92788 213748 92792
rect 204852 92652 204916 92716
rect 91692 92380 91756 92444
rect 203196 92380 203260 92444
rect 226564 92380 226628 92444
rect 186820 92244 186884 92308
rect 97396 92108 97460 92172
rect 224356 92108 224420 92172
rect 190316 91836 190380 91900
rect 192340 91156 192404 91220
rect 71636 91020 71700 91084
rect 100708 91080 100772 91084
rect 100708 91024 100758 91080
rect 100758 91024 100772 91080
rect 100708 91020 100772 91024
rect 68876 88164 68940 88228
rect 193812 87484 193876 87548
rect 226380 85308 226444 85372
rect 66484 84084 66548 84148
rect 69612 80004 69676 80068
rect 224908 80004 224972 80068
rect 192708 73748 192772 73812
rect 233372 62732 233436 62796
rect 230428 61372 230492 61436
rect 196572 58516 196636 58580
rect 234660 55796 234724 55860
rect 197124 24108 197188 24172
rect 233188 17172 233252 17236
rect 232268 15812 232332 15876
rect 230796 14452 230860 14516
rect 178540 10236 178604 10300
rect 160692 8876 160756 8940
rect 168972 4796 169036 4860
rect 65380 3980 65444 4044
rect 105492 3436 105556 3500
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 529174 60134 564618
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 59514 493174 60134 528618
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59514 457174 60134 492618
rect 59514 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 60134 457174
rect 59514 456854 60134 456938
rect 59514 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 60134 456854
rect 59514 421174 60134 456618
rect 59514 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 60134 421174
rect 59514 420854 60134 420938
rect 59514 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 60134 420854
rect 57099 388924 57165 388925
rect 57099 388860 57100 388924
rect 57164 388860 57165 388924
rect 57099 388859 57165 388860
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 50843 285836 50909 285837
rect 50843 285772 50844 285836
rect 50908 285772 50909 285836
rect 50843 285771 50909 285772
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 50846 153101 50906 285771
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 57102 242997 57162 388859
rect 59514 385174 60134 420618
rect 59514 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 60134 385174
rect 59514 384854 60134 384938
rect 59514 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 60134 384854
rect 59514 349174 60134 384618
rect 59514 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 60134 349174
rect 59514 348854 60134 348938
rect 59514 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 60134 348854
rect 59514 313174 60134 348618
rect 59514 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 60134 313174
rect 59514 312854 60134 312938
rect 59514 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 60134 312854
rect 59514 277174 60134 312618
rect 59514 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 60134 277174
rect 59514 276854 60134 276938
rect 59514 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 60134 276854
rect 57099 242996 57165 242997
rect 57099 242932 57100 242996
rect 57164 242932 57165 242996
rect 57099 242931 57165 242932
rect 57835 242996 57901 242997
rect 57835 242932 57836 242996
rect 57900 242932 57901 242996
rect 57835 242931 57901 242932
rect 57838 241365 57898 242931
rect 57835 241364 57901 241365
rect 57835 241300 57836 241364
rect 57900 241300 57901 241364
rect 57835 241299 57901 241300
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 50843 153100 50909 153101
rect 50843 153036 50844 153100
rect 50908 153036 50909 153100
rect 50843 153035 50909 153036
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 241174 60134 276618
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 583166 67574 608058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 74579 621620 74645 621621
rect 74579 621556 74580 621620
rect 74644 621556 74645 621620
rect 74579 621555 74645 621556
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 583166 74414 614898
rect 74582 582453 74642 621555
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 76051 584900 76117 584901
rect 76051 584836 76052 584900
rect 76116 584836 76117 584900
rect 76051 584835 76117 584836
rect 74579 582452 74645 582453
rect 74579 582388 74580 582452
rect 74644 582388 74645 582452
rect 74579 582387 74645 582388
rect 75683 580956 75749 580957
rect 75683 580892 75684 580956
rect 75748 580892 75749 580956
rect 75683 580891 75749 580892
rect 70531 580820 70597 580821
rect 70531 580756 70532 580820
rect 70596 580756 70597 580820
rect 70531 580755 70597 580756
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 532894 63854 568338
rect 69059 548316 69125 548317
rect 69059 548252 69060 548316
rect 69124 548252 69125 548316
rect 69059 548251 69125 548252
rect 67771 542468 67837 542469
rect 67771 542404 67772 542468
rect 67836 542404 67837 542468
rect 67771 542403 67837 542404
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 63234 460894 63854 496338
rect 63234 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 63854 460894
rect 63234 460574 63854 460658
rect 63234 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 63854 460574
rect 63234 424894 63854 460338
rect 66954 536614 67574 537166
rect 66954 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 67574 536614
rect 66954 536294 67574 536378
rect 66954 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 67574 536294
rect 66954 500614 67574 536058
rect 66954 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 67574 500614
rect 66954 500294 67574 500378
rect 66954 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 67574 500294
rect 66954 464614 67574 500058
rect 66954 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 67574 464614
rect 66954 464294 67574 464378
rect 66954 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 67574 464294
rect 66954 436356 67574 464058
rect 67774 449989 67834 542403
rect 67771 449988 67837 449989
rect 67771 449924 67772 449988
rect 67836 449924 67837 449988
rect 67771 449923 67837 449924
rect 67771 442916 67837 442917
rect 67771 442852 67772 442916
rect 67836 442852 67837 442916
rect 67771 442851 67837 442852
rect 64643 425236 64709 425237
rect 64643 425172 64644 425236
rect 64708 425172 64709 425236
rect 64643 425171 64709 425172
rect 63234 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 63854 424894
rect 63234 424574 63854 424658
rect 63234 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 63854 424574
rect 63234 388894 63854 424338
rect 63234 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 63854 388894
rect 63234 388574 63854 388658
rect 63234 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 63854 388574
rect 63234 352894 63854 388338
rect 63234 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 63854 352894
rect 63234 352574 63854 352658
rect 63234 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 63854 352574
rect 63234 316894 63854 352338
rect 63234 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 63854 316894
rect 63234 316574 63854 316658
rect 63234 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 63854 316574
rect 63234 280894 63854 316338
rect 63234 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 63854 280894
rect 63234 280574 63854 280658
rect 63234 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 63854 280574
rect 61883 248300 61949 248301
rect 61883 248236 61884 248300
rect 61948 248236 61949 248300
rect 61883 248235 61949 248236
rect 59514 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 60134 241174
rect 59514 240854 60134 240938
rect 59514 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 60134 240854
rect 59514 205174 60134 240618
rect 61886 216749 61946 248235
rect 63234 244894 63854 280338
rect 64646 269789 64706 425171
rect 66851 422244 66917 422245
rect 66851 422180 66852 422244
rect 66916 422180 66917 422244
rect 66851 422179 66917 422180
rect 66854 420885 66914 422179
rect 66851 420884 66917 420885
rect 66851 420820 66852 420884
rect 66916 420820 66917 420884
rect 66851 420819 66917 420820
rect 66115 415988 66181 415989
rect 66115 415924 66116 415988
rect 66180 415924 66181 415988
rect 66115 415923 66181 415924
rect 64643 269788 64709 269789
rect 64643 269724 64644 269788
rect 64708 269724 64709 269788
rect 64643 269723 64709 269724
rect 65747 265164 65813 265165
rect 65747 265100 65748 265164
rect 65812 265100 65813 265164
rect 65747 265099 65813 265100
rect 64643 258772 64709 258773
rect 64643 258708 64644 258772
rect 64708 258708 64709 258772
rect 64643 258707 64709 258708
rect 63234 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 63854 244894
rect 63234 244574 63854 244658
rect 63234 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 63854 244574
rect 61883 216748 61949 216749
rect 61883 216684 61884 216748
rect 61948 216684 61949 216748
rect 61883 216683 61949 216684
rect 59514 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 60134 205174
rect 59514 204854 60134 204938
rect 59514 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 60134 204854
rect 59514 169174 60134 204618
rect 59514 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 60134 169174
rect 59514 168854 60134 168938
rect 59514 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 60134 168854
rect 59514 133174 60134 168618
rect 59514 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 60134 133174
rect 59514 132854 60134 132938
rect 59514 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 60134 132854
rect 59514 97174 60134 132618
rect 59514 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 60134 97174
rect 59514 96854 60134 96938
rect 59514 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 60134 96854
rect 59514 61174 60134 96618
rect 59514 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 60134 61174
rect 59514 60854 60134 60938
rect 59514 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 60134 60854
rect 59514 25174 60134 60618
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 208894 63854 244338
rect 64646 237965 64706 258707
rect 64643 237964 64709 237965
rect 64643 237900 64644 237964
rect 64708 237900 64709 237964
rect 64643 237899 64709 237900
rect 63234 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 63854 208894
rect 63234 208574 63854 208658
rect 63234 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 63854 208574
rect 63234 172894 63854 208338
rect 65379 184244 65445 184245
rect 65379 184180 65380 184244
rect 65444 184180 65445 184244
rect 65379 184179 65445 184180
rect 63234 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 63854 172894
rect 63234 172574 63854 172658
rect 63234 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 63854 172574
rect 63234 136894 63854 172338
rect 63234 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 63854 136894
rect 63234 136574 63854 136658
rect 63234 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 63854 136574
rect 63234 100894 63854 136338
rect 63234 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 63854 100894
rect 63234 100574 63854 100658
rect 63234 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 63854 100574
rect 63234 64894 63854 100338
rect 63234 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 63854 64894
rect 63234 64574 63854 64658
rect 63234 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 63854 64574
rect 63234 28894 63854 64338
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 65382 4045 65442 184179
rect 65750 144805 65810 265099
rect 66118 261765 66178 415923
rect 67774 409733 67834 442851
rect 69062 436117 69122 548251
rect 69427 542196 69493 542197
rect 69427 542132 69428 542196
rect 69492 542132 69493 542196
rect 69427 542131 69493 542132
rect 69430 538230 69490 542131
rect 69430 538170 69674 538230
rect 69614 468485 69674 538170
rect 69611 468484 69677 468485
rect 69611 468420 69612 468484
rect 69676 468420 69677 468484
rect 69611 468419 69677 468420
rect 70534 442917 70594 580755
rect 73679 543454 73999 543486
rect 73679 543218 73721 543454
rect 73957 543218 73999 543454
rect 73679 543134 73999 543218
rect 73679 542898 73721 543134
rect 73957 542898 73999 543134
rect 73679 542866 73999 542898
rect 73475 525060 73541 525061
rect 73475 524996 73476 525060
rect 73540 524996 73541 525060
rect 73475 524995 73541 524996
rect 72371 474060 72437 474061
rect 72371 473996 72372 474060
rect 72436 473996 72437 474060
rect 72371 473995 72437 473996
rect 70531 442916 70597 442917
rect 70531 442852 70532 442916
rect 70596 442852 70597 442916
rect 70531 442851 70597 442852
rect 71451 441692 71517 441693
rect 71451 441628 71452 441692
rect 71516 441628 71517 441692
rect 71451 441627 71517 441628
rect 69059 436116 69125 436117
rect 69059 436052 69060 436116
rect 69124 436052 69125 436116
rect 69059 436051 69125 436052
rect 69611 433668 69677 433669
rect 69611 433604 69612 433668
rect 69676 433604 69677 433668
rect 69611 433603 69677 433604
rect 66667 409732 66733 409733
rect 66667 409668 66668 409732
rect 66732 409668 66733 409732
rect 66667 409667 66733 409668
rect 67771 409732 67837 409733
rect 67771 409668 67772 409732
rect 67836 409668 67837 409732
rect 67771 409667 67837 409668
rect 66483 312220 66549 312221
rect 66483 312156 66484 312220
rect 66548 312156 66549 312220
rect 66483 312155 66549 312156
rect 66486 306390 66546 312155
rect 66670 312085 66730 409667
rect 68139 394636 68205 394637
rect 68139 394572 68140 394636
rect 68204 394572 68205 394636
rect 68139 394571 68205 394572
rect 66954 356614 67574 388356
rect 68142 383621 68202 394571
rect 68139 383620 68205 383621
rect 68139 383556 68140 383620
rect 68204 383556 68205 383620
rect 68139 383555 68205 383556
rect 66954 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 67574 356614
rect 66954 356294 67574 356378
rect 66954 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 67574 356294
rect 66954 320614 67574 356058
rect 66954 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 67574 320614
rect 66954 320294 67574 320378
rect 66954 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 67574 320294
rect 66667 312084 66733 312085
rect 66667 312020 66668 312084
rect 66732 312020 66733 312084
rect 66667 312019 66733 312020
rect 66486 306330 66730 306390
rect 66299 277676 66365 277677
rect 66299 277612 66300 277676
rect 66364 277612 66365 277676
rect 66299 277611 66365 277612
rect 66302 274821 66362 277611
rect 66299 274820 66365 274821
rect 66299 274756 66300 274820
rect 66364 274756 66365 274820
rect 66299 274755 66365 274756
rect 66115 261764 66181 261765
rect 66115 261700 66116 261764
rect 66180 261700 66181 261764
rect 66115 261699 66181 261700
rect 66118 258090 66178 261699
rect 65934 258030 66178 258090
rect 65934 226405 65994 258030
rect 66670 253877 66730 306330
rect 66954 285592 67574 320058
rect 69614 285701 69674 433603
rect 71454 389061 71514 441627
rect 71635 436388 71701 436389
rect 71635 436324 71636 436388
rect 71700 436324 71701 436388
rect 71635 436323 71701 436324
rect 71451 389060 71517 389061
rect 71451 388996 71452 389060
rect 71516 388996 71517 389060
rect 71451 388995 71517 388996
rect 70899 387836 70965 387837
rect 70899 387772 70900 387836
rect 70964 387772 70965 387836
rect 70899 387771 70965 387772
rect 70163 292636 70229 292637
rect 70163 292572 70164 292636
rect 70228 292572 70229 292636
rect 70163 292571 70229 292572
rect 69611 285700 69677 285701
rect 69611 285636 69612 285700
rect 69676 285636 69677 285700
rect 69611 285635 69677 285636
rect 68875 283660 68941 283661
rect 68875 283596 68876 283660
rect 68940 283596 68941 283660
rect 68875 283595 68941 283596
rect 69979 283660 70045 283661
rect 69979 283596 69980 283660
rect 70044 283596 70045 283660
rect 69979 283595 70045 283596
rect 66667 253876 66733 253877
rect 66667 253812 66668 253876
rect 66732 253812 66733 253876
rect 66667 253811 66733 253812
rect 65931 226404 65997 226405
rect 65931 226340 65932 226404
rect 65996 226340 65997 226404
rect 65931 226339 65997 226340
rect 66670 147933 66730 253811
rect 66954 212614 67574 239592
rect 68878 230621 68938 283595
rect 69982 241637 70042 283595
rect 70166 241773 70226 292571
rect 70347 282980 70413 282981
rect 70347 282916 70348 282980
rect 70412 282916 70413 282980
rect 70347 282915 70413 282916
rect 70163 241772 70229 241773
rect 70163 241708 70164 241772
rect 70228 241708 70229 241772
rect 70163 241707 70229 241708
rect 69979 241636 70045 241637
rect 69979 241572 69980 241636
rect 70044 241572 70045 241636
rect 69979 241571 70045 241572
rect 68875 230620 68941 230621
rect 68875 230556 68876 230620
rect 68940 230556 68941 230620
rect 68875 230555 68941 230556
rect 66954 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 67574 212614
rect 66954 212294 67574 212378
rect 66954 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 67574 212294
rect 66954 176614 67574 212058
rect 68875 203556 68941 203557
rect 68875 203492 68876 203556
rect 68940 203492 68941 203556
rect 68875 203491 68941 203492
rect 66954 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 67574 176614
rect 66954 176294 67574 176378
rect 66954 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 67574 176294
rect 66667 147932 66733 147933
rect 66667 147868 66668 147932
rect 66732 147868 66733 147932
rect 66667 147867 66733 147868
rect 65747 144804 65813 144805
rect 65747 144740 65748 144804
rect 65812 144740 65813 144804
rect 65747 144739 65813 144740
rect 66483 109444 66549 109445
rect 66483 109380 66484 109444
rect 66548 109380 66549 109444
rect 66483 109379 66549 109380
rect 66486 84149 66546 109379
rect 66670 104005 66730 147867
rect 66954 140614 67574 176058
rect 66954 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 67574 140614
rect 66954 140294 67574 140378
rect 66954 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 67574 140294
rect 66954 136782 67574 140058
rect 68139 136916 68205 136917
rect 68139 136852 68140 136916
rect 68204 136852 68205 136916
rect 68139 136851 68205 136852
rect 68142 126853 68202 136851
rect 68139 126852 68205 126853
rect 68139 126788 68140 126852
rect 68204 126788 68205 126852
rect 68139 126787 68205 126788
rect 66667 104004 66733 104005
rect 66667 103940 66668 104004
rect 66732 103940 66733 104004
rect 66667 103939 66733 103940
rect 66851 95844 66917 95845
rect 66851 95780 66852 95844
rect 66916 95780 66917 95844
rect 66851 95779 66917 95780
rect 66854 95029 66914 95779
rect 66851 95028 66917 95029
rect 66851 94964 66852 95028
rect 66916 94964 66917 95028
rect 66851 94963 66917 94964
rect 66483 84148 66549 84149
rect 66483 84084 66484 84148
rect 66548 84084 66549 84148
rect 66483 84083 66549 84084
rect 66954 68614 67574 90782
rect 68878 88229 68938 203491
rect 69611 164388 69677 164389
rect 69611 164324 69612 164388
rect 69676 164324 69677 164388
rect 69611 164323 69677 164324
rect 69614 142170 69674 164323
rect 69246 142110 69674 142170
rect 69246 125629 69306 142110
rect 70350 141405 70410 282915
rect 70902 241773 70962 387771
rect 71638 286109 71698 436323
rect 72374 390421 72434 473995
rect 72739 436252 72805 436253
rect 72739 436188 72740 436252
rect 72804 436188 72805 436252
rect 72739 436187 72805 436188
rect 72371 390420 72437 390421
rect 72371 390356 72372 390420
rect 72436 390356 72437 390420
rect 72371 390355 72437 390356
rect 72742 298757 72802 436187
rect 72978 399454 73298 399486
rect 72978 399218 73020 399454
rect 73256 399218 73298 399454
rect 72978 399134 73298 399218
rect 72978 398898 73020 399134
rect 73256 398898 73298 399134
rect 72978 398866 73298 398898
rect 73478 390421 73538 524995
rect 73794 507454 74414 537166
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 436356 74414 470898
rect 75686 462909 75746 580891
rect 76054 539613 76114 584835
rect 77514 583166 78134 618618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 586894 81854 622338
rect 81234 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 81854 586894
rect 81234 586574 81854 586658
rect 81234 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 81854 586574
rect 81234 583166 81854 586338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 590614 85574 626058
rect 84954 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 85574 590614
rect 84954 590294 85574 590378
rect 84954 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 85574 590294
rect 84954 583166 85574 590058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 583166 92414 596898
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 95514 583166 96134 600618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 79731 580820 79797 580821
rect 79731 580756 79732 580820
rect 79796 580756 79797 580820
rect 79731 580755 79797 580756
rect 83963 580820 84029 580821
rect 83963 580756 83964 580820
rect 84028 580756 84029 580820
rect 83963 580755 84029 580756
rect 88379 580820 88445 580821
rect 88379 580756 88380 580820
rect 88444 580756 88445 580820
rect 88379 580755 88445 580756
rect 91507 580820 91573 580821
rect 91507 580756 91508 580820
rect 91572 580756 91573 580820
rect 91507 580755 91573 580756
rect 77644 561454 77964 561486
rect 77644 561218 77686 561454
rect 77922 561218 77964 561454
rect 77644 561134 77964 561218
rect 77644 560898 77686 561134
rect 77922 560898 77964 561134
rect 77644 560866 77964 560898
rect 76051 539612 76117 539613
rect 76051 539548 76052 539612
rect 76116 539548 76117 539612
rect 76051 539547 76117 539548
rect 77155 523700 77221 523701
rect 77155 523636 77156 523700
rect 77220 523636 77221 523700
rect 77155 523635 77221 523636
rect 75683 462908 75749 462909
rect 75683 462844 75684 462908
rect 75748 462844 75749 462908
rect 75683 462843 75749 462844
rect 73659 435300 73725 435301
rect 73659 435236 73660 435300
rect 73724 435236 73725 435300
rect 73659 435235 73725 435236
rect 73475 390420 73541 390421
rect 73475 390356 73476 390420
rect 73540 390356 73541 390420
rect 73475 390355 73541 390356
rect 73662 388650 73722 435235
rect 74579 434348 74645 434349
rect 74579 434284 74580 434348
rect 74644 434284 74645 434348
rect 74579 434283 74645 434284
rect 75867 434348 75933 434349
rect 75867 434284 75868 434348
rect 75932 434284 75933 434348
rect 75867 434283 75933 434284
rect 73478 388590 73722 388650
rect 73478 387701 73538 388590
rect 73475 387700 73541 387701
rect 73475 387636 73476 387700
rect 73540 387636 73541 387700
rect 73475 387635 73541 387636
rect 73475 387564 73541 387565
rect 73475 387500 73476 387564
rect 73540 387500 73541 387564
rect 73475 387499 73541 387500
rect 72923 385796 72989 385797
rect 72923 385732 72924 385796
rect 72988 385732 72989 385796
rect 72923 385731 72989 385732
rect 72739 298756 72805 298757
rect 72739 298692 72740 298756
rect 72804 298692 72805 298756
rect 72739 298691 72805 298692
rect 71635 286108 71701 286109
rect 71635 286044 71636 286108
rect 71700 286044 71701 286108
rect 71635 286043 71701 286044
rect 72371 284204 72437 284205
rect 72371 284140 72372 284204
rect 72436 284140 72437 284204
rect 72371 284139 72437 284140
rect 72374 241773 72434 284139
rect 70899 241772 70965 241773
rect 70899 241708 70900 241772
rect 70964 241708 70965 241772
rect 70899 241707 70965 241708
rect 72371 241772 72437 241773
rect 72371 241708 72372 241772
rect 72436 241708 72437 241772
rect 72371 241707 72437 241708
rect 72926 241637 72986 385731
rect 73107 283524 73173 283525
rect 73107 283460 73108 283524
rect 73172 283460 73173 283524
rect 73107 283459 73173 283460
rect 72923 241636 72989 241637
rect 72923 241572 72924 241636
rect 72988 241572 72989 241636
rect 72923 241571 72989 241572
rect 72555 240004 72621 240005
rect 72555 239940 72556 240004
rect 72620 239940 72621 240004
rect 72555 239939 72621 239940
rect 72558 229110 72618 239939
rect 72558 229050 72986 229110
rect 72926 215933 72986 229050
rect 72923 215932 72989 215933
rect 72923 215868 72924 215932
rect 72988 215868 72989 215932
rect 72923 215867 72989 215868
rect 71635 208452 71701 208453
rect 71635 208388 71636 208452
rect 71700 208388 71701 208452
rect 71635 208387 71701 208388
rect 70347 141404 70413 141405
rect 70347 141340 70348 141404
rect 70412 141340 70413 141404
rect 70347 141339 70413 141340
rect 69427 138140 69493 138141
rect 69427 138076 69428 138140
rect 69492 138076 69493 138140
rect 69427 138075 69493 138076
rect 69430 131069 69490 138075
rect 70350 138005 70410 141339
rect 70347 138004 70413 138005
rect 70347 137940 70348 138004
rect 70412 137940 70413 138004
rect 70347 137939 70413 137940
rect 69427 131068 69493 131069
rect 69427 131004 69428 131068
rect 69492 131004 69493 131068
rect 69427 131003 69493 131004
rect 69243 125628 69309 125629
rect 69243 125564 69244 125628
rect 69308 125564 69309 125628
rect 69243 125563 69309 125564
rect 69427 99924 69493 99925
rect 69427 99860 69428 99924
rect 69492 99860 69493 99924
rect 69427 99859 69493 99860
rect 69430 93870 69490 99859
rect 69430 93810 69674 93870
rect 68875 88228 68941 88229
rect 68875 88164 68876 88228
rect 68940 88164 68941 88228
rect 68875 88163 68941 88164
rect 69614 80069 69674 93810
rect 71638 91085 71698 208387
rect 72926 92717 72986 215867
rect 73110 140861 73170 283459
rect 73478 241773 73538 387499
rect 73794 363454 74414 388356
rect 74582 364445 74642 434283
rect 75683 433804 75749 433805
rect 75683 433740 75684 433804
rect 75748 433740 75749 433804
rect 75683 433739 75749 433740
rect 74579 364444 74645 364445
rect 74579 364380 74580 364444
rect 74644 364380 74645 364444
rect 74579 364379 74645 364380
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 75686 321605 75746 433739
rect 75683 321604 75749 321605
rect 75683 321540 75684 321604
rect 75748 321540 75749 321604
rect 75683 321539 75749 321540
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 285592 74414 290898
rect 75686 283253 75746 321539
rect 75870 317525 75930 434283
rect 77158 390421 77218 523635
rect 77514 511174 78134 537166
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 475174 78134 510618
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 439174 78134 474618
rect 79734 456109 79794 580755
rect 81609 543454 81929 543486
rect 81609 543218 81651 543454
rect 81887 543218 81929 543454
rect 81609 543134 81929 543218
rect 81609 542898 81651 543134
rect 81887 542898 81929 543134
rect 81609 542866 81929 542898
rect 79915 530772 79981 530773
rect 79915 530708 79916 530772
rect 79980 530708 79981 530772
rect 79915 530707 79981 530708
rect 79731 456108 79797 456109
rect 79731 456044 79732 456108
rect 79796 456044 79797 456108
rect 79731 456043 79797 456044
rect 77514 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 78134 439174
rect 77514 438854 78134 438938
rect 77514 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 78134 438854
rect 77514 436356 78134 438618
rect 78443 437476 78509 437477
rect 78443 437412 78444 437476
rect 78508 437412 78509 437476
rect 78443 437411 78509 437412
rect 78446 436117 78506 437411
rect 78443 436116 78509 436117
rect 78443 436052 78444 436116
rect 78508 436052 78509 436116
rect 78443 436051 78509 436052
rect 77339 433668 77405 433669
rect 77339 433604 77340 433668
rect 77404 433604 77405 433668
rect 77339 433603 77405 433604
rect 77155 390420 77221 390421
rect 77155 390356 77156 390420
rect 77220 390356 77221 390420
rect 77155 390355 77221 390356
rect 77342 318749 77402 433603
rect 77514 367174 78134 388356
rect 78446 387973 78506 436051
rect 78627 433668 78693 433669
rect 78627 433604 78628 433668
rect 78692 433604 78693 433668
rect 78627 433603 78693 433604
rect 78443 387972 78509 387973
rect 78443 387908 78444 387972
rect 78508 387908 78509 387972
rect 78443 387907 78509 387908
rect 78630 380221 78690 433603
rect 79918 390421 79978 530707
rect 81234 514894 81854 537166
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 81234 478894 81854 514338
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 80099 456108 80165 456109
rect 80099 456044 80100 456108
rect 80164 456044 80165 456108
rect 80099 456043 80165 456044
rect 79915 390420 79981 390421
rect 79915 390356 79916 390420
rect 79980 390356 79981 390420
rect 79915 390355 79981 390356
rect 80102 389061 80162 456043
rect 81234 442894 81854 478338
rect 83966 471885 84026 580755
rect 85575 561454 85895 561486
rect 85575 561218 85617 561454
rect 85853 561218 85895 561454
rect 85575 561134 85895 561218
rect 85575 560898 85617 561134
rect 85853 560898 85895 561134
rect 85575 560866 85895 560898
rect 84954 518614 85574 537166
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 84954 482614 85574 518058
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 81939 471884 82005 471885
rect 81939 471820 81940 471884
rect 82004 471820 82005 471884
rect 81939 471819 82005 471820
rect 83963 471884 84029 471885
rect 83963 471820 83964 471884
rect 84028 471820 84029 471884
rect 83963 471819 84029 471820
rect 81234 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 81854 442894
rect 81234 442574 81854 442658
rect 81234 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 81854 442574
rect 81234 436356 81854 442338
rect 80651 434484 80717 434485
rect 80651 434420 80652 434484
rect 80716 434420 80717 434484
rect 80651 434419 80717 434420
rect 78811 389060 78877 389061
rect 78811 388996 78812 389060
rect 78876 388996 78877 389060
rect 78811 388995 78877 388996
rect 80099 389060 80165 389061
rect 80099 388996 80100 389060
rect 80164 388996 80165 389060
rect 80099 388995 80165 388996
rect 78814 384301 78874 388995
rect 78811 384300 78877 384301
rect 78811 384236 78812 384300
rect 78876 384236 78877 384300
rect 78811 384235 78877 384236
rect 78627 380220 78693 380221
rect 78627 380156 78628 380220
rect 78692 380156 78693 380220
rect 78627 380155 78693 380156
rect 77514 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 78134 367174
rect 77514 366854 78134 366938
rect 77514 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 78134 366854
rect 77514 331174 78134 366618
rect 77514 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 78134 331174
rect 77514 330854 78134 330938
rect 77514 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 78134 330854
rect 77339 318748 77405 318749
rect 77339 318684 77340 318748
rect 77404 318684 77405 318748
rect 77339 318683 77405 318684
rect 75867 317524 75933 317525
rect 75867 317460 75868 317524
rect 75932 317460 75933 317524
rect 75867 317459 75933 317460
rect 77514 295174 78134 330618
rect 80654 304197 80714 434419
rect 81942 390421 82002 471819
rect 84954 446614 85574 482058
rect 84954 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 85574 446614
rect 84954 446294 85574 446378
rect 84954 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 85574 446294
rect 84954 436356 85574 446058
rect 88382 438157 88442 580755
rect 89540 543454 89860 543486
rect 89540 543218 89582 543454
rect 89818 543218 89860 543454
rect 89540 543134 89860 543218
rect 89540 542898 89582 543134
rect 89818 542898 89860 543134
rect 89540 542866 89860 542898
rect 91510 525061 91570 580755
rect 99234 568894 99854 604338
rect 99234 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 99854 568894
rect 99234 568574 99854 568658
rect 99234 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 99854 568574
rect 94083 567084 94149 567085
rect 94083 567020 94084 567084
rect 94148 567020 94149 567084
rect 94083 567019 94149 567020
rect 94086 547890 94146 567019
rect 93902 547830 94146 547890
rect 91794 525454 92414 537166
rect 93902 530773 93962 547830
rect 96659 547092 96725 547093
rect 96659 547028 96660 547092
rect 96724 547028 96725 547092
rect 96659 547027 96725 547028
rect 93899 530772 93965 530773
rect 93899 530708 93900 530772
rect 93964 530708 93965 530772
rect 93899 530707 93965 530708
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91507 525060 91573 525061
rect 91507 524996 91508 525060
rect 91572 524996 91573 525060
rect 91507 524995 91573 524996
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 88747 468484 88813 468485
rect 88747 468420 88748 468484
rect 88812 468420 88813 468484
rect 88747 468419 88813 468420
rect 88379 438156 88445 438157
rect 88379 438092 88380 438156
rect 88444 438092 88445 438156
rect 88379 438091 88445 438092
rect 83411 436252 83477 436253
rect 83411 436188 83412 436252
rect 83476 436188 83477 436252
rect 83411 436187 83477 436188
rect 82675 433940 82741 433941
rect 82675 433876 82676 433940
rect 82740 433876 82741 433940
rect 82675 433875 82741 433876
rect 81939 390420 82005 390421
rect 81939 390356 81940 390420
rect 82004 390356 82005 390420
rect 81939 390355 82005 390356
rect 81234 370894 81854 388356
rect 81234 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 81854 370894
rect 81234 370574 81854 370658
rect 81234 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 81854 370574
rect 81234 334894 81854 370338
rect 81234 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 81854 334894
rect 81234 334574 81854 334658
rect 81234 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 81854 334574
rect 80651 304196 80717 304197
rect 80651 304132 80652 304196
rect 80716 304132 80717 304196
rect 80651 304131 80717 304132
rect 77514 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 78134 295174
rect 77514 294854 78134 294938
rect 77514 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 78134 294854
rect 77514 285592 78134 294618
rect 81234 298894 81854 334338
rect 81234 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 81854 298894
rect 81234 298574 81854 298658
rect 81234 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 81854 298574
rect 81234 285592 81854 298338
rect 82678 289101 82738 433875
rect 82859 339556 82925 339557
rect 82859 339492 82860 339556
rect 82924 339492 82925 339556
rect 82859 339491 82925 339492
rect 82862 327045 82922 339491
rect 82859 327044 82925 327045
rect 82859 326980 82860 327044
rect 82924 326980 82925 327044
rect 82859 326979 82925 326980
rect 83414 303653 83474 436187
rect 86171 433804 86237 433805
rect 86171 433740 86172 433804
rect 86236 433740 86237 433804
rect 86171 433739 86237 433740
rect 83595 433668 83661 433669
rect 83595 433604 83596 433668
rect 83660 433604 83661 433668
rect 83595 433603 83661 433604
rect 84147 433668 84213 433669
rect 84147 433604 84148 433668
rect 84212 433604 84213 433668
rect 84147 433603 84213 433604
rect 85251 433668 85317 433669
rect 85251 433604 85252 433668
rect 85316 433604 85317 433668
rect 85251 433603 85317 433604
rect 85803 433668 85869 433669
rect 85803 433604 85804 433668
rect 85868 433604 85869 433668
rect 85803 433603 85869 433604
rect 83598 339557 83658 433603
rect 84150 427830 84210 433603
rect 83966 427770 84210 427830
rect 83966 365669 84026 427770
rect 85254 390693 85314 433603
rect 85251 390692 85317 390693
rect 85251 390628 85252 390692
rect 85316 390628 85317 390692
rect 85251 390627 85317 390628
rect 84954 374614 85574 388356
rect 85806 383757 85866 433603
rect 85803 383756 85869 383757
rect 85803 383692 85804 383756
rect 85868 383692 85869 383756
rect 85803 383691 85869 383692
rect 84954 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 85574 374614
rect 84954 374294 85574 374378
rect 84954 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 85574 374294
rect 83963 365668 84029 365669
rect 83963 365604 83964 365668
rect 84028 365604 84029 365668
rect 83963 365603 84029 365604
rect 83595 339556 83661 339557
rect 83595 339492 83596 339556
rect 83660 339492 83661 339556
rect 83595 339491 83661 339492
rect 84954 338614 85574 374058
rect 84954 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 85574 338614
rect 84954 338294 85574 338378
rect 84954 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 85574 338294
rect 83411 303652 83477 303653
rect 83411 303588 83412 303652
rect 83476 303588 83477 303652
rect 83411 303587 83477 303588
rect 84954 302614 85574 338058
rect 86174 323645 86234 433739
rect 87091 433668 87157 433669
rect 87091 433604 87092 433668
rect 87156 433604 87157 433668
rect 87091 433603 87157 433604
rect 87459 433668 87525 433669
rect 87459 433604 87460 433668
rect 87524 433604 87525 433668
rect 87459 433603 87525 433604
rect 86171 323644 86237 323645
rect 86171 323580 86172 323644
rect 86236 323580 86237 323644
rect 86171 323579 86237 323580
rect 86723 322964 86789 322965
rect 86723 322900 86724 322964
rect 86788 322900 86789 322964
rect 86723 322899 86789 322900
rect 84954 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 85574 302614
rect 84954 302294 85574 302378
rect 84954 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 85574 302294
rect 83411 293180 83477 293181
rect 83411 293116 83412 293180
rect 83476 293116 83477 293180
rect 83411 293115 83477 293116
rect 82675 289100 82741 289101
rect 82675 289036 82676 289100
rect 82740 289036 82741 289100
rect 82675 289035 82741 289036
rect 82678 285701 82738 289035
rect 82675 285700 82741 285701
rect 82675 285636 82676 285700
rect 82740 285636 82741 285700
rect 82675 285635 82741 285636
rect 75683 283252 75749 283253
rect 75683 283188 75684 283252
rect 75748 283188 75749 283252
rect 75683 283187 75749 283188
rect 78977 273454 79297 273486
rect 78977 273218 79019 273454
rect 79255 273218 79297 273454
rect 78977 273134 79297 273218
rect 78977 272898 79019 273134
rect 79255 272898 79297 273134
rect 78977 272866 79297 272898
rect 74345 255454 74665 255486
rect 74345 255218 74387 255454
rect 74623 255218 74665 255454
rect 74345 255134 74665 255218
rect 74345 254898 74387 255134
rect 74623 254898 74665 255134
rect 74345 254866 74665 254898
rect 83414 241773 83474 293115
rect 84954 285592 85574 302058
rect 86171 300796 86237 300797
rect 86171 300732 86172 300796
rect 86236 300732 86237 300796
rect 86171 300731 86237 300732
rect 84699 283660 84765 283661
rect 84699 283596 84700 283660
rect 84764 283596 84765 283660
rect 84699 283595 84765 283596
rect 83963 282980 84029 282981
rect 83963 282916 83964 282980
rect 84028 282916 84029 282980
rect 83963 282915 84029 282916
rect 83966 281890 84026 282915
rect 83966 281830 84394 281890
rect 83609 255454 83929 255486
rect 83609 255218 83651 255454
rect 83887 255218 83929 255454
rect 83609 255134 83929 255218
rect 83609 254898 83651 255134
rect 83887 254898 83929 255134
rect 83609 254866 83929 254898
rect 84334 243130 84394 281830
rect 83966 243070 84394 243130
rect 73475 241772 73541 241773
rect 73475 241708 73476 241772
rect 73540 241708 73541 241772
rect 73475 241707 73541 241708
rect 83411 241772 83477 241773
rect 83411 241708 83412 241772
rect 83476 241708 83477 241772
rect 83411 241707 83477 241708
rect 73794 219454 74414 239592
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73107 140860 73173 140861
rect 73107 140796 73108 140860
rect 73172 140796 73173 140860
rect 73107 140795 73173 140796
rect 73794 136782 74414 146898
rect 77514 223174 78134 239592
rect 77514 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 78134 223174
rect 77514 222854 78134 222938
rect 77514 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 78134 222854
rect 77514 187174 78134 222618
rect 77514 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 78134 187174
rect 77514 186854 78134 186938
rect 77514 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 78134 186854
rect 77514 151174 78134 186618
rect 77514 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 78134 151174
rect 77514 150854 78134 150938
rect 77514 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 78134 150854
rect 77514 136782 78134 150618
rect 81234 226894 81854 239592
rect 83414 238770 83474 241707
rect 83966 241365 84026 243070
rect 84702 241773 84762 283595
rect 86174 241773 86234 300731
rect 86726 241773 86786 322899
rect 87094 318341 87154 433603
rect 87462 378725 87522 433603
rect 88338 417454 88658 417486
rect 88338 417218 88380 417454
rect 88616 417218 88658 417454
rect 88338 417134 88658 417218
rect 88338 416898 88380 417134
rect 88616 416898 88658 417134
rect 88338 416866 88658 416898
rect 88750 389061 88810 468419
rect 91794 453454 92414 488898
rect 95514 529174 96134 537166
rect 96662 530637 96722 547027
rect 96843 541652 96909 541653
rect 96843 541588 96844 541652
rect 96908 541588 96909 541652
rect 96843 541587 96909 541588
rect 96846 531997 96906 541587
rect 99234 532894 99854 568338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102954 572614 103574 608058
rect 102954 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 103574 572614
rect 102954 572294 103574 572378
rect 102954 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 103574 572294
rect 100707 549404 100773 549405
rect 100707 549340 100708 549404
rect 100772 549340 100773 549404
rect 100707 549339 100773 549340
rect 99234 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 99854 532894
rect 99234 532574 99854 532658
rect 99234 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 99854 532574
rect 96843 531996 96909 531997
rect 96843 531932 96844 531996
rect 96908 531932 96909 531996
rect 96843 531931 96909 531932
rect 96659 530636 96725 530637
rect 96659 530572 96660 530636
rect 96724 530572 96725 530636
rect 96659 530571 96725 530572
rect 95514 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 96134 529174
rect 95514 528854 96134 528938
rect 95514 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 96134 528854
rect 95514 493174 96134 528618
rect 95514 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 96134 493174
rect 95514 492854 96134 492938
rect 95514 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 96134 492854
rect 93899 462908 93965 462909
rect 93899 462844 93900 462908
rect 93964 462844 93965 462908
rect 93899 462843 93965 462844
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 90219 436388 90285 436389
rect 90219 436324 90220 436388
rect 90284 436324 90285 436388
rect 91794 436356 92414 452898
rect 90219 436323 90285 436324
rect 89851 433668 89917 433669
rect 89851 433604 89852 433668
rect 89916 433604 89917 433668
rect 89851 433603 89917 433604
rect 88747 389060 88813 389061
rect 88747 388996 88748 389060
rect 88812 388996 88813 389060
rect 88747 388995 88813 388996
rect 87459 378724 87525 378725
rect 87459 378660 87460 378724
rect 87524 378660 87525 378724
rect 87459 378659 87525 378660
rect 88011 351932 88077 351933
rect 88011 351868 88012 351932
rect 88076 351868 88077 351932
rect 88011 351867 88077 351868
rect 87091 318340 87157 318341
rect 87091 318276 87092 318340
rect 87156 318276 87157 318340
rect 87091 318275 87157 318276
rect 87827 282980 87893 282981
rect 87827 282916 87828 282980
rect 87892 282916 87893 282980
rect 87827 282915 87893 282916
rect 84699 241772 84765 241773
rect 84699 241708 84700 241772
rect 84764 241708 84765 241772
rect 84699 241707 84765 241708
rect 86171 241772 86237 241773
rect 86171 241708 86172 241772
rect 86236 241708 86237 241772
rect 86171 241707 86237 241708
rect 86723 241772 86789 241773
rect 86723 241708 86724 241772
rect 86788 241708 86789 241772
rect 86723 241707 86789 241708
rect 83963 241364 84029 241365
rect 83963 241300 83964 241364
rect 84028 241300 84029 241364
rect 83963 241299 84029 241300
rect 84702 240141 84762 241707
rect 84699 240140 84765 240141
rect 84699 240076 84700 240140
rect 84764 240076 84765 240140
rect 84699 240075 84765 240076
rect 81234 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 81854 226894
rect 81234 226574 81854 226658
rect 81234 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 81854 226574
rect 81234 190894 81854 226338
rect 82862 238710 83474 238770
rect 82862 203557 82922 238710
rect 84954 230614 85574 239592
rect 84954 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 85574 230614
rect 84954 230294 85574 230378
rect 84954 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 85574 230294
rect 82859 203556 82925 203557
rect 82859 203492 82860 203556
rect 82924 203492 82925 203556
rect 82859 203491 82925 203492
rect 81234 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 81854 190894
rect 81234 190574 81854 190658
rect 81234 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 81854 190574
rect 81234 154894 81854 190338
rect 81234 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 81854 154894
rect 81234 154574 81854 154658
rect 81234 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 81854 154574
rect 81234 136782 81854 154338
rect 84954 194614 85574 230058
rect 84954 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 85574 194614
rect 84954 194294 85574 194378
rect 84954 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 85574 194294
rect 84954 158614 85574 194058
rect 87830 177309 87890 282915
rect 88014 241773 88074 351867
rect 89854 320789 89914 433603
rect 89851 320788 89917 320789
rect 89851 320724 89852 320788
rect 89916 320724 89917 320788
rect 89851 320723 89917 320724
rect 90222 288421 90282 436323
rect 93902 436117 93962 462843
rect 95514 457174 96134 492618
rect 95514 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 96134 457174
rect 95514 456854 96134 456938
rect 95514 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 96134 456854
rect 95514 436356 96134 456618
rect 99234 496894 99854 532338
rect 99234 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 99854 496894
rect 99234 496574 99854 496658
rect 99234 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 99854 496574
rect 99234 460894 99854 496338
rect 100155 476780 100221 476781
rect 100155 476716 100156 476780
rect 100220 476716 100221 476780
rect 100155 476715 100221 476716
rect 99234 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 99854 460894
rect 99234 460574 99854 460658
rect 99234 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 99854 460574
rect 99234 436356 99854 460338
rect 95003 436252 95069 436253
rect 95003 436188 95004 436252
rect 95068 436188 95069 436252
rect 95003 436187 95069 436188
rect 93899 436116 93965 436117
rect 93899 436052 93900 436116
rect 93964 436052 93965 436116
rect 93899 436051 93965 436052
rect 92979 434620 93045 434621
rect 92979 434556 92980 434620
rect 93044 434556 93045 434620
rect 92979 434555 93045 434556
rect 92611 434212 92677 434213
rect 92611 434148 92612 434212
rect 92676 434148 92677 434212
rect 92611 434147 92677 434148
rect 91323 433804 91389 433805
rect 91323 433740 91324 433804
rect 91388 433740 91389 433804
rect 91323 433739 91389 433740
rect 91326 376005 91386 433739
rect 91507 433668 91573 433669
rect 91507 433604 91508 433668
rect 91572 433604 91573 433668
rect 91507 433603 91573 433604
rect 91510 387837 91570 433603
rect 91507 387836 91573 387837
rect 91507 387772 91508 387836
rect 91572 387772 91573 387836
rect 91507 387771 91573 387772
rect 91794 381454 92414 388356
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91323 376004 91389 376005
rect 91323 375940 91324 376004
rect 91388 375940 91389 376004
rect 91323 375939 91389 375940
rect 91507 376004 91573 376005
rect 91507 375940 91508 376004
rect 91572 375940 91573 376004
rect 91507 375939 91573 375940
rect 90955 321468 91021 321469
rect 90955 321404 90956 321468
rect 91020 321404 91021 321468
rect 90955 321403 91021 321404
rect 90219 288420 90285 288421
rect 90219 288356 90220 288420
rect 90284 288356 90285 288420
rect 90219 288355 90285 288356
rect 88747 285700 88813 285701
rect 88747 285636 88748 285700
rect 88812 285636 88813 285700
rect 88747 285635 88813 285636
rect 88750 282981 88810 285635
rect 89851 283524 89917 283525
rect 89851 283460 89852 283524
rect 89916 283460 89917 283524
rect 89851 283459 89917 283460
rect 88747 282980 88813 282981
rect 88747 282916 88748 282980
rect 88812 282916 88813 282980
rect 88747 282915 88813 282916
rect 88241 273454 88561 273486
rect 88241 273218 88283 273454
rect 88519 273218 88561 273454
rect 88241 273134 88561 273218
rect 88241 272898 88283 273134
rect 88519 272898 88561 273134
rect 88241 272866 88561 272898
rect 88011 241772 88077 241773
rect 88011 241708 88012 241772
rect 88076 241708 88077 241772
rect 88011 241707 88077 241708
rect 87827 177308 87893 177309
rect 87827 177244 87828 177308
rect 87892 177244 87893 177308
rect 87827 177243 87893 177244
rect 87830 176765 87890 177243
rect 87827 176764 87893 176765
rect 87827 176700 87828 176764
rect 87892 176700 87893 176764
rect 87827 176699 87893 176700
rect 84954 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 85574 158614
rect 84954 158294 85574 158378
rect 84954 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 85574 158294
rect 84954 136782 85574 158058
rect 88750 143717 88810 282915
rect 89854 156637 89914 283459
rect 90958 239733 91018 321403
rect 91323 284204 91389 284205
rect 91323 284140 91324 284204
rect 91388 284140 91389 284204
rect 91323 284139 91389 284140
rect 91326 241637 91386 284139
rect 91323 241636 91389 241637
rect 91323 241572 91324 241636
rect 91388 241572 91389 241636
rect 91323 241571 91389 241572
rect 91510 240141 91570 375939
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 92614 330445 92674 434147
rect 92611 330444 92677 330445
rect 92611 330380 92612 330444
rect 92676 330380 92677 330444
rect 92611 330379 92677 330380
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 285592 92414 308898
rect 92982 293317 93042 434555
rect 94819 434348 94885 434349
rect 94819 434284 94820 434348
rect 94884 434284 94885 434348
rect 94819 434283 94885 434284
rect 94822 318885 94882 434283
rect 95006 382261 95066 436187
rect 96291 434348 96357 434349
rect 96291 434284 96292 434348
rect 96356 434284 96357 434348
rect 96291 434283 96357 434284
rect 96294 389605 96354 434283
rect 96843 434212 96909 434213
rect 96843 434148 96844 434212
rect 96908 434148 96909 434212
rect 96843 434147 96909 434148
rect 96475 434076 96541 434077
rect 96475 434012 96476 434076
rect 96540 434012 96541 434076
rect 96475 434011 96541 434012
rect 96291 389604 96357 389605
rect 96291 389540 96292 389604
rect 96356 389540 96357 389604
rect 96291 389539 96357 389540
rect 95514 385174 96134 388356
rect 95514 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 96134 385174
rect 95514 384854 96134 384938
rect 95514 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 96134 384854
rect 95003 382260 95069 382261
rect 95003 382196 95004 382260
rect 95068 382196 95069 382260
rect 95003 382195 95069 382196
rect 95187 381036 95253 381037
rect 95187 380972 95188 381036
rect 95252 380972 95253 381036
rect 95187 380971 95253 380972
rect 95190 374010 95250 380971
rect 95006 373950 95250 374010
rect 94819 318884 94885 318885
rect 94819 318820 94820 318884
rect 94884 318820 94885 318884
rect 94819 318819 94885 318820
rect 94822 316050 94882 318819
rect 94454 315990 94882 316050
rect 94454 294677 94514 315990
rect 94451 294676 94517 294677
rect 94451 294612 94452 294676
rect 94516 294612 94517 294676
rect 94451 294611 94517 294612
rect 92979 293316 93045 293317
rect 92979 293252 92980 293316
rect 93044 293252 93045 293316
rect 92979 293251 93045 293252
rect 92611 283524 92677 283525
rect 92611 283460 92612 283524
rect 92676 283460 92677 283524
rect 92611 283459 92677 283460
rect 91507 240140 91573 240141
rect 91507 240076 91508 240140
rect 91572 240076 91573 240140
rect 91507 240075 91573 240076
rect 90955 239732 91021 239733
rect 90955 239668 90956 239732
rect 91020 239668 91021 239732
rect 90955 239667 91021 239668
rect 91510 219450 91570 240075
rect 91142 219390 91570 219450
rect 91794 237454 92414 239592
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 89851 156636 89917 156637
rect 89851 156572 89852 156636
rect 89916 156572 89917 156636
rect 89851 156571 89917 156572
rect 88747 143716 88813 143717
rect 88747 143652 88748 143716
rect 88812 143652 88813 143716
rect 88747 143651 88813 143652
rect 90955 142220 91021 142221
rect 90955 142156 90956 142220
rect 91020 142156 91021 142220
rect 90955 142155 91021 142156
rect 90958 135285 91018 142155
rect 90955 135284 91021 135285
rect 90955 135220 90956 135284
rect 91020 135220 91021 135284
rect 90955 135219 91021 135220
rect 91142 132970 91202 219390
rect 91794 201454 92414 236898
rect 92614 235789 92674 283459
rect 92873 255454 93193 255486
rect 92873 255218 92915 255454
rect 93151 255218 93193 255454
rect 92873 255134 93193 255218
rect 92873 254898 92915 255134
rect 93151 254898 93193 255134
rect 92873 254866 93193 254898
rect 95006 240141 95066 373950
rect 95514 349174 96134 384618
rect 95514 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 96134 349174
rect 95514 348854 96134 348938
rect 95514 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 96134 348854
rect 95514 313174 96134 348618
rect 95514 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 96134 313174
rect 95514 312854 96134 312938
rect 95514 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 96134 312854
rect 95514 285592 96134 312618
rect 96478 283797 96538 434011
rect 96846 380221 96906 434147
rect 97211 433940 97277 433941
rect 97211 433876 97212 433940
rect 97276 433876 97277 433940
rect 97211 433875 97277 433876
rect 97214 385661 97274 433875
rect 98499 433804 98565 433805
rect 98499 433740 98500 433804
rect 98564 433740 98565 433804
rect 98499 433739 98565 433740
rect 98315 433668 98381 433669
rect 98315 433604 98316 433668
rect 98380 433604 98381 433668
rect 98315 433603 98381 433604
rect 97211 385660 97277 385661
rect 97211 385596 97212 385660
rect 97276 385596 97277 385660
rect 97211 385595 97277 385596
rect 96843 380220 96909 380221
rect 96843 380156 96844 380220
rect 96908 380156 96909 380220
rect 96843 380155 96909 380156
rect 98131 332620 98197 332621
rect 98131 332556 98132 332620
rect 98196 332556 98197 332620
rect 98131 332555 98197 332556
rect 98134 316709 98194 332555
rect 98318 319565 98378 433603
rect 98502 332621 98562 433739
rect 99971 433668 100037 433669
rect 99971 433604 99972 433668
rect 100036 433604 100037 433668
rect 99971 433603 100037 433604
rect 99234 352894 99854 388356
rect 99234 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 99854 352894
rect 99234 352574 99854 352658
rect 99234 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 99854 352574
rect 98499 332620 98565 332621
rect 98499 332556 98500 332620
rect 98564 332556 98565 332620
rect 98499 332555 98565 332556
rect 98315 319564 98381 319565
rect 98315 319500 98316 319564
rect 98380 319500 98381 319564
rect 98315 319499 98381 319500
rect 99234 316894 99854 352338
rect 99974 326365 100034 433603
rect 100158 389061 100218 476715
rect 100710 389061 100770 549339
rect 102954 536614 103574 572058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 104939 571436 105005 571437
rect 104939 571372 104940 571436
rect 105004 571372 105005 571436
rect 104939 571371 105005 571372
rect 102954 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 103574 536614
rect 102954 536294 103574 536378
rect 102954 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 103574 536294
rect 102179 522340 102245 522341
rect 102179 522276 102180 522340
rect 102244 522276 102245 522340
rect 102179 522275 102245 522276
rect 102182 433669 102242 522275
rect 102954 500614 103574 536058
rect 102954 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 103574 500614
rect 102954 500294 103574 500378
rect 102954 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 103574 500294
rect 102954 464614 103574 500058
rect 102954 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 103574 464614
rect 102954 464294 103574 464378
rect 102954 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 103574 464294
rect 102954 436356 103574 464058
rect 103283 436116 103349 436117
rect 103283 436052 103284 436116
rect 103348 436052 103349 436116
rect 103283 436051 103349 436052
rect 100891 433668 100957 433669
rect 100891 433604 100892 433668
rect 100956 433604 100957 433668
rect 100891 433603 100957 433604
rect 102179 433668 102245 433669
rect 102179 433604 102180 433668
rect 102244 433604 102245 433668
rect 102179 433603 102245 433604
rect 100155 389060 100221 389061
rect 100155 388996 100156 389060
rect 100220 388996 100221 389060
rect 100155 388995 100221 388996
rect 100707 389060 100773 389061
rect 100707 388996 100708 389060
rect 100772 388996 100773 389060
rect 100707 388995 100773 388996
rect 100710 381037 100770 388995
rect 100707 381036 100773 381037
rect 100707 380972 100708 381036
rect 100772 380972 100773 381036
rect 100707 380971 100773 380972
rect 100894 373285 100954 433603
rect 102182 387021 102242 433603
rect 103286 390965 103346 436051
rect 104203 433668 104269 433669
rect 104203 433604 104204 433668
rect 104268 433604 104269 433668
rect 104203 433603 104269 433604
rect 103698 399454 104018 399486
rect 103698 399218 103740 399454
rect 103976 399218 104018 399454
rect 103698 399134 104018 399218
rect 103698 398898 103740 399134
rect 103976 398898 104018 399134
rect 103698 398866 104018 398898
rect 103283 390964 103349 390965
rect 103283 390900 103284 390964
rect 103348 390900 103349 390964
rect 103283 390899 103349 390900
rect 102179 387020 102245 387021
rect 102179 386956 102180 387020
rect 102244 386956 102245 387020
rect 102179 386955 102245 386956
rect 100891 373284 100957 373285
rect 100891 373220 100892 373284
rect 100956 373220 100957 373284
rect 100891 373219 100957 373220
rect 102954 356614 103574 388356
rect 102954 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 103574 356614
rect 102954 356294 103574 356378
rect 102954 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 103574 356294
rect 99971 326364 100037 326365
rect 99971 326300 99972 326364
rect 100036 326300 100037 326364
rect 99971 326299 100037 326300
rect 98131 316708 98197 316709
rect 98131 316644 98132 316708
rect 98196 316644 98197 316708
rect 98131 316643 98197 316644
rect 99234 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 99854 316894
rect 99234 316574 99854 316658
rect 99234 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 99854 316574
rect 97947 287332 98013 287333
rect 97947 287268 97948 287332
rect 98012 287268 98013 287332
rect 97947 287267 98013 287268
rect 97950 284885 98010 287267
rect 99234 285592 99854 316338
rect 102954 320614 103574 356058
rect 104206 353973 104266 433603
rect 104942 389061 105002 571371
rect 109794 543454 110414 578898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 110643 559468 110709 559469
rect 110643 559404 110644 559468
rect 110708 559404 110709 559468
rect 110643 559403 110709 559404
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 107699 479500 107765 479501
rect 107699 479436 107700 479500
rect 107764 479436 107765 479500
rect 107699 479435 107765 479436
rect 106411 468620 106477 468621
rect 106411 468556 106412 468620
rect 106476 468556 106477 468620
rect 106411 468555 106477 468556
rect 106414 441630 106474 468555
rect 106230 441570 106474 441630
rect 105123 436116 105189 436117
rect 105123 436052 105124 436116
rect 105188 436052 105189 436116
rect 105123 436051 105189 436052
rect 105126 433669 105186 436051
rect 105123 433668 105189 433669
rect 105123 433604 105124 433668
rect 105188 433604 105189 433668
rect 105123 433603 105189 433604
rect 104939 389060 105005 389061
rect 104939 388996 104940 389060
rect 105004 388996 105005 389060
rect 104939 388995 105005 388996
rect 104203 353972 104269 353973
rect 104203 353908 104204 353972
rect 104268 353908 104269 353972
rect 104203 353907 104269 353908
rect 102954 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 103574 320614
rect 102954 320294 103574 320378
rect 102954 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 103574 320294
rect 101259 294676 101325 294677
rect 101259 294612 101260 294676
rect 101324 294612 101325 294676
rect 101259 294611 101325 294612
rect 100707 291956 100773 291957
rect 100707 291892 100708 291956
rect 100772 291892 100773 291956
rect 100707 291891 100773 291892
rect 97947 284884 98013 284885
rect 97947 284820 97948 284884
rect 98012 284820 98013 284884
rect 97947 284819 98013 284820
rect 95187 283796 95253 283797
rect 95187 283732 95188 283796
rect 95252 283732 95253 283796
rect 95187 283731 95253 283732
rect 96475 283796 96541 283797
rect 96475 283732 96476 283796
rect 96540 283732 96541 283796
rect 96475 283731 96541 283732
rect 95003 240140 95069 240141
rect 95003 240076 95004 240140
rect 95068 240076 95069 240140
rect 95003 240075 95069 240076
rect 93715 238236 93781 238237
rect 93715 238172 93716 238236
rect 93780 238172 93781 238236
rect 93715 238171 93781 238172
rect 92611 235788 92677 235789
rect 92611 235724 92612 235788
rect 92676 235724 92677 235788
rect 92611 235723 92677 235724
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 136782 92414 164898
rect 91142 132910 91754 132970
rect 77644 129454 77964 129486
rect 77644 129218 77686 129454
rect 77922 129218 77964 129454
rect 77644 129134 77964 129218
rect 77644 128898 77686 129134
rect 77922 128898 77964 129134
rect 77644 128866 77964 128898
rect 85575 129454 85895 129486
rect 85575 129218 85617 129454
rect 85853 129218 85895 129454
rect 85575 129134 85895 129218
rect 85575 128898 85617 129134
rect 85853 128898 85895 129134
rect 85575 128866 85895 128898
rect 73679 111454 73999 111486
rect 73679 111218 73721 111454
rect 73957 111218 73999 111454
rect 73679 111134 73999 111218
rect 73679 110898 73721 111134
rect 73957 110898 73999 111134
rect 73679 110866 73999 110898
rect 81609 111454 81929 111486
rect 81609 111218 81651 111454
rect 81887 111218 81929 111454
rect 81609 111134 81929 111218
rect 81609 110898 81651 111134
rect 81887 110898 81929 111134
rect 81609 110866 81929 110898
rect 89540 111454 89860 111486
rect 89540 111218 89582 111454
rect 89818 111218 89860 111454
rect 89540 111134 89860 111218
rect 89540 110898 89582 111134
rect 89818 110898 89860 111134
rect 89540 110866 89860 110898
rect 72923 92716 72989 92717
rect 72923 92652 72924 92716
rect 72988 92652 72989 92716
rect 72923 92651 72989 92652
rect 91694 92445 91754 132910
rect 93718 92717 93778 238171
rect 95190 237013 95250 283731
rect 98867 282980 98933 282981
rect 98867 282916 98868 282980
rect 98932 282916 98933 282980
rect 98867 282915 98933 282916
rect 98870 277405 98930 282915
rect 100710 282709 100770 291891
rect 100707 282708 100773 282709
rect 100707 282644 100708 282708
rect 100772 282644 100773 282708
rect 100707 282643 100773 282644
rect 101262 278629 101322 294611
rect 102954 284614 103574 320058
rect 102954 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 103574 284614
rect 102954 284294 103574 284378
rect 102954 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 103574 284294
rect 101259 278628 101325 278629
rect 101259 278564 101260 278628
rect 101324 278564 101325 278628
rect 101259 278563 101325 278564
rect 98867 277404 98933 277405
rect 98867 277340 98868 277404
rect 98932 277340 98933 277404
rect 98867 277339 98933 277340
rect 99971 256732 100037 256733
rect 99971 256668 99972 256732
rect 100036 256668 100037 256732
rect 99971 256667 100037 256668
rect 98131 255372 98197 255373
rect 98131 255308 98132 255372
rect 98196 255308 98197 255372
rect 98131 255307 98197 255308
rect 97763 240140 97829 240141
rect 97763 240076 97764 240140
rect 97828 240076 97829 240140
rect 97763 240075 97829 240076
rect 95187 237012 95253 237013
rect 95187 236948 95188 237012
rect 95252 236948 95253 237012
rect 95187 236947 95253 236948
rect 95514 205174 96134 239592
rect 97766 209790 97826 240075
rect 98134 234630 98194 255307
rect 99974 242589 100034 256667
rect 102954 248614 103574 284058
rect 102954 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 103574 248614
rect 102954 248294 103574 248378
rect 102954 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 103574 248294
rect 99971 242588 100037 242589
rect 99971 242524 99972 242588
rect 100036 242524 100037 242588
rect 99971 242523 100037 242524
rect 97214 209730 97826 209790
rect 97950 234570 98194 234630
rect 97214 207093 97274 209730
rect 97211 207092 97277 207093
rect 97211 207028 97212 207092
rect 97276 207028 97277 207092
rect 97211 207027 97277 207028
rect 95514 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 96134 205174
rect 95514 204854 96134 204938
rect 95514 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 96134 204854
rect 95514 169174 96134 204618
rect 95514 168938 95546 169174
rect 95782 168938 95866 169174
rect 96102 168938 96134 169174
rect 95514 168854 96134 168938
rect 95514 168618 95546 168854
rect 95782 168618 95866 168854
rect 96102 168618 96134 168854
rect 94819 136916 94885 136917
rect 94819 136852 94820 136916
rect 94884 136852 94885 136916
rect 94819 136851 94885 136852
rect 94822 133789 94882 136851
rect 95514 136782 96134 168618
rect 95739 135284 95805 135285
rect 95739 135220 95740 135284
rect 95804 135220 95805 135284
rect 95739 135219 95805 135220
rect 94819 133788 94885 133789
rect 94819 133724 94820 133788
rect 94884 133724 94885 133788
rect 94819 133723 94885 133724
rect 95742 118557 95802 135219
rect 95739 118556 95805 118557
rect 95739 118492 95740 118556
rect 95804 118492 95805 118556
rect 95739 118491 95805 118492
rect 97214 92853 97274 207027
rect 97395 124268 97461 124269
rect 97395 124204 97396 124268
rect 97460 124204 97461 124268
rect 97395 124203 97461 124204
rect 97211 92852 97277 92853
rect 97211 92788 97212 92852
rect 97276 92788 97277 92852
rect 97211 92787 97277 92788
rect 93715 92716 93781 92717
rect 93715 92652 93716 92716
rect 93780 92652 93781 92716
rect 93715 92651 93781 92652
rect 91691 92444 91757 92445
rect 91691 92380 91692 92444
rect 91756 92380 91757 92444
rect 91691 92379 91757 92380
rect 97398 92173 97458 124203
rect 97950 108901 98010 234570
rect 99234 208894 99854 239592
rect 99234 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 99854 208894
rect 99234 208574 99854 208658
rect 99234 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 99854 208574
rect 99234 172894 99854 208338
rect 99234 172658 99266 172894
rect 99502 172658 99586 172894
rect 99822 172658 99854 172894
rect 99234 172574 99854 172658
rect 99234 172338 99266 172574
rect 99502 172338 99586 172574
rect 99822 172338 99854 172574
rect 99234 136894 99854 172338
rect 102954 212614 103574 248058
rect 104942 241501 105002 388995
rect 105126 384301 105186 433603
rect 106230 390965 106290 441570
rect 106411 433668 106477 433669
rect 106411 433604 106412 433668
rect 106476 433604 106477 433668
rect 106411 433603 106477 433604
rect 106227 390964 106293 390965
rect 106227 390900 106228 390964
rect 106292 390900 106293 390964
rect 106227 390899 106293 390900
rect 105123 384300 105189 384301
rect 105123 384236 105124 384300
rect 105188 384236 105189 384300
rect 105123 384235 105189 384236
rect 106414 374645 106474 433603
rect 107702 390557 107762 479435
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109539 439516 109605 439517
rect 109539 439452 109540 439516
rect 109604 439452 109605 439516
rect 109539 439451 109605 439452
rect 108987 434348 109053 434349
rect 108987 434284 108988 434348
rect 109052 434284 109053 434348
rect 108987 434283 109053 434284
rect 108990 434210 109050 434283
rect 108806 434150 109050 434210
rect 108435 433804 108501 433805
rect 108435 433740 108436 433804
rect 108500 433740 108501 433804
rect 108435 433739 108501 433740
rect 108438 427830 108498 433739
rect 108806 428770 108866 434150
rect 109542 434077 109602 439451
rect 109794 436356 110414 470898
rect 109539 434076 109605 434077
rect 109539 434012 109540 434076
rect 109604 434012 109605 434076
rect 109539 434011 109605 434012
rect 110646 433669 110706 559403
rect 113514 547174 114134 582618
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 111747 534716 111813 534717
rect 111747 534652 111748 534716
rect 111812 534652 111813 534716
rect 111747 534651 111813 534652
rect 110643 433668 110709 433669
rect 110643 433604 110644 433668
rect 110708 433604 110709 433668
rect 110643 433603 110709 433604
rect 108806 428710 109050 428770
rect 108438 427770 108866 427830
rect 108806 398850 108866 427770
rect 108622 398790 108866 398850
rect 107699 390556 107765 390557
rect 107699 390492 107700 390556
rect 107764 390492 107765 390556
rect 107699 390491 107765 390492
rect 108622 390285 108682 398790
rect 108990 398170 109050 428710
rect 108806 398110 109050 398170
rect 108619 390284 108685 390285
rect 108619 390220 108620 390284
rect 108684 390220 108685 390284
rect 108619 390219 108685 390220
rect 108806 389190 108866 398110
rect 111750 390421 111810 534651
rect 113514 511174 114134 546618
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 113514 475174 114134 510618
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 113514 439174 114134 474618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117234 550894 117854 586338
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 514894 117854 550338
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 117234 478894 117854 514338
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 114323 450532 114389 450533
rect 114323 450468 114324 450532
rect 114388 450468 114389 450532
rect 114323 450467 114389 450468
rect 113514 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 114134 439174
rect 113514 438854 114134 438938
rect 113514 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 114134 438854
rect 113514 436356 114134 438618
rect 112115 434076 112181 434077
rect 112115 434012 112116 434076
rect 112180 434012 112181 434076
rect 112115 434011 112181 434012
rect 111931 433668 111997 433669
rect 111931 433604 111932 433668
rect 111996 433604 111997 433668
rect 111931 433603 111997 433604
rect 111747 390420 111813 390421
rect 111747 390356 111748 390420
rect 111812 390356 111813 390420
rect 111747 390355 111813 390356
rect 108806 389130 109050 389190
rect 108251 384300 108317 384301
rect 108251 384236 108252 384300
rect 108316 384236 108317 384300
rect 108251 384235 108317 384236
rect 106411 374644 106477 374645
rect 106411 374580 106412 374644
rect 106476 374580 106477 374644
rect 106411 374579 106477 374580
rect 108254 268565 108314 384235
rect 108990 376005 109050 389130
rect 108987 376004 109053 376005
rect 108987 375940 108988 376004
rect 109052 375940 109053 376004
rect 108987 375939 109053 375940
rect 109794 363454 110414 388356
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 111934 327725 111994 433603
rect 112118 432853 112178 434011
rect 112115 432852 112181 432853
rect 112115 432788 112116 432852
rect 112180 432788 112181 432852
rect 112115 432787 112181 432788
rect 114326 399533 114386 450467
rect 117234 442894 117854 478338
rect 117234 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 117854 442894
rect 117234 442574 117854 442658
rect 117234 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 117854 442574
rect 115979 440332 116045 440333
rect 115979 440268 115980 440332
rect 116044 440268 116045 440332
rect 115979 440267 116045 440268
rect 114507 417892 114573 417893
rect 114507 417828 114508 417892
rect 114572 417828 114573 417892
rect 114507 417827 114573 417828
rect 114323 399532 114389 399533
rect 114323 399468 114324 399532
rect 114388 399468 114389 399532
rect 114323 399467 114389 399468
rect 113514 367174 114134 388356
rect 113514 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 114134 367174
rect 113514 366854 114134 366938
rect 113514 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 114134 366854
rect 113514 331174 114134 366618
rect 113514 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 114134 331174
rect 113514 330854 114134 330938
rect 113514 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 114134 330854
rect 111931 327724 111997 327725
rect 111931 327660 111932 327724
rect 111996 327660 111997 327724
rect 111931 327659 111997 327660
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 108251 268564 108317 268565
rect 108251 268500 108252 268564
rect 108316 268500 108317 268564
rect 108251 268499 108317 268500
rect 108251 266388 108317 266389
rect 108251 266324 108252 266388
rect 108316 266324 108317 266388
rect 108251 266323 108317 266324
rect 108254 260813 108314 266323
rect 108435 262852 108501 262853
rect 108435 262788 108436 262852
rect 108500 262788 108501 262852
rect 108435 262787 108501 262788
rect 108251 260812 108317 260813
rect 108251 260748 108252 260812
rect 108316 260748 108317 260812
rect 108251 260747 108317 260748
rect 108438 258090 108498 262787
rect 108254 258030 108498 258090
rect 108254 254557 108314 258030
rect 109794 255454 110414 290898
rect 113514 295174 114134 330618
rect 113514 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 114134 295174
rect 113514 294854 114134 294938
rect 113514 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 114134 294854
rect 110643 267068 110709 267069
rect 110643 267004 110644 267068
rect 110708 267004 110709 267068
rect 110643 267003 110709 267004
rect 110646 265029 110706 267003
rect 110643 265028 110709 265029
rect 110643 264964 110644 265028
rect 110708 264964 110709 265028
rect 110643 264963 110709 264964
rect 113514 259174 114134 294618
rect 114510 271149 114570 417827
rect 114691 408644 114757 408645
rect 114691 408580 114692 408644
rect 114756 408580 114757 408644
rect 114691 408579 114757 408580
rect 114694 318341 114754 408579
rect 115982 319429 116042 440267
rect 117234 406894 117854 442338
rect 117234 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 117854 406894
rect 117234 406574 117854 406658
rect 117234 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 117854 406574
rect 117234 370894 117854 406338
rect 117234 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 117854 370894
rect 117234 370574 117854 370658
rect 117234 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 117854 370574
rect 117234 334894 117854 370338
rect 117234 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 117854 334894
rect 117234 334574 117854 334658
rect 117234 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 117854 334574
rect 115979 319428 116045 319429
rect 115979 319364 115980 319428
rect 116044 319364 116045 319428
rect 115979 319363 116045 319364
rect 114691 318340 114757 318341
rect 114691 318276 114692 318340
rect 114756 318276 114757 318340
rect 114691 318275 114757 318276
rect 117234 298894 117854 334338
rect 117234 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 117854 298894
rect 117234 298574 117854 298658
rect 117234 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 117854 298574
rect 114507 271148 114573 271149
rect 114507 271084 114508 271148
rect 114572 271084 114573 271148
rect 114507 271083 114573 271084
rect 113514 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 114134 259174
rect 113514 258854 114134 258938
rect 111011 258772 111077 258773
rect 111011 258708 111012 258772
rect 111076 258708 111077 258772
rect 111011 258707 111077 258708
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 108251 254556 108317 254557
rect 108251 254492 108252 254556
rect 108316 254492 108317 254556
rect 108251 254491 108317 254492
rect 104939 241500 105005 241501
rect 104939 241436 104940 241500
rect 105004 241436 105005 241500
rect 104939 241435 105005 241436
rect 108254 221645 108314 254491
rect 108251 221644 108317 221645
rect 108251 221580 108252 221644
rect 108316 221580 108317 221644
rect 108251 221579 108317 221580
rect 102954 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 103574 212614
rect 102954 212294 103574 212378
rect 102954 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 103574 212294
rect 102954 176614 103574 212058
rect 109794 219454 110414 254898
rect 111014 241365 111074 258707
rect 113514 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 114134 258854
rect 111011 241364 111077 241365
rect 111011 241300 111012 241364
rect 111076 241300 111077 241364
rect 111011 241299 111077 241300
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 105491 196756 105557 196757
rect 105491 196692 105492 196756
rect 105556 196692 105557 196756
rect 105491 196691 105557 196692
rect 102954 176378 102986 176614
rect 103222 176378 103306 176614
rect 103542 176378 103574 176614
rect 102954 176294 103574 176378
rect 102954 176058 102986 176294
rect 103222 176058 103306 176294
rect 103542 176058 103574 176294
rect 100707 145620 100773 145621
rect 100707 145556 100708 145620
rect 100772 145556 100773 145620
rect 100707 145555 100773 145556
rect 99234 136658 99266 136894
rect 99502 136658 99586 136894
rect 99822 136658 99854 136894
rect 99234 136574 99854 136658
rect 99234 136338 99266 136574
rect 99502 136338 99586 136574
rect 99822 136338 99854 136574
rect 97947 108900 98013 108901
rect 97947 108836 97948 108900
rect 98012 108836 98013 108900
rect 97947 108835 98013 108836
rect 99234 100894 99854 136338
rect 99234 100658 99266 100894
rect 99502 100658 99586 100894
rect 99822 100658 99854 100894
rect 99234 100574 99854 100658
rect 99234 100338 99266 100574
rect 99502 100338 99586 100574
rect 99822 100338 99854 100574
rect 97395 92172 97461 92173
rect 97395 92108 97396 92172
rect 97460 92108 97461 92172
rect 97395 92107 97461 92108
rect 71635 91084 71701 91085
rect 71635 91020 71636 91084
rect 71700 91020 71701 91084
rect 71635 91019 71701 91020
rect 69611 80068 69677 80069
rect 69611 80004 69612 80068
rect 69676 80004 69677 80068
rect 69611 80003 69677 80004
rect 66954 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 67574 68614
rect 66954 68294 67574 68378
rect 66954 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 67574 68294
rect 66954 32614 67574 68058
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 65379 4044 65445 4045
rect 65379 3980 65380 4044
rect 65444 3980 65445 4044
rect 65379 3979 65445 3980
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 75454 74414 90782
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 79174 78134 90782
rect 77514 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 78134 79174
rect 77514 78854 78134 78938
rect 77514 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 78134 78854
rect 77514 43174 78134 78618
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 82894 81854 90782
rect 81234 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 81854 82894
rect 81234 82574 81854 82658
rect 81234 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 81854 82574
rect 81234 46894 81854 82338
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 86614 85574 90782
rect 84954 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 85574 86614
rect 84954 86294 85574 86378
rect 84954 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 85574 86294
rect 84954 50614 85574 86058
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 57454 92414 90782
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 61174 96134 90782
rect 95514 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 96134 61174
rect 95514 60854 96134 60938
rect 95514 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 96134 60854
rect 95514 25174 96134 60618
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 64894 99854 100338
rect 100710 91085 100770 145555
rect 102954 140614 103574 176058
rect 102954 140378 102986 140614
rect 103222 140378 103306 140614
rect 103542 140378 103574 140614
rect 102954 140294 103574 140378
rect 102954 140058 102986 140294
rect 103222 140058 103306 140294
rect 103542 140058 103574 140294
rect 102954 104614 103574 140058
rect 102954 104378 102986 104614
rect 103222 104378 103306 104614
rect 103542 104378 103574 104614
rect 102954 104294 103574 104378
rect 102954 104058 102986 104294
rect 103222 104058 103306 104294
rect 103542 104058 103574 104294
rect 100707 91084 100773 91085
rect 100707 91020 100708 91084
rect 100772 91020 100773 91084
rect 100707 91019 100773 91020
rect 99234 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 99854 64894
rect 99234 64574 99854 64658
rect 99234 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 99854 64574
rect 99234 28894 99854 64338
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 68614 103574 104058
rect 102954 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 103574 68614
rect 102954 68294 103574 68378
rect 102954 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 103574 68294
rect 102954 32614 103574 68058
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 105494 3501 105554 196691
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 105491 3500 105557 3501
rect 105491 3436 105492 3500
rect 105556 3436 105557 3500
rect 105491 3435 105557 3436
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 223174 114134 258618
rect 113514 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 114134 223174
rect 113514 222854 114134 222938
rect 113514 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 114134 222854
rect 113514 187174 114134 222618
rect 113514 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 114134 187174
rect 113514 186854 114134 186938
rect 113514 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 114134 186854
rect 113514 151174 114134 186618
rect 113514 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 114134 151174
rect 113514 150854 114134 150938
rect 113514 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 114134 150854
rect 113514 115174 114134 150618
rect 113514 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 114134 115174
rect 113514 114854 114134 114938
rect 113514 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 114134 114854
rect 113514 79174 114134 114618
rect 113514 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 114134 79174
rect 113514 78854 114134 78938
rect 113514 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 114134 78854
rect 113514 43174 114134 78618
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 262894 117854 298338
rect 117234 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 117854 262894
rect 117234 262574 117854 262658
rect 117234 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 117854 262574
rect 117234 226894 117854 262338
rect 117234 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 117854 226894
rect 117234 226574 117854 226658
rect 117234 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 117854 226574
rect 117234 190894 117854 226338
rect 117234 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 117854 190894
rect 117234 190574 117854 190658
rect 117234 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 117854 190574
rect 117234 154894 117854 190338
rect 117234 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 117854 154894
rect 117234 154574 117854 154658
rect 117234 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 117854 154574
rect 117234 118894 117854 154338
rect 117234 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 117854 118894
rect 117234 118574 117854 118658
rect 117234 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 117854 118574
rect 117234 82894 117854 118338
rect 117234 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 117854 82894
rect 117234 82574 117854 82658
rect 117234 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 117854 82574
rect 117234 46894 117854 82338
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 125731 590748 125797 590749
rect 125731 590684 125732 590748
rect 125796 590684 125797 590748
rect 125731 590683 125797 590684
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 120954 554614 121574 590058
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 518614 121574 554058
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 120954 482614 121574 518058
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120954 446614 121574 482058
rect 120954 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 121574 446614
rect 120954 446294 121574 446378
rect 120954 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 121574 446294
rect 120954 410614 121574 446058
rect 120954 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 121574 410614
rect 120954 410294 121574 410378
rect 120954 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 121574 410294
rect 120954 374614 121574 410058
rect 125734 389061 125794 590683
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 125731 389060 125797 389061
rect 125731 388996 125732 389060
rect 125796 388996 125797 389060
rect 125731 388995 125797 388996
rect 120954 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 121574 374614
rect 120954 374294 121574 374378
rect 120954 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 121574 374294
rect 120954 338614 121574 374058
rect 120954 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 121574 338614
rect 120954 338294 121574 338378
rect 120954 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 121574 338294
rect 120954 302614 121574 338058
rect 120954 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 121574 302614
rect 120954 302294 121574 302378
rect 120954 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 121574 302294
rect 120954 266614 121574 302058
rect 120954 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 121574 266614
rect 120954 266294 121574 266378
rect 120954 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 121574 266294
rect 120954 230614 121574 266058
rect 125734 234565 125794 388995
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 125731 234564 125797 234565
rect 125731 234500 125732 234564
rect 125796 234500 125797 234564
rect 125731 234499 125797 234500
rect 120954 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 121574 230614
rect 120954 230294 121574 230378
rect 120954 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 121574 230294
rect 120954 194614 121574 230058
rect 120954 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 121574 194614
rect 120954 194294 121574 194378
rect 120954 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 121574 194294
rect 120954 158614 121574 194058
rect 120954 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 121574 158614
rect 120954 158294 121574 158378
rect 120954 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 121574 158294
rect 120954 122614 121574 158058
rect 120954 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 121574 122614
rect 120954 122294 121574 122378
rect 120954 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 121574 122294
rect 120954 86614 121574 122058
rect 120954 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 121574 86614
rect 120954 86294 121574 86378
rect 120954 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 121574 86294
rect 120954 50614 121574 86058
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 127794 165454 128414 200898
rect 127794 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 128414 165454
rect 127794 165134 128414 165218
rect 127794 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 128414 165134
rect 127794 129454 128414 164898
rect 127794 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 128414 129454
rect 127794 129134 128414 129218
rect 127794 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 128414 129134
rect 127794 93454 128414 128898
rect 127794 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 128414 93454
rect 127794 93134 128414 93218
rect 127794 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 128414 93134
rect 127794 57454 128414 92898
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 529174 132134 564618
rect 131514 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 132134 529174
rect 131514 528854 132134 528938
rect 131514 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 132134 528854
rect 131514 493174 132134 528618
rect 131514 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 132134 493174
rect 131514 492854 132134 492938
rect 131514 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 132134 492854
rect 131514 457174 132134 492618
rect 131514 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 132134 457174
rect 131514 456854 132134 456938
rect 131514 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 132134 456854
rect 131514 421174 132134 456618
rect 131514 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 132134 421174
rect 131514 420854 132134 420938
rect 131514 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 132134 420854
rect 131514 385174 132134 420618
rect 131514 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 132134 385174
rect 131514 384854 132134 384938
rect 131514 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 132134 384854
rect 131514 349174 132134 384618
rect 131514 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 132134 349174
rect 131514 348854 132134 348938
rect 131514 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 132134 348854
rect 131514 313174 132134 348618
rect 131514 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 132134 313174
rect 131514 312854 132134 312938
rect 131514 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 132134 312854
rect 131514 277174 132134 312618
rect 131514 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 132134 277174
rect 131514 276854 132134 276938
rect 131514 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 132134 276854
rect 131514 241174 132134 276618
rect 131514 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 132134 241174
rect 131514 240854 132134 240938
rect 131514 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 132134 240854
rect 131514 205174 132134 240618
rect 131514 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 132134 205174
rect 131514 204854 132134 204938
rect 131514 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 132134 204854
rect 131514 169174 132134 204618
rect 131514 168938 131546 169174
rect 131782 168938 131866 169174
rect 132102 168938 132134 169174
rect 131514 168854 132134 168938
rect 131514 168618 131546 168854
rect 131782 168618 131866 168854
rect 132102 168618 132134 168854
rect 131514 133174 132134 168618
rect 131514 132938 131546 133174
rect 131782 132938 131866 133174
rect 132102 132938 132134 133174
rect 131514 132854 132134 132938
rect 131514 132618 131546 132854
rect 131782 132618 131866 132854
rect 132102 132618 132134 132854
rect 131514 97174 132134 132618
rect 131514 96938 131546 97174
rect 131782 96938 131866 97174
rect 132102 96938 132134 97174
rect 131514 96854 132134 96938
rect 131514 96618 131546 96854
rect 131782 96618 131866 96854
rect 132102 96618 132134 96854
rect 131514 61174 132134 96618
rect 131514 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 132134 61174
rect 131514 60854 132134 60938
rect 131514 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 132134 60854
rect 131514 25174 132134 60618
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 532894 135854 568338
rect 135234 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 135854 532894
rect 135234 532574 135854 532658
rect 135234 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 135854 532574
rect 135234 496894 135854 532338
rect 135234 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 135854 496894
rect 135234 496574 135854 496658
rect 135234 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 135854 496574
rect 135234 460894 135854 496338
rect 135234 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 135854 460894
rect 135234 460574 135854 460658
rect 135234 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 135854 460574
rect 135234 424894 135854 460338
rect 135234 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 135854 424894
rect 135234 424574 135854 424658
rect 135234 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 135854 424574
rect 135234 388894 135854 424338
rect 135234 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 135854 388894
rect 135234 388574 135854 388658
rect 135234 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 135854 388574
rect 135234 352894 135854 388338
rect 135234 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 135854 352894
rect 135234 352574 135854 352658
rect 135234 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 135854 352574
rect 135234 316894 135854 352338
rect 135234 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 135854 316894
rect 135234 316574 135854 316658
rect 135234 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 135854 316574
rect 135234 280894 135854 316338
rect 135234 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 135854 280894
rect 135234 280574 135854 280658
rect 135234 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 135854 280574
rect 135234 244894 135854 280338
rect 135234 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 135854 244894
rect 135234 244574 135854 244658
rect 135234 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 135854 244574
rect 135234 208894 135854 244338
rect 135234 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 135854 208894
rect 135234 208574 135854 208658
rect 135234 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 135854 208574
rect 135234 172894 135854 208338
rect 135234 172658 135266 172894
rect 135502 172658 135586 172894
rect 135822 172658 135854 172894
rect 135234 172574 135854 172658
rect 135234 172338 135266 172574
rect 135502 172338 135586 172574
rect 135822 172338 135854 172574
rect 135234 136894 135854 172338
rect 135234 136658 135266 136894
rect 135502 136658 135586 136894
rect 135822 136658 135854 136894
rect 135234 136574 135854 136658
rect 135234 136338 135266 136574
rect 135502 136338 135586 136574
rect 135822 136338 135854 136574
rect 135234 100894 135854 136338
rect 135234 100658 135266 100894
rect 135502 100658 135586 100894
rect 135822 100658 135854 100894
rect 135234 100574 135854 100658
rect 135234 100338 135266 100574
rect 135502 100338 135586 100574
rect 135822 100338 135854 100574
rect 135234 64894 135854 100338
rect 135234 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 135854 64894
rect 135234 64574 135854 64658
rect 135234 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 135854 64574
rect 135234 28894 135854 64338
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 536614 139574 572058
rect 138954 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 139574 536614
rect 138954 536294 139574 536378
rect 138954 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 139574 536294
rect 138954 500614 139574 536058
rect 138954 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 139574 500614
rect 138954 500294 139574 500378
rect 138954 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 139574 500294
rect 138954 464614 139574 500058
rect 138954 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 139574 464614
rect 138954 464294 139574 464378
rect 138954 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 139574 464294
rect 138954 428614 139574 464058
rect 138954 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 139574 428614
rect 138954 428294 139574 428378
rect 138954 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 139574 428294
rect 138954 392614 139574 428058
rect 138954 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 139574 392614
rect 138954 392294 139574 392378
rect 138954 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 139574 392294
rect 138954 356614 139574 392058
rect 138954 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 139574 356614
rect 138954 356294 139574 356378
rect 138954 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 139574 356294
rect 138954 320614 139574 356058
rect 138954 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 139574 320614
rect 138954 320294 139574 320378
rect 138954 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 139574 320294
rect 138954 284614 139574 320058
rect 138954 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 139574 284614
rect 138954 284294 139574 284378
rect 138954 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 139574 284294
rect 138954 248614 139574 284058
rect 138954 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 139574 248614
rect 138954 248294 139574 248378
rect 138954 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 139574 248294
rect 138954 212614 139574 248058
rect 138954 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 139574 212614
rect 138954 212294 139574 212378
rect 138954 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 139574 212294
rect 138954 176614 139574 212058
rect 138954 176378 138986 176614
rect 139222 176378 139306 176614
rect 139542 176378 139574 176614
rect 138954 176294 139574 176378
rect 138954 176058 138986 176294
rect 139222 176058 139306 176294
rect 139542 176058 139574 176294
rect 138954 140614 139574 176058
rect 138954 140378 138986 140614
rect 139222 140378 139306 140614
rect 139542 140378 139574 140614
rect 138954 140294 139574 140378
rect 138954 140058 138986 140294
rect 139222 140058 139306 140294
rect 139542 140058 139574 140294
rect 138954 104614 139574 140058
rect 138954 104378 138986 104614
rect 139222 104378 139306 104614
rect 139542 104378 139574 104614
rect 138954 104294 139574 104378
rect 138954 104058 138986 104294
rect 139222 104058 139306 104294
rect 139542 104058 139574 104294
rect 138954 68614 139574 104058
rect 138954 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 139574 68614
rect 138954 68294 139574 68378
rect 138954 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 139574 68294
rect 138954 32614 139574 68058
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 147454 146414 182898
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 111454 146414 146898
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 145794 75454 146414 110898
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 149514 475174 150134 510618
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 439174 150134 474618
rect 149514 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 150134 439174
rect 149514 438854 150134 438938
rect 149514 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 150134 438854
rect 149514 403174 150134 438618
rect 149514 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 150134 403174
rect 149514 402854 150134 402938
rect 149514 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 150134 402854
rect 149514 367174 150134 402618
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 149514 331174 150134 366618
rect 149514 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 150134 331174
rect 149514 330854 150134 330938
rect 149514 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 150134 330854
rect 149514 295174 150134 330618
rect 149514 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 150134 295174
rect 149514 294854 150134 294938
rect 149514 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 150134 294854
rect 149514 259174 150134 294618
rect 149514 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 150134 259174
rect 149514 258854 150134 258938
rect 149514 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 150134 258854
rect 149514 223174 150134 258618
rect 149514 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 150134 223174
rect 149514 222854 150134 222938
rect 149514 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 150134 222854
rect 149514 187174 150134 222618
rect 149514 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 150134 187174
rect 149514 186854 150134 186938
rect 149514 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 150134 186854
rect 149514 151174 150134 186618
rect 149514 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 150134 151174
rect 149514 150854 150134 150938
rect 149514 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 150134 150854
rect 149514 115174 150134 150618
rect 149514 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 150134 115174
rect 149514 114854 150134 114938
rect 149514 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 150134 114854
rect 149514 79174 150134 114618
rect 149514 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 150134 79174
rect 149514 78854 150134 78938
rect 149514 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 150134 78854
rect 149514 43174 150134 78618
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 514894 153854 550338
rect 153234 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 153854 514894
rect 153234 514574 153854 514658
rect 153234 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 153854 514574
rect 153234 478894 153854 514338
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 442894 153854 478338
rect 153234 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 153854 442894
rect 153234 442574 153854 442658
rect 153234 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 153854 442574
rect 153234 406894 153854 442338
rect 153234 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 153854 406894
rect 153234 406574 153854 406658
rect 153234 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 153854 406574
rect 153234 370894 153854 406338
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 153234 334894 153854 370338
rect 153234 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 153854 334894
rect 153234 334574 153854 334658
rect 153234 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 153854 334574
rect 153234 298894 153854 334338
rect 153234 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 153854 298894
rect 153234 298574 153854 298658
rect 153234 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 153854 298574
rect 153234 262894 153854 298338
rect 153234 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 153854 262894
rect 153234 262574 153854 262658
rect 153234 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 153854 262574
rect 153234 226894 153854 262338
rect 153234 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 153854 226894
rect 153234 226574 153854 226658
rect 153234 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 153854 226574
rect 153234 190894 153854 226338
rect 153234 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 153854 190894
rect 153234 190574 153854 190658
rect 153234 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 153854 190574
rect 153234 154894 153854 190338
rect 153234 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 153854 154894
rect 153234 154574 153854 154658
rect 153234 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 153854 154574
rect 153234 118894 153854 154338
rect 153234 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 153854 118894
rect 153234 118574 153854 118658
rect 153234 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 153854 118574
rect 153234 82894 153854 118338
rect 153234 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 153854 82894
rect 153234 82574 153854 82658
rect 153234 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 153854 82574
rect 153234 46894 153854 82338
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 518614 157574 554058
rect 156954 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 157574 518614
rect 156954 518294 157574 518378
rect 156954 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 157574 518294
rect 156954 482614 157574 518058
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156954 446614 157574 482058
rect 156954 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 157574 446614
rect 156954 446294 157574 446378
rect 156954 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 157574 446294
rect 156954 410614 157574 446058
rect 156954 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 157574 410614
rect 156954 410294 157574 410378
rect 156954 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 157574 410294
rect 156954 374614 157574 410058
rect 156954 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 157574 374614
rect 156954 374294 157574 374378
rect 156954 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 157574 374294
rect 156954 338614 157574 374058
rect 156954 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 157574 338614
rect 156954 338294 157574 338378
rect 156954 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 157574 338294
rect 156954 302614 157574 338058
rect 156954 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 157574 302614
rect 156954 302294 157574 302378
rect 156954 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 157574 302294
rect 156954 266614 157574 302058
rect 156954 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 157574 266614
rect 156954 266294 157574 266378
rect 156954 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 157574 266294
rect 156954 230614 157574 266058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 160691 263668 160757 263669
rect 160691 263604 160692 263668
rect 160756 263604 160757 263668
rect 160691 263603 160757 263604
rect 156954 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 157574 230614
rect 156954 230294 157574 230378
rect 156954 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 157574 230294
rect 156954 194614 157574 230058
rect 156954 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 157574 194614
rect 156954 194294 157574 194378
rect 156954 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 157574 194294
rect 156954 158614 157574 194058
rect 156954 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 157574 158614
rect 156954 158294 157574 158378
rect 156954 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 157574 158294
rect 156954 122614 157574 158058
rect 156954 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 157574 122614
rect 156954 122294 157574 122378
rect 156954 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 157574 122294
rect 156954 86614 157574 122058
rect 156954 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 157574 86614
rect 156954 86294 157574 86378
rect 156954 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 157574 86294
rect 156954 50614 157574 86058
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 160694 8941 160754 263603
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 163794 165454 164414 200898
rect 163794 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 164414 165454
rect 163794 165134 164414 165218
rect 163794 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 164414 165134
rect 163794 129454 164414 164898
rect 163794 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 164414 129454
rect 163794 129134 164414 129218
rect 163794 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 164414 129134
rect 163794 93454 164414 128898
rect 163794 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 164414 93454
rect 163794 93134 164414 93218
rect 163794 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 164414 93134
rect 163794 57454 164414 92898
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 160691 8940 160757 8941
rect 160691 8876 160692 8940
rect 160756 8876 160757 8940
rect 160691 8875 160757 8876
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 565174 168134 600618
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 529174 168134 564618
rect 167514 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 168134 529174
rect 167514 528854 168134 528938
rect 167514 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 168134 528854
rect 167514 493174 168134 528618
rect 167514 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 168134 493174
rect 167514 492854 168134 492938
rect 167514 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 168134 492854
rect 167514 457174 168134 492618
rect 167514 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 168134 457174
rect 167514 456854 168134 456938
rect 167514 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 168134 456854
rect 167514 421174 168134 456618
rect 167514 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 168134 421174
rect 167514 420854 168134 420938
rect 167514 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 168134 420854
rect 167514 385174 168134 420618
rect 167514 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 168134 385174
rect 167514 384854 168134 384938
rect 167514 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 168134 384854
rect 167514 349174 168134 384618
rect 167514 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 168134 349174
rect 167514 348854 168134 348938
rect 167514 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 168134 348854
rect 167514 313174 168134 348618
rect 167514 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 168134 313174
rect 167514 312854 168134 312938
rect 167514 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 168134 312854
rect 167514 277174 168134 312618
rect 167514 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 168134 277174
rect 167514 276854 168134 276938
rect 167514 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 168134 276854
rect 167514 241174 168134 276618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 171234 568894 171854 604338
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 171234 532894 171854 568338
rect 171234 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 171854 532894
rect 171234 532574 171854 532658
rect 171234 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 171854 532574
rect 171234 496894 171854 532338
rect 171234 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 171854 496894
rect 171234 496574 171854 496658
rect 171234 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 171854 496574
rect 171234 460894 171854 496338
rect 171234 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 171854 460894
rect 171234 460574 171854 460658
rect 171234 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 171854 460574
rect 171234 424894 171854 460338
rect 171234 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 171854 424894
rect 171234 424574 171854 424658
rect 171234 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 171854 424574
rect 171234 388894 171854 424338
rect 171234 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 171854 388894
rect 171234 388574 171854 388658
rect 171234 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 171854 388574
rect 171234 352894 171854 388338
rect 171234 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 171854 352894
rect 171234 352574 171854 352658
rect 171234 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 171854 352574
rect 171234 316894 171854 352338
rect 171234 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 171854 316894
rect 171234 316574 171854 316658
rect 171234 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 171854 316574
rect 171234 280894 171854 316338
rect 171234 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 171854 280894
rect 171234 280574 171854 280658
rect 171234 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 171854 280574
rect 171234 244894 171854 280338
rect 171234 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 171854 244894
rect 171234 244574 171854 244658
rect 168971 244356 169037 244357
rect 168971 244292 168972 244356
rect 169036 244292 169037 244356
rect 168971 244291 169037 244292
rect 171234 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 171854 244574
rect 167514 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 168134 241174
rect 167514 240854 168134 240938
rect 167514 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 168134 240854
rect 167514 205174 168134 240618
rect 167514 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 168134 205174
rect 167514 204854 168134 204938
rect 167514 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 168134 204854
rect 167514 169174 168134 204618
rect 167514 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 168134 169174
rect 167514 168854 168134 168938
rect 167514 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 168134 168854
rect 167514 133174 168134 168618
rect 167514 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 168134 133174
rect 167514 132854 168134 132938
rect 167514 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 168134 132854
rect 167514 97174 168134 132618
rect 167514 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 168134 97174
rect 167514 96854 168134 96938
rect 167514 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 168134 96854
rect 167514 61174 168134 96618
rect 167514 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 168134 61174
rect 167514 60854 168134 60938
rect 167514 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 168134 60854
rect 167514 25174 168134 60618
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 168974 4861 169034 244291
rect 171234 208894 171854 244338
rect 171234 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 171854 208894
rect 171234 208574 171854 208658
rect 171234 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 171854 208574
rect 171234 172894 171854 208338
rect 171234 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 171854 172894
rect 171234 172574 171854 172658
rect 171234 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 171854 172574
rect 171234 136894 171854 172338
rect 171234 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 171854 136894
rect 171234 136574 171854 136658
rect 171234 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 171854 136574
rect 171234 100894 171854 136338
rect 171234 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 171854 100894
rect 171234 100574 171854 100658
rect 171234 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 171854 100574
rect 171234 64894 171854 100338
rect 171234 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 171854 64894
rect 171234 64574 171854 64658
rect 171234 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 171854 64574
rect 171234 28894 171854 64338
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 168971 4860 169037 4861
rect 168971 4796 168972 4860
rect 169036 4796 169037 4860
rect 168971 4795 169037 4796
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 572614 175574 608058
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 536614 175574 572058
rect 174954 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 175574 536614
rect 174954 536294 175574 536378
rect 174954 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 175574 536294
rect 174954 500614 175574 536058
rect 174954 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 175574 500614
rect 174954 500294 175574 500378
rect 174954 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 175574 500294
rect 174954 464614 175574 500058
rect 174954 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 175574 464614
rect 174954 464294 175574 464378
rect 174954 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 175574 464294
rect 174954 428614 175574 464058
rect 174954 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 175574 428614
rect 174954 428294 175574 428378
rect 174954 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 175574 428294
rect 174954 392614 175574 428058
rect 174954 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 175574 392614
rect 174954 392294 175574 392378
rect 174954 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 175574 392294
rect 174954 356614 175574 392058
rect 174954 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 175574 356614
rect 174954 356294 175574 356378
rect 174954 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 175574 356294
rect 174954 320614 175574 356058
rect 174954 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 175574 320614
rect 174954 320294 175574 320378
rect 174954 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 175574 320294
rect 174954 284614 175574 320058
rect 174954 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 175574 284614
rect 174954 284294 175574 284378
rect 174954 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 175574 284294
rect 174954 248614 175574 284058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 178539 258228 178605 258229
rect 178539 258164 178540 258228
rect 178604 258164 178605 258228
rect 178539 258163 178605 258164
rect 174954 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 175574 248614
rect 174954 248294 175574 248378
rect 174954 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 175574 248294
rect 174954 212614 175574 248058
rect 174954 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 175574 212614
rect 174954 212294 175574 212378
rect 174954 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 175574 212294
rect 174954 176614 175574 212058
rect 174954 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 175574 176614
rect 174954 176294 175574 176378
rect 174954 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 175574 176294
rect 174954 140614 175574 176058
rect 174954 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 175574 140614
rect 174954 140294 175574 140378
rect 174954 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 175574 140294
rect 174954 104614 175574 140058
rect 174954 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 175574 104614
rect 174954 104294 175574 104378
rect 174954 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 175574 104294
rect 174954 68614 175574 104058
rect 174954 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 175574 68614
rect 174954 68294 175574 68378
rect 174954 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 175574 68294
rect 174954 32614 175574 68058
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 178542 10301 178602 258163
rect 181794 255454 182414 290898
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 547174 186134 582618
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 475174 186134 510618
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 439174 186134 474618
rect 185514 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 186134 439174
rect 185514 438854 186134 438938
rect 185514 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 186134 438854
rect 185514 403174 186134 438618
rect 185514 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 186134 403174
rect 185514 402854 186134 402938
rect 185514 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 186134 402854
rect 185514 367174 186134 402618
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 185514 331174 186134 366618
rect 185514 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 186134 331174
rect 185514 330854 186134 330938
rect 185514 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 186134 330854
rect 185514 295174 186134 330618
rect 185514 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 186134 295174
rect 185514 294854 186134 294938
rect 185514 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 186134 294854
rect 184059 274684 184125 274685
rect 184059 274620 184060 274684
rect 184124 274620 184125 274684
rect 184059 274619 184125 274620
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 184062 144125 184122 274619
rect 185514 259174 186134 294618
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 185514 223174 186134 258618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 550894 189854 586338
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 514894 189854 550338
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 189234 478894 189854 514338
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 189234 442894 189854 478338
rect 189234 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 189854 442894
rect 189234 442574 189854 442658
rect 189234 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 189854 442574
rect 189234 406894 189854 442338
rect 189234 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 189854 406894
rect 189234 406574 189854 406658
rect 189234 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 189854 406574
rect 189234 370894 189854 406338
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 189234 334894 189854 370338
rect 189234 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 189854 334894
rect 189234 334574 189854 334658
rect 189234 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 189854 334574
rect 189234 298894 189854 334338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 554614 193574 590058
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 518614 193574 554058
rect 192954 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 193574 518614
rect 192954 518294 193574 518378
rect 192954 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 193574 518294
rect 192954 482614 193574 518058
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 192954 446614 193574 482058
rect 192954 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 193574 446614
rect 192954 446294 193574 446378
rect 192954 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 193574 446294
rect 192954 410614 193574 446058
rect 192954 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 193574 410614
rect 192954 410294 193574 410378
rect 192954 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 193574 410294
rect 192954 374614 193574 410058
rect 192954 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 193574 374614
rect 192954 374294 193574 374378
rect 192954 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 193574 374294
rect 192954 338614 193574 374058
rect 192954 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 193574 338614
rect 192954 338294 193574 338378
rect 192954 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 193574 338294
rect 192954 303592 193574 338058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 203514 565174 204134 600618
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 203514 529174 204134 564618
rect 203514 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 204134 529174
rect 203514 528854 204134 528938
rect 203514 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 204134 528854
rect 203514 493174 204134 528618
rect 203514 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 204134 493174
rect 203514 492854 204134 492938
rect 203514 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 204134 492854
rect 203514 457174 204134 492618
rect 203514 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 204134 457174
rect 203514 456854 204134 456938
rect 203514 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 204134 456854
rect 203514 421174 204134 456618
rect 203514 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 204134 421174
rect 203514 420854 204134 420938
rect 203514 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 204134 420854
rect 203514 385174 204134 420618
rect 203514 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 204134 385174
rect 203514 384854 204134 384938
rect 203514 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 204134 384854
rect 203514 349174 204134 384618
rect 203514 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 204134 349174
rect 203514 348854 204134 348938
rect 203514 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 204134 348854
rect 203514 313174 204134 348618
rect 203514 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 204134 313174
rect 203514 312854 204134 312938
rect 203514 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 204134 312854
rect 201539 310860 201605 310861
rect 201539 310796 201540 310860
rect 201604 310796 201605 310860
rect 201539 310795 201605 310796
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 197307 306508 197373 306509
rect 197307 306444 197308 306508
rect 197372 306444 197373 306508
rect 197307 306443 197373 306444
rect 193443 302292 193509 302293
rect 193443 302228 193444 302292
rect 193508 302228 193509 302292
rect 193443 302227 193509 302228
rect 193259 301884 193325 301885
rect 193259 301820 193260 301884
rect 193324 301820 193325 301884
rect 193259 301819 193325 301820
rect 189234 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 189854 298894
rect 189234 298574 189854 298658
rect 189234 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 189854 298574
rect 189234 262894 189854 298338
rect 193262 296717 193322 301819
rect 193446 298893 193506 302227
rect 194547 300932 194613 300933
rect 194547 300868 194548 300932
rect 194612 300868 194613 300932
rect 194547 300867 194613 300868
rect 193443 298892 193509 298893
rect 193443 298828 193444 298892
rect 193508 298828 193509 298892
rect 193443 298827 193509 298828
rect 193259 296716 193325 296717
rect 193259 296652 193260 296716
rect 193324 296652 193325 296716
rect 193259 296651 193325 296652
rect 193075 296580 193141 296581
rect 193075 296516 193076 296580
rect 193140 296516 193141 296580
rect 193075 296515 193141 296516
rect 191603 295220 191669 295221
rect 191603 295156 191604 295220
rect 191668 295156 191669 295220
rect 191603 295155 191669 295156
rect 189234 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 189854 262894
rect 189234 262574 189854 262658
rect 189234 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 189854 262574
rect 188291 253196 188357 253197
rect 188291 253132 188292 253196
rect 188356 253132 188357 253196
rect 188291 253131 188357 253132
rect 185514 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 186134 223174
rect 185514 222854 186134 222938
rect 185514 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 186134 222854
rect 184795 213348 184861 213349
rect 184795 213284 184796 213348
rect 184860 213284 184861 213348
rect 184795 213283 184861 213284
rect 184798 212669 184858 213283
rect 184795 212668 184861 212669
rect 184795 212604 184796 212668
rect 184860 212604 184861 212668
rect 184795 212603 184861 212604
rect 184059 144124 184125 144125
rect 184059 144060 184060 144124
rect 184124 144060 184125 144124
rect 184059 144059 184125 144060
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 184798 96661 184858 212603
rect 185514 187174 186134 222618
rect 188294 212533 188354 253131
rect 189234 226894 189854 262338
rect 189234 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 189854 226894
rect 189234 226574 189854 226658
rect 189234 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 189854 226574
rect 188291 212532 188357 212533
rect 188291 212468 188292 212532
rect 188356 212468 188357 212532
rect 188291 212467 188357 212468
rect 188843 211172 188909 211173
rect 188843 211108 188844 211172
rect 188908 211108 188909 211172
rect 188843 211107 188909 211108
rect 185514 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 186134 187174
rect 185514 186854 186134 186938
rect 185514 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 186134 186854
rect 185514 151174 186134 186618
rect 187555 164388 187621 164389
rect 187555 164324 187556 164388
rect 187620 164324 187621 164388
rect 187555 164323 187621 164324
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 185514 115174 186134 150618
rect 187558 131205 187618 164323
rect 187555 131204 187621 131205
rect 187555 131140 187556 131204
rect 187620 131140 187621 131204
rect 187555 131139 187621 131140
rect 185514 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 186134 115174
rect 185514 114854 186134 114938
rect 185514 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 186134 114854
rect 184795 96660 184861 96661
rect 184795 96596 184796 96660
rect 184860 96596 184861 96660
rect 184795 96595 184861 96596
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 178539 10300 178605 10301
rect 178539 10236 178540 10300
rect 178604 10236 178605 10300
rect 178539 10235 178605 10236
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 79174 186134 114618
rect 186819 109172 186885 109173
rect 186819 109108 186820 109172
rect 186884 109108 186885 109172
rect 186819 109107 186885 109108
rect 186822 92309 186882 109107
rect 188846 95301 188906 211107
rect 189234 190894 189854 226338
rect 190315 208452 190381 208453
rect 190315 208388 190316 208452
rect 190380 208388 190381 208452
rect 190315 208387 190381 208388
rect 189234 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 189854 190894
rect 189234 190574 189854 190658
rect 189234 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 189854 190574
rect 189234 154894 189854 190338
rect 189234 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 189854 154894
rect 189234 154574 189854 154658
rect 189234 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 189854 154574
rect 189234 118894 189854 154338
rect 189234 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 189854 118894
rect 189234 118574 189854 118658
rect 189234 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 189854 118574
rect 188843 95300 188909 95301
rect 188843 95236 188844 95300
rect 188908 95236 188909 95300
rect 188843 95235 188909 95236
rect 186819 92308 186885 92309
rect 186819 92244 186820 92308
rect 186884 92244 186885 92308
rect 186819 92243 186885 92244
rect 185514 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 186134 79174
rect 185514 78854 186134 78938
rect 185514 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 186134 78854
rect 185514 43174 186134 78618
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 82894 189854 118338
rect 190318 91901 190378 208387
rect 191606 129301 191666 295155
rect 192891 242180 192957 242181
rect 192891 242116 192892 242180
rect 192956 242116 192957 242180
rect 192891 242115 192957 242116
rect 192894 240957 192954 242115
rect 193078 241501 193138 296515
rect 193995 286516 194061 286517
rect 193995 286452 193996 286516
rect 194060 286452 194061 286516
rect 193995 286451 194061 286452
rect 193259 247620 193325 247621
rect 193259 247556 193260 247620
rect 193324 247556 193325 247620
rect 193259 247555 193325 247556
rect 193262 242861 193322 247555
rect 193259 242860 193325 242861
rect 193259 242796 193260 242860
rect 193324 242796 193325 242860
rect 193259 242795 193325 242796
rect 193075 241500 193141 241501
rect 193075 241436 193076 241500
rect 193140 241436 193141 241500
rect 193075 241435 193141 241436
rect 192891 240956 192957 240957
rect 192891 240892 192892 240956
rect 192956 240892 192957 240956
rect 192891 240891 192957 240892
rect 192954 230614 193574 239592
rect 192954 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 193574 230614
rect 192954 230294 193574 230378
rect 192954 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 193574 230294
rect 192954 194614 193574 230058
rect 192954 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 193574 194614
rect 192954 194294 193574 194378
rect 192954 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 193574 194294
rect 192954 158614 193574 194058
rect 192954 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 193574 158614
rect 192954 158294 193574 158378
rect 192954 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 193574 158294
rect 192707 147116 192773 147117
rect 192707 147052 192708 147116
rect 192772 147052 192773 147116
rect 192707 147051 192773 147052
rect 191603 129300 191669 129301
rect 191603 129236 191604 129300
rect 191668 129236 191669 129300
rect 191603 129235 191669 129236
rect 192339 124268 192405 124269
rect 192339 124204 192340 124268
rect 192404 124204 192405 124268
rect 192339 124203 192405 124204
rect 192155 118692 192221 118693
rect 192155 118628 192156 118692
rect 192220 118628 192221 118692
rect 192155 118627 192221 118628
rect 192158 117333 192218 118627
rect 192155 117332 192221 117333
rect 192155 117268 192156 117332
rect 192220 117268 192221 117332
rect 192155 117267 192221 117268
rect 190315 91900 190381 91901
rect 190315 91836 190316 91900
rect 190380 91836 190381 91900
rect 190315 91835 190381 91836
rect 192342 91221 192402 124203
rect 192710 120325 192770 147051
rect 192954 143035 193574 158058
rect 193259 139636 193325 139637
rect 193259 139572 193260 139636
rect 193324 139572 193325 139636
rect 193259 139571 193325 139572
rect 193262 125765 193322 139571
rect 193259 125764 193325 125765
rect 193259 125700 193260 125764
rect 193324 125700 193325 125764
rect 193259 125699 193325 125700
rect 193811 125628 193877 125629
rect 193811 125564 193812 125628
rect 193876 125564 193877 125628
rect 193811 125563 193877 125564
rect 192707 120324 192773 120325
rect 192707 120260 192708 120324
rect 192772 120260 192773 120324
rect 192707 120259 192773 120260
rect 192707 117332 192773 117333
rect 192707 117268 192708 117332
rect 192772 117268 192773 117332
rect 192707 117267 192773 117268
rect 192339 91220 192405 91221
rect 192339 91156 192340 91220
rect 192404 91156 192405 91220
rect 192339 91155 192405 91156
rect 189234 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 189854 82894
rect 189234 82574 189854 82658
rect 189234 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 189854 82574
rect 189234 46894 189854 82338
rect 192710 73813 192770 117267
rect 192954 86614 193574 90782
rect 193814 87549 193874 125563
rect 193998 92853 194058 286451
rect 194550 196621 194610 300867
rect 196571 300796 196637 300797
rect 196571 300732 196572 300796
rect 196636 300732 196637 300796
rect 196571 300731 196637 300732
rect 195835 231164 195901 231165
rect 195835 231100 195836 231164
rect 195900 231100 195901 231164
rect 195835 231099 195901 231100
rect 194547 196620 194613 196621
rect 194547 196556 194548 196620
rect 194612 196556 194613 196620
rect 194547 196555 194613 196556
rect 195838 92853 195898 231099
rect 196574 202197 196634 300731
rect 197310 300661 197370 306443
rect 199794 303592 200414 308898
rect 201542 308277 201602 310795
rect 201539 308276 201605 308277
rect 201539 308212 201540 308276
rect 201604 308212 201605 308276
rect 201539 308211 201605 308212
rect 198779 300932 198845 300933
rect 198779 300868 198780 300932
rect 198844 300868 198845 300932
rect 198779 300867 198845 300868
rect 197307 300660 197373 300661
rect 197307 300596 197308 300660
rect 197372 300596 197373 300660
rect 197307 300595 197373 300596
rect 197776 291454 198096 291486
rect 197776 291218 197818 291454
rect 198054 291218 198096 291454
rect 197776 291134 198096 291218
rect 197776 290898 197818 291134
rect 198054 290898 198096 291134
rect 197776 290866 198096 290898
rect 197776 255454 198096 255486
rect 197776 255218 197818 255454
rect 198054 255218 198096 255454
rect 197776 255134 198096 255218
rect 197776 254898 197818 255134
rect 198054 254898 198096 255134
rect 197776 254866 198096 254898
rect 198782 237285 198842 300867
rect 201542 240277 201602 308211
rect 203514 303592 204134 312618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 532894 207854 568338
rect 207234 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 207854 532894
rect 207234 532574 207854 532658
rect 207234 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 207854 532574
rect 207234 496894 207854 532338
rect 207234 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 207854 496894
rect 207234 496574 207854 496658
rect 207234 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 207854 496574
rect 207234 460894 207854 496338
rect 207234 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 207854 460894
rect 207234 460574 207854 460658
rect 207234 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 207854 460574
rect 207234 424894 207854 460338
rect 207234 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 207854 424894
rect 207234 424574 207854 424658
rect 207234 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 207854 424574
rect 207234 388894 207854 424338
rect 207234 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 207854 388894
rect 207234 388574 207854 388658
rect 207234 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 207854 388574
rect 207234 352894 207854 388338
rect 207234 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 207854 352894
rect 207234 352574 207854 352658
rect 207234 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 207854 352574
rect 207234 316894 207854 352338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 536614 211574 572058
rect 210954 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 211574 536614
rect 210954 536294 211574 536378
rect 210954 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 211574 536294
rect 210954 500614 211574 536058
rect 210954 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 211574 500614
rect 210954 500294 211574 500378
rect 210954 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 211574 500294
rect 210954 464614 211574 500058
rect 210954 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 211574 464614
rect 210954 464294 211574 464378
rect 210954 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 211574 464294
rect 210954 428614 211574 464058
rect 210954 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 211574 428614
rect 210954 428294 211574 428378
rect 210954 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 211574 428294
rect 210954 392614 211574 428058
rect 210954 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 211574 392614
rect 210954 392294 211574 392378
rect 210954 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 211574 392294
rect 210954 356614 211574 392058
rect 210954 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 211574 356614
rect 210954 356294 211574 356378
rect 210954 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 211574 356294
rect 210954 320614 211574 356058
rect 210954 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 211574 320614
rect 210954 320294 211574 320378
rect 210371 320244 210437 320245
rect 210371 320180 210372 320244
rect 210436 320180 210437 320244
rect 210371 320179 210437 320180
rect 207234 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 207854 316894
rect 207234 316574 207854 316658
rect 207234 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 207854 316574
rect 207234 303592 207854 316338
rect 204851 300932 204917 300933
rect 204851 300868 204852 300932
rect 204916 300868 204917 300932
rect 204851 300867 204917 300868
rect 205771 300932 205837 300933
rect 205771 300868 205772 300932
rect 205836 300868 205837 300932
rect 205771 300867 205837 300868
rect 207059 300932 207125 300933
rect 207059 300868 207060 300932
rect 207124 300868 207125 300932
rect 207059 300867 207125 300868
rect 201539 240276 201605 240277
rect 201539 240212 201540 240276
rect 201604 240212 201605 240276
rect 201539 240211 201605 240212
rect 199794 237454 200414 239592
rect 198779 237284 198845 237285
rect 198779 237220 198780 237284
rect 198844 237220 198845 237284
rect 198779 237219 198845 237220
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 196571 202196 196637 202197
rect 196571 202132 196572 202196
rect 196636 202132 196637 202196
rect 196571 202131 196637 202132
rect 199794 201454 200414 236898
rect 201539 223548 201605 223549
rect 201539 223484 201540 223548
rect 201604 223484 201605 223548
rect 201539 223483 201605 223484
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 201355 186964 201421 186965
rect 201355 186900 201356 186964
rect 201420 186900 201421 186964
rect 201355 186899 201421 186900
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 198779 143716 198845 143717
rect 198779 143652 198780 143716
rect 198844 143652 198845 143716
rect 198779 143651 198845 143652
rect 196571 142356 196637 142357
rect 196571 142292 196572 142356
rect 196636 142292 196637 142356
rect 196571 142291 196637 142292
rect 193995 92852 194061 92853
rect 193995 92788 193996 92852
rect 194060 92788 194061 92852
rect 193995 92787 194061 92788
rect 195835 92852 195901 92853
rect 195835 92788 195836 92852
rect 195900 92788 195901 92852
rect 195835 92787 195901 92788
rect 193811 87548 193877 87549
rect 193811 87484 193812 87548
rect 193876 87484 193877 87548
rect 193811 87483 193877 87484
rect 192954 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 193574 86614
rect 192954 86294 193574 86378
rect 192954 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 193574 86294
rect 192707 73812 192773 73813
rect 192707 73748 192708 73812
rect 192772 73748 192773 73812
rect 192707 73747 192773 73748
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 50614 193574 86058
rect 196574 58581 196634 142291
rect 197123 142220 197189 142221
rect 197123 142156 197124 142220
rect 197188 142156 197189 142220
rect 197123 142155 197189 142156
rect 196571 58580 196637 58581
rect 196571 58516 196572 58580
rect 196636 58516 196637 58580
rect 196571 58515 196637 58516
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 197126 24173 197186 142155
rect 198782 141133 198842 143651
rect 199794 143035 200414 164898
rect 200619 142220 200685 142221
rect 200619 142156 200620 142220
rect 200684 142156 200685 142220
rect 200619 142155 200685 142156
rect 198779 141132 198845 141133
rect 198779 141068 198780 141132
rect 198844 141068 198845 141132
rect 198779 141067 198845 141068
rect 199388 111454 199708 111486
rect 199388 111218 199430 111454
rect 199666 111218 199708 111454
rect 199388 111134 199708 111218
rect 199388 110898 199430 111134
rect 199666 110898 199708 111134
rect 199388 110866 199708 110898
rect 200622 92853 200682 142155
rect 201358 92989 201418 186899
rect 201355 92988 201421 92989
rect 201355 92924 201356 92988
rect 201420 92924 201421 92988
rect 201355 92923 201421 92924
rect 201542 92853 201602 223483
rect 203195 205732 203261 205733
rect 203195 205668 203196 205732
rect 203260 205668 203261 205732
rect 203195 205667 203261 205668
rect 203198 202877 203258 205667
rect 203514 205174 204134 239592
rect 203514 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 204134 205174
rect 203514 204854 204134 204938
rect 204854 204917 204914 300867
rect 203514 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 204134 204854
rect 204851 204916 204917 204917
rect 204851 204852 204852 204916
rect 204916 204852 204917 204916
rect 204851 204851 204917 204852
rect 203195 202876 203261 202877
rect 203195 202812 203196 202876
rect 203260 202812 203261 202876
rect 203195 202811 203261 202812
rect 200619 92852 200685 92853
rect 200619 92788 200620 92852
rect 200684 92788 200685 92852
rect 200619 92787 200685 92788
rect 201539 92852 201605 92853
rect 201539 92788 201540 92852
rect 201604 92788 201605 92852
rect 201539 92787 201605 92788
rect 203198 92445 203258 202811
rect 203514 169174 204134 204618
rect 205774 199341 205834 300867
rect 207062 206277 207122 300867
rect 208531 300796 208597 300797
rect 208531 300732 208532 300796
rect 208596 300732 208597 300796
rect 208531 300731 208597 300732
rect 207234 208894 207854 239592
rect 207234 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 207854 208894
rect 207234 208574 207854 208658
rect 207234 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 207854 208574
rect 207059 206276 207125 206277
rect 207059 206212 207060 206276
rect 207124 206212 207125 206276
rect 207059 206211 207125 206212
rect 205771 199340 205837 199341
rect 205771 199276 205772 199340
rect 205836 199276 205837 199340
rect 205771 199275 205837 199276
rect 204851 194036 204917 194037
rect 204851 193972 204852 194036
rect 204916 193972 204917 194036
rect 204851 193971 204917 193972
rect 203514 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 204134 169174
rect 203514 168854 204134 168938
rect 203514 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 204134 168854
rect 203514 143035 204134 168618
rect 204264 129454 204584 129486
rect 204264 129218 204306 129454
rect 204542 129218 204584 129454
rect 204264 129134 204584 129218
rect 204264 128898 204306 129134
rect 204542 128898 204584 129134
rect 204264 128866 204584 128898
rect 204854 92717 204914 193971
rect 207059 173908 207125 173909
rect 207059 173844 207060 173908
rect 207124 173844 207125 173908
rect 207059 173843 207125 173844
rect 207062 92853 207122 173843
rect 207234 172894 207854 208338
rect 208534 193901 208594 300731
rect 210374 300661 210434 320179
rect 210954 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 211574 320294
rect 210954 303592 211574 320058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 213683 303652 213749 303653
rect 213683 303588 213684 303652
rect 213748 303588 213749 303652
rect 217794 303592 218414 326898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 547174 222134 582618
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 511174 222134 546618
rect 221514 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 222134 511174
rect 221514 510854 222134 510938
rect 221514 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 222134 510854
rect 221514 475174 222134 510618
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 221514 439174 222134 474618
rect 221514 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 222134 439174
rect 221514 438854 222134 438938
rect 221514 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 222134 438854
rect 221514 403174 222134 438618
rect 221514 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 222134 403174
rect 221514 402854 222134 402938
rect 221514 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 222134 402854
rect 221514 367174 222134 402618
rect 221514 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 222134 367174
rect 221514 366854 222134 366938
rect 221514 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 222134 366854
rect 221514 331174 222134 366618
rect 221514 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 222134 331174
rect 221514 330854 222134 330938
rect 221514 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 222134 330854
rect 219939 303652 220005 303653
rect 213683 303587 213749 303588
rect 219939 303588 219940 303652
rect 220004 303588 220005 303652
rect 221514 303592 222134 330618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 550894 225854 586338
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 514894 225854 550338
rect 225234 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 225854 514894
rect 225234 514574 225854 514658
rect 225234 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 225854 514574
rect 225234 478894 225854 514338
rect 225234 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 225854 478894
rect 225234 478574 225854 478658
rect 225234 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 225854 478574
rect 225234 442894 225854 478338
rect 225234 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 225854 442894
rect 225234 442574 225854 442658
rect 225234 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 225854 442574
rect 225234 406894 225854 442338
rect 225234 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 225854 406894
rect 225234 406574 225854 406658
rect 225234 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 225854 406574
rect 225234 370894 225854 406338
rect 225234 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 225854 370894
rect 225234 370574 225854 370658
rect 225234 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 225854 370574
rect 225234 334894 225854 370338
rect 225234 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 225854 334894
rect 225234 334574 225854 334658
rect 225234 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 225854 334574
rect 225234 303592 225854 334338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 554614 229574 590058
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 518614 229574 554058
rect 228954 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 229574 518614
rect 228954 518294 229574 518378
rect 228954 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 229574 518294
rect 228954 482614 229574 518058
rect 228954 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 229574 482614
rect 228954 482294 229574 482378
rect 228954 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 229574 482294
rect 228954 446614 229574 482058
rect 228954 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 229574 446614
rect 228954 446294 229574 446378
rect 228954 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 229574 446294
rect 228954 410614 229574 446058
rect 228954 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 229574 410614
rect 228954 410294 229574 410378
rect 228954 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 229574 410294
rect 228954 374614 229574 410058
rect 228954 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 229574 374614
rect 228954 374294 229574 374378
rect 228954 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 229574 374294
rect 228954 338614 229574 374058
rect 228954 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 229574 338614
rect 228954 338294 229574 338378
rect 228954 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 229574 338294
rect 228954 303592 229574 338058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 601174 240134 636618
rect 239514 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 240134 601174
rect 239514 600854 240134 600938
rect 239514 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 240134 600854
rect 239514 565174 240134 600618
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 239514 529174 240134 564618
rect 239514 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 240134 529174
rect 239514 528854 240134 528938
rect 239514 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 240134 528854
rect 239514 493174 240134 528618
rect 239514 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 240134 493174
rect 239514 492854 240134 492938
rect 239514 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 240134 492854
rect 239514 457174 240134 492618
rect 239514 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 240134 457174
rect 239514 456854 240134 456938
rect 239514 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 240134 456854
rect 239514 421174 240134 456618
rect 239514 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 240134 421174
rect 239514 420854 240134 420938
rect 239514 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 240134 420854
rect 239514 385174 240134 420618
rect 239514 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 240134 385174
rect 239514 384854 240134 384938
rect 239514 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 240134 384854
rect 239514 349174 240134 384618
rect 239514 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 240134 349174
rect 239514 348854 240134 348938
rect 239514 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 240134 348854
rect 237971 335476 238037 335477
rect 237971 335412 237972 335476
rect 238036 335412 238037 335476
rect 237971 335411 238037 335412
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 303592 236414 308898
rect 237974 303653 238034 335411
rect 239514 313174 240134 348618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 604894 243854 640338
rect 243234 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 243854 604894
rect 243234 604574 243854 604658
rect 243234 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 243854 604574
rect 243234 568894 243854 604338
rect 243234 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 243854 568894
rect 243234 568574 243854 568658
rect 243234 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 243854 568574
rect 243234 532894 243854 568338
rect 243234 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 243854 532894
rect 243234 532574 243854 532658
rect 243234 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 243854 532574
rect 243234 496894 243854 532338
rect 243234 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 243854 496894
rect 243234 496574 243854 496658
rect 243234 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 243854 496574
rect 243234 460894 243854 496338
rect 243234 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 243854 460894
rect 243234 460574 243854 460658
rect 243234 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 243854 460574
rect 243234 424894 243854 460338
rect 243234 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 243854 424894
rect 243234 424574 243854 424658
rect 243234 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 243854 424574
rect 243234 388894 243854 424338
rect 243234 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 243854 388894
rect 243234 388574 243854 388658
rect 243234 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 243854 388574
rect 243234 352894 243854 388338
rect 243234 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 243854 352894
rect 243234 352574 243854 352658
rect 243234 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 243854 352574
rect 242019 329900 242085 329901
rect 242019 329836 242020 329900
rect 242084 329836 242085 329900
rect 242019 329835 242085 329836
rect 239514 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 240134 313174
rect 239514 312854 240134 312938
rect 239514 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 240134 312854
rect 239259 303924 239325 303925
rect 239259 303860 239260 303924
rect 239324 303860 239325 303924
rect 239259 303859 239325 303860
rect 237971 303652 238037 303653
rect 219939 303587 220005 303588
rect 237971 303588 237972 303652
rect 238036 303588 238037 303652
rect 237971 303587 238037 303588
rect 212395 301204 212461 301205
rect 212395 301140 212396 301204
rect 212460 301140 212461 301204
rect 212395 301139 212461 301140
rect 210371 300660 210437 300661
rect 210371 300596 210372 300660
rect 210436 300596 210437 300660
rect 210371 300595 210437 300596
rect 210374 235925 210434 300595
rect 210371 235924 210437 235925
rect 210371 235860 210372 235924
rect 210436 235860 210437 235924
rect 210371 235859 210437 235860
rect 209819 233204 209885 233205
rect 209819 233140 209820 233204
rect 209884 233140 209885 233204
rect 209819 233139 209885 233140
rect 208715 227764 208781 227765
rect 208715 227700 208716 227764
rect 208780 227700 208781 227764
rect 208715 227699 208781 227700
rect 208531 193900 208597 193901
rect 208531 193836 208532 193900
rect 208596 193836 208597 193900
rect 208531 193835 208597 193836
rect 207234 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 207854 172894
rect 207234 172574 207854 172658
rect 207234 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 207854 172574
rect 207234 143035 207854 172338
rect 208718 92853 208778 227699
rect 209140 111454 209460 111486
rect 209140 111218 209182 111454
rect 209418 111218 209460 111454
rect 209140 111134 209460 111218
rect 209140 110898 209182 111134
rect 209418 110898 209460 111134
rect 209140 110866 209460 110898
rect 209822 92853 209882 233139
rect 210954 212614 211574 239592
rect 210954 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 211574 212614
rect 210954 212294 211574 212378
rect 210954 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 211574 212294
rect 210954 176614 211574 212058
rect 210954 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 211574 176614
rect 210954 176294 211574 176378
rect 210954 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 211574 176294
rect 210954 143035 211574 176058
rect 212398 160717 212458 301139
rect 213136 273454 213456 273486
rect 213136 273218 213178 273454
rect 213414 273218 213456 273454
rect 213136 273134 213456 273218
rect 213136 272898 213178 273134
rect 213414 272898 213456 273134
rect 213136 272866 213456 272898
rect 212395 160716 212461 160717
rect 212395 160652 212396 160716
rect 212460 160652 212461 160716
rect 212395 160651 212461 160652
rect 213686 155277 213746 303587
rect 215891 301068 215957 301069
rect 215891 301004 215892 301068
rect 215956 301004 215957 301068
rect 215891 301003 215957 301004
rect 218651 301068 218717 301069
rect 218651 301004 218652 301068
rect 218716 301004 218717 301068
rect 218651 301003 218717 301004
rect 214419 300932 214485 300933
rect 214419 300868 214420 300932
rect 214484 300868 214485 300932
rect 214419 300867 214485 300868
rect 214422 203557 214482 300867
rect 215339 240140 215405 240141
rect 215339 240076 215340 240140
rect 215404 240076 215405 240140
rect 215339 240075 215405 240076
rect 215342 239869 215402 240075
rect 215339 239868 215405 239869
rect 215339 239804 215340 239868
rect 215404 239804 215405 239868
rect 215339 239803 215405 239804
rect 214419 203556 214485 203557
rect 214419 203492 214420 203556
rect 214484 203492 214485 203556
rect 214419 203491 214485 203492
rect 213683 155276 213749 155277
rect 213683 155212 213684 155276
rect 213748 155212 213749 155276
rect 213683 155211 213749 155212
rect 213683 148476 213749 148477
rect 213683 148412 213684 148476
rect 213748 148412 213749 148476
rect 213683 148411 213749 148412
rect 213686 92853 213746 148411
rect 214016 129454 214336 129486
rect 214016 129218 214058 129454
rect 214294 129218 214336 129454
rect 214016 129134 214336 129218
rect 214016 128898 214058 129134
rect 214294 128898 214336 129134
rect 214016 128866 214336 128898
rect 215342 93397 215402 239803
rect 215894 216069 215954 301003
rect 217179 300932 217245 300933
rect 217179 300868 217180 300932
rect 217244 300868 217245 300932
rect 217179 300867 217245 300868
rect 217182 220149 217242 300867
rect 217179 220148 217245 220149
rect 217179 220084 217180 220148
rect 217244 220084 217245 220148
rect 217179 220083 217245 220084
rect 217794 219454 218414 239592
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 215891 216068 215957 216069
rect 215891 216004 215892 216068
rect 215956 216004 215957 216068
rect 215891 216003 215957 216004
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 147454 218414 182898
rect 218654 178669 218714 301003
rect 219203 300932 219269 300933
rect 219203 300868 219204 300932
rect 219268 300868 219269 300932
rect 219203 300867 219269 300868
rect 218651 178668 218717 178669
rect 218651 178604 218652 178668
rect 218716 178604 218717 178668
rect 218651 178603 218717 178604
rect 219206 147690 219266 300867
rect 219942 210357 220002 303587
rect 224171 301340 224237 301341
rect 224171 301276 224172 301340
rect 224236 301276 224237 301340
rect 224171 301275 224237 301276
rect 233187 301340 233253 301341
rect 233187 301276 233188 301340
rect 233252 301276 233253 301340
rect 233187 301275 233253 301276
rect 234659 301340 234725 301341
rect 234659 301276 234660 301340
rect 234724 301276 234725 301340
rect 234659 301275 234725 301276
rect 236499 301340 236565 301341
rect 236499 301276 236500 301340
rect 236564 301276 236565 301340
rect 236499 301275 236565 301276
rect 220859 300932 220925 300933
rect 220859 300868 220860 300932
rect 220924 300868 220925 300932
rect 220859 300867 220925 300868
rect 222331 300932 222397 300933
rect 222331 300868 222332 300932
rect 222396 300868 222397 300932
rect 222331 300867 222397 300868
rect 220862 226949 220922 300867
rect 220859 226948 220925 226949
rect 220859 226884 220860 226948
rect 220924 226884 220925 226948
rect 220859 226883 220925 226884
rect 221514 223174 222134 239592
rect 221514 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 222134 223174
rect 221514 222854 222134 222938
rect 221514 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 222134 222854
rect 219939 210356 220005 210357
rect 219939 210292 219940 210356
rect 220004 210292 220005 210356
rect 219939 210291 220005 210292
rect 221514 187174 222134 222618
rect 222334 211853 222394 300867
rect 223619 227084 223685 227085
rect 223619 227020 223620 227084
rect 223684 227020 223685 227084
rect 223619 227019 223685 227020
rect 222331 211852 222397 211853
rect 222331 211788 222332 211852
rect 222396 211788 222397 211852
rect 222331 211787 222397 211788
rect 221514 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 222134 187174
rect 221514 186854 222134 186938
rect 221514 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 222134 186854
rect 221514 151174 222134 186618
rect 221514 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 222134 151174
rect 221514 150854 222134 150938
rect 221514 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 222134 150854
rect 219206 147630 219450 147690
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 143035 218414 146898
rect 219390 145757 219450 147630
rect 219387 145756 219453 145757
rect 219387 145692 219388 145756
rect 219452 145692 219453 145756
rect 219387 145691 219453 145692
rect 221514 143035 222134 150618
rect 223622 132510 223682 227019
rect 224174 222869 224234 301275
rect 224355 300932 224421 300933
rect 224355 300868 224356 300932
rect 224420 300868 224421 300932
rect 224355 300867 224421 300868
rect 226011 300932 226077 300933
rect 226011 300868 226012 300932
rect 226076 300868 226077 300932
rect 226011 300867 226077 300868
rect 226563 300932 226629 300933
rect 226563 300868 226564 300932
rect 226628 300868 226629 300932
rect 226563 300867 226629 300868
rect 226747 300932 226813 300933
rect 226747 300868 226748 300932
rect 226812 300868 226813 300932
rect 226747 300867 226813 300868
rect 229691 300932 229757 300933
rect 229691 300868 229692 300932
rect 229756 300868 229757 300932
rect 229691 300867 229757 300868
rect 230427 300932 230493 300933
rect 230427 300868 230428 300932
rect 230492 300868 230493 300932
rect 230427 300867 230493 300868
rect 230795 300932 230861 300933
rect 230795 300868 230796 300932
rect 230860 300868 230861 300932
rect 230795 300867 230861 300868
rect 232083 300932 232149 300933
rect 232083 300868 232084 300932
rect 232148 300868 232149 300932
rect 232083 300867 232149 300868
rect 232267 300932 232333 300933
rect 232267 300868 232268 300932
rect 232332 300868 232333 300932
rect 232267 300867 232333 300868
rect 224358 226541 224418 300867
rect 225234 226894 225854 239592
rect 225234 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 225854 226894
rect 225234 226574 225854 226658
rect 224355 226540 224421 226541
rect 224355 226476 224356 226540
rect 224420 226476 224421 226540
rect 224355 226475 224421 226476
rect 225234 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 225854 226574
rect 224171 222868 224237 222869
rect 224171 222804 224172 222868
rect 224236 222804 224237 222868
rect 224171 222803 224237 222804
rect 224907 207636 224973 207637
rect 224907 207572 224908 207636
rect 224972 207572 224973 207636
rect 224907 207571 224973 207572
rect 224910 147690 224970 207571
rect 224726 147630 224970 147690
rect 225234 190894 225854 226338
rect 226014 207093 226074 300867
rect 226566 218653 226626 300867
rect 226563 218652 226629 218653
rect 226563 218588 226564 218652
rect 226628 218588 226629 218652
rect 226563 218587 226629 218588
rect 226750 217293 226810 300867
rect 228496 291454 228816 291486
rect 228496 291218 228538 291454
rect 228774 291218 228816 291454
rect 228496 291134 228816 291218
rect 228496 290898 228538 291134
rect 228774 290898 228816 291134
rect 228496 290866 228816 290898
rect 228496 255454 228816 255486
rect 228496 255218 228538 255454
rect 228774 255218 228816 255454
rect 228496 255134 228816 255218
rect 228496 254898 228538 255134
rect 228774 254898 228816 255134
rect 228496 254866 228816 254898
rect 228219 234428 228285 234429
rect 228219 234364 228220 234428
rect 228284 234364 228285 234428
rect 228219 234363 228285 234364
rect 226747 217292 226813 217293
rect 226747 217228 226748 217292
rect 226812 217228 226813 217292
rect 226747 217227 226813 217228
rect 226011 207092 226077 207093
rect 226011 207028 226012 207092
rect 226076 207028 226077 207092
rect 226011 207027 226077 207028
rect 225234 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 225854 190894
rect 225234 190574 225854 190658
rect 225234 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 225854 190574
rect 225234 154894 225854 190338
rect 227667 164252 227733 164253
rect 227667 164188 227668 164252
rect 227732 164188 227733 164252
rect 227667 164187 227733 164188
rect 227670 162893 227730 164187
rect 227667 162892 227733 162893
rect 227667 162828 227668 162892
rect 227732 162828 227733 162892
rect 227667 162827 227733 162828
rect 225234 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 225854 154894
rect 226379 154732 226445 154733
rect 226379 154668 226380 154732
rect 226444 154668 226445 154732
rect 226379 154667 226445 154668
rect 225234 154574 225854 154658
rect 225234 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 225854 154574
rect 224355 142084 224421 142085
rect 224355 142020 224356 142084
rect 224420 142020 224421 142084
rect 224355 142019 224421 142020
rect 224358 136645 224418 142019
rect 224726 138030 224786 147630
rect 225234 143035 225854 154338
rect 224726 137970 224970 138030
rect 224355 136644 224421 136645
rect 224355 136580 224356 136644
rect 224420 136580 224421 136644
rect 224355 136579 224421 136580
rect 223622 132450 224418 132510
rect 224358 114477 224418 132450
rect 224355 114476 224421 114477
rect 224355 114412 224356 114476
rect 224420 114412 224421 114476
rect 224355 114411 224421 114412
rect 218892 111454 219212 111486
rect 218892 111218 218934 111454
rect 219170 111218 219212 111454
rect 218892 111134 219212 111218
rect 218892 110898 218934 111134
rect 219170 110898 219212 111134
rect 218892 110866 219212 110898
rect 224355 94348 224421 94349
rect 224355 94284 224356 94348
rect 224420 94284 224421 94348
rect 224355 94283 224421 94284
rect 215339 93396 215405 93397
rect 215339 93332 215340 93396
rect 215404 93332 215405 93396
rect 215339 93331 215405 93332
rect 207059 92852 207125 92853
rect 207059 92788 207060 92852
rect 207124 92788 207125 92852
rect 207059 92787 207125 92788
rect 208715 92852 208781 92853
rect 208715 92788 208716 92852
rect 208780 92788 208781 92852
rect 208715 92787 208781 92788
rect 209819 92852 209885 92853
rect 209819 92788 209820 92852
rect 209884 92788 209885 92852
rect 209819 92787 209885 92788
rect 213683 92852 213749 92853
rect 213683 92788 213684 92852
rect 213748 92788 213749 92852
rect 213683 92787 213749 92788
rect 204851 92716 204917 92717
rect 204851 92652 204852 92716
rect 204916 92652 204917 92716
rect 204851 92651 204917 92652
rect 203195 92444 203261 92445
rect 203195 92380 203196 92444
rect 203260 92380 203261 92444
rect 203195 92379 203261 92380
rect 224358 92173 224418 94283
rect 224910 93397 224970 137970
rect 226382 130117 226442 154667
rect 227670 139093 227730 162827
rect 228222 154597 228282 234363
rect 228954 230614 229574 239592
rect 228954 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 229574 230614
rect 228954 230294 229574 230378
rect 228954 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 229574 230294
rect 228954 194614 229574 230058
rect 228954 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 229574 194614
rect 228954 194294 229574 194378
rect 228954 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 229574 194294
rect 228954 158614 229574 194058
rect 229694 184245 229754 300867
rect 229691 184244 229757 184245
rect 229691 184180 229692 184244
rect 229756 184180 229757 184244
rect 229691 184179 229757 184180
rect 228954 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 229574 158614
rect 228954 158294 229574 158378
rect 228954 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 229574 158294
rect 228219 154596 228285 154597
rect 228219 154532 228220 154596
rect 228284 154532 228285 154596
rect 228219 154531 228285 154532
rect 228222 142170 228282 154531
rect 227854 142110 228282 142170
rect 227667 139092 227733 139093
rect 227667 139028 227668 139092
rect 227732 139028 227733 139092
rect 227667 139027 227733 139028
rect 227854 136645 227914 142110
rect 226931 136644 226997 136645
rect 226931 136580 226932 136644
rect 226996 136580 226997 136644
rect 226931 136579 226997 136580
rect 227851 136644 227917 136645
rect 227851 136580 227852 136644
rect 227916 136580 227917 136644
rect 227851 136579 227917 136580
rect 226379 130116 226445 130117
rect 226379 130052 226380 130116
rect 226444 130052 226445 130116
rect 226379 130051 226445 130052
rect 226934 121141 226994 136579
rect 228954 122614 229574 158058
rect 228954 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 229574 122614
rect 228954 122294 229574 122378
rect 228954 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 229574 122294
rect 226931 121140 226997 121141
rect 226931 121076 226932 121140
rect 226996 121076 226997 121140
rect 226931 121075 226997 121076
rect 225091 98292 225157 98293
rect 225091 98228 225092 98292
rect 225156 98228 225157 98292
rect 225091 98227 225157 98228
rect 224907 93396 224973 93397
rect 224907 93332 224908 93396
rect 224972 93332 224973 93396
rect 224907 93331 224973 93332
rect 224355 92172 224421 92173
rect 224355 92108 224356 92172
rect 224420 92108 224421 92172
rect 224355 92107 224421 92108
rect 199794 57454 200414 90782
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 197123 24172 197189 24173
rect 197123 24108 197124 24172
rect 197188 24108 197189 24172
rect 197123 24107 197189 24108
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 61174 204134 90782
rect 203514 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 204134 61174
rect 203514 60854 204134 60938
rect 203514 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 204134 60854
rect 203514 25174 204134 60618
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 64894 207854 90782
rect 207234 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 207854 64894
rect 207234 64574 207854 64658
rect 207234 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 207854 64574
rect 207234 28894 207854 64338
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 68614 211574 90782
rect 210954 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 211574 68614
rect 210954 68294 211574 68378
rect 210954 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 211574 68294
rect 210954 32614 211574 68058
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 75454 218414 90782
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 79174 222134 90782
rect 225094 84210 225154 98227
rect 226379 97204 226445 97205
rect 226379 97140 226380 97204
rect 226444 97140 226445 97204
rect 226379 97139 226445 97140
rect 224910 84150 225154 84210
rect 224910 80069 224970 84150
rect 225234 82894 225854 90782
rect 226382 85373 226442 97139
rect 226563 95300 226629 95301
rect 226563 95236 226564 95300
rect 226628 95236 226629 95300
rect 226563 95235 226629 95236
rect 226566 92445 226626 95235
rect 226563 92444 226629 92445
rect 226563 92380 226564 92444
rect 226628 92380 226629 92444
rect 226563 92379 226629 92380
rect 228954 86614 229574 122058
rect 228954 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 229574 86614
rect 228954 86294 229574 86378
rect 228954 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 229574 86294
rect 226379 85372 226445 85373
rect 226379 85308 226380 85372
rect 226444 85308 226445 85372
rect 226379 85307 226445 85308
rect 225234 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 225854 82894
rect 225234 82574 225854 82658
rect 225234 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 225854 82574
rect 224907 80068 224973 80069
rect 224907 80004 224908 80068
rect 224972 80004 224973 80068
rect 224907 80003 224973 80004
rect 221514 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 222134 79174
rect 221514 78854 222134 78938
rect 221514 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 222134 78854
rect 221514 43174 222134 78618
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 46894 225854 82338
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 50614 229574 86058
rect 230430 61437 230490 300867
rect 230427 61436 230493 61437
rect 230427 61372 230428 61436
rect 230492 61372 230493 61436
rect 230427 61371 230493 61372
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 230798 14517 230858 300867
rect 232086 196757 232146 300867
rect 232083 196756 232149 196757
rect 232083 196692 232084 196756
rect 232148 196692 232149 196756
rect 232083 196691 232149 196692
rect 232270 15877 232330 300867
rect 233190 17237 233250 301275
rect 233371 300932 233437 300933
rect 233371 300868 233372 300932
rect 233436 300868 233437 300932
rect 233371 300867 233437 300868
rect 233374 62797 233434 300867
rect 233371 62796 233437 62797
rect 233371 62732 233372 62796
rect 233436 62732 233437 62796
rect 233371 62731 233437 62732
rect 234662 55861 234722 301275
rect 234843 300932 234909 300933
rect 234843 300868 234844 300932
rect 234908 300868 234909 300932
rect 234843 300867 234909 300868
rect 234846 240141 234906 300867
rect 234843 240140 234909 240141
rect 234843 240076 234844 240140
rect 234908 240076 234909 240140
rect 234843 240075 234909 240076
rect 235794 237454 236414 239592
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 235794 201454 236414 236898
rect 236502 213213 236562 301275
rect 236683 300932 236749 300933
rect 236683 300868 236684 300932
rect 236748 300868 236749 300932
rect 236683 300867 236749 300868
rect 236686 240141 236746 300867
rect 236683 240140 236749 240141
rect 236683 240076 236684 240140
rect 236748 240076 236749 240140
rect 236683 240075 236749 240076
rect 236499 213212 236565 213213
rect 236499 213148 236500 213212
rect 236564 213148 236565 213212
rect 236499 213147 236565 213148
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 165454 236414 200898
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 235794 129454 236414 164898
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 237974 113117 238034 303587
rect 238155 301340 238221 301341
rect 238155 301276 238156 301340
rect 238220 301276 238221 301340
rect 238155 301275 238221 301276
rect 238158 214573 238218 301275
rect 238707 300932 238773 300933
rect 238707 300930 238708 300932
rect 238526 300870 238708 300930
rect 238526 238770 238586 300870
rect 238707 300868 238708 300870
rect 238772 300868 238773 300932
rect 238707 300867 238773 300868
rect 238707 238780 238773 238781
rect 238707 238770 238708 238780
rect 238526 238716 238708 238770
rect 238772 238716 238773 238780
rect 238526 238715 238773 238716
rect 238526 238710 238770 238715
rect 238155 214572 238221 214573
rect 238155 214508 238156 214572
rect 238220 214508 238221 214572
rect 238155 214507 238221 214508
rect 239262 173229 239322 303859
rect 239514 303592 240134 312618
rect 242022 303653 242082 329835
rect 243234 316894 243854 352338
rect 243234 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 243854 316894
rect 243234 316574 243854 316658
rect 243234 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 243854 316574
rect 240731 303652 240797 303653
rect 240731 303588 240732 303652
rect 240796 303588 240797 303652
rect 240731 303587 240797 303588
rect 242019 303652 242085 303653
rect 242019 303588 242020 303652
rect 242084 303588 242085 303652
rect 243234 303592 243854 316338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 608614 247574 644058
rect 246954 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 247574 608614
rect 246954 608294 247574 608378
rect 246954 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 247574 608294
rect 246954 572614 247574 608058
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 536614 247574 572058
rect 246954 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 247574 536614
rect 246954 536294 247574 536378
rect 246954 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 247574 536294
rect 246954 500614 247574 536058
rect 246954 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 247574 500614
rect 246954 500294 247574 500378
rect 246954 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 247574 500294
rect 246954 464614 247574 500058
rect 246954 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 247574 464614
rect 246954 464294 247574 464378
rect 246954 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 247574 464294
rect 246954 428614 247574 464058
rect 246954 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 247574 428614
rect 246954 428294 247574 428378
rect 246954 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 247574 428294
rect 246954 392614 247574 428058
rect 246954 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 247574 392614
rect 246954 392294 247574 392378
rect 246954 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 247574 392294
rect 246954 356614 247574 392058
rect 246954 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 247574 356614
rect 246954 356294 247574 356378
rect 246954 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 247574 356294
rect 246954 320614 247574 356058
rect 246954 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 247574 320614
rect 246954 320294 247574 320378
rect 246954 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 247574 320294
rect 246954 303592 247574 320058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253059 318204 253125 318205
rect 253059 318140 253060 318204
rect 253124 318140 253125 318204
rect 253059 318139 253125 318140
rect 253062 306390 253122 318139
rect 253062 306330 253674 306390
rect 242019 303587 242085 303588
rect 239514 205174 240134 239592
rect 239514 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 240134 205174
rect 239514 204854 240134 204938
rect 239514 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 240134 204854
rect 239259 173228 239325 173229
rect 239259 173164 239260 173228
rect 239324 173164 239325 173228
rect 239259 173163 239325 173164
rect 239514 169174 240134 204618
rect 239514 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 240134 169174
rect 239514 168854 240134 168938
rect 239514 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 240134 168854
rect 239514 133174 240134 168618
rect 239514 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 240134 133174
rect 239514 132854 240134 132938
rect 239514 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 240134 132854
rect 237971 113116 238037 113117
rect 237971 113052 237972 113116
rect 238036 113052 238037 113116
rect 237971 113051 238037 113052
rect 237974 111893 238034 113051
rect 237971 111892 238037 111893
rect 237971 111828 237972 111892
rect 238036 111828 238037 111892
rect 237971 111827 238037 111828
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 234659 55860 234725 55861
rect 234659 55796 234660 55860
rect 234724 55796 234725 55860
rect 234659 55795 234725 55796
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 233187 17236 233253 17237
rect 233187 17172 233188 17236
rect 233252 17172 233253 17236
rect 233187 17171 233253 17172
rect 232267 15876 232333 15877
rect 232267 15812 232268 15876
rect 232332 15812 232333 15876
rect 232267 15811 232333 15812
rect 230795 14516 230861 14517
rect 230795 14452 230796 14516
rect 230860 14452 230861 14516
rect 230795 14451 230861 14452
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 97174 240134 132618
rect 240734 111893 240794 303587
rect 240915 300932 240981 300933
rect 240915 300868 240916 300932
rect 240980 300868 240981 300932
rect 240915 300867 240981 300868
rect 241651 300932 241717 300933
rect 241651 300868 241652 300932
rect 241716 300868 241717 300932
rect 241651 300867 241717 300868
rect 240918 186965 240978 300867
rect 240915 186964 240981 186965
rect 240915 186900 240916 186964
rect 240980 186900 240981 186964
rect 240915 186899 240981 186900
rect 241654 171733 241714 300867
rect 242022 238101 242082 303587
rect 242939 300932 243005 300933
rect 242939 300868 242940 300932
rect 243004 300868 243005 300932
rect 242939 300867 243005 300868
rect 244411 300932 244477 300933
rect 244411 300868 244412 300932
rect 244476 300868 244477 300932
rect 244411 300867 244477 300868
rect 245699 300932 245765 300933
rect 245699 300868 245700 300932
rect 245764 300868 245765 300932
rect 245699 300867 245765 300868
rect 247723 300932 247789 300933
rect 247723 300868 247724 300932
rect 247788 300868 247789 300932
rect 247723 300867 247789 300868
rect 248459 300932 248525 300933
rect 248459 300868 248460 300932
rect 248524 300868 248525 300932
rect 248459 300867 248525 300868
rect 251219 300932 251285 300933
rect 251219 300868 251220 300932
rect 251284 300868 251285 300932
rect 251219 300867 251285 300868
rect 252507 300932 252573 300933
rect 252507 300868 252508 300932
rect 252572 300868 252573 300932
rect 252507 300867 252573 300868
rect 242019 238100 242085 238101
rect 242019 238036 242020 238100
rect 242084 238036 242085 238100
rect 242019 238035 242085 238036
rect 241651 171732 241717 171733
rect 241651 171668 241652 171732
rect 241716 171668 241717 171732
rect 241651 171667 241717 171668
rect 242942 148341 243002 300867
rect 243856 273454 244176 273486
rect 243856 273218 243898 273454
rect 244134 273218 244176 273454
rect 243856 273134 244176 273218
rect 243856 272898 243898 273134
rect 244134 272898 244176 273134
rect 243856 272866 244176 272898
rect 243234 208894 243854 239592
rect 243234 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 243854 208894
rect 243234 208574 243854 208658
rect 243234 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 243854 208574
rect 243234 172894 243854 208338
rect 243234 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 243854 172894
rect 243234 172574 243854 172658
rect 243234 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 243854 172574
rect 242939 148340 243005 148341
rect 242939 148276 242940 148340
rect 243004 148276 243005 148340
rect 242939 148275 243005 148276
rect 243234 136894 243854 172338
rect 244414 147117 244474 300867
rect 245702 206277 245762 300867
rect 246954 212614 247574 239592
rect 246954 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 247574 212614
rect 246954 212294 247574 212378
rect 246954 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 247574 212294
rect 245699 206276 245765 206277
rect 245699 206212 245700 206276
rect 245764 206212 245765 206276
rect 245699 206211 245765 206212
rect 246954 176614 247574 212058
rect 247726 181389 247786 300867
rect 248462 213485 248522 300867
rect 248459 213484 248525 213485
rect 248459 213420 248460 213484
rect 248524 213420 248525 213484
rect 248459 213419 248525 213420
rect 251222 194037 251282 300867
rect 252510 248430 252570 300867
rect 253614 292773 253674 306330
rect 253794 303592 254414 326898
rect 257514 691174 258134 706202
rect 260051 699820 260117 699821
rect 260051 699756 260052 699820
rect 260116 699756 260117 699820
rect 260051 699755 260117 699756
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 547174 258134 582618
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257514 511174 258134 546618
rect 257514 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 258134 511174
rect 257514 510854 258134 510938
rect 257514 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 258134 510854
rect 257514 475174 258134 510618
rect 257514 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 258134 475174
rect 257514 474854 258134 474938
rect 257514 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 258134 474854
rect 257514 439174 258134 474618
rect 257514 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 258134 439174
rect 257514 438854 258134 438938
rect 257514 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 258134 438854
rect 257514 403174 258134 438618
rect 257514 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 258134 403174
rect 257514 402854 258134 402938
rect 257514 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 258134 402854
rect 257514 367174 258134 402618
rect 257514 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 258134 367174
rect 257514 366854 258134 366938
rect 257514 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 258134 366854
rect 257514 331174 258134 366618
rect 257514 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 258134 331174
rect 257514 330854 258134 330938
rect 257514 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 258134 330854
rect 254531 307052 254597 307053
rect 254531 306988 254532 307052
rect 254596 306988 254597 307052
rect 254531 306987 254597 306988
rect 254163 301748 254229 301749
rect 254163 301684 254164 301748
rect 254228 301684 254229 301748
rect 254163 301683 254229 301684
rect 254166 294269 254226 301683
rect 254534 299029 254594 306987
rect 255451 300388 255517 300389
rect 255451 300324 255452 300388
rect 255516 300324 255517 300388
rect 255451 300323 255517 300324
rect 255267 299572 255333 299573
rect 255267 299508 255268 299572
rect 255332 299508 255333 299572
rect 255267 299507 255333 299508
rect 254531 299028 254597 299029
rect 254531 298964 254532 299028
rect 254596 298964 254597 299028
rect 254531 298963 254597 298964
rect 255270 298621 255330 299507
rect 255454 298757 255514 300323
rect 256739 300252 256805 300253
rect 256739 300188 256740 300252
rect 256804 300188 256805 300252
rect 256739 300187 256805 300188
rect 256555 299436 256621 299437
rect 256555 299372 256556 299436
rect 256620 299372 256621 299436
rect 256555 299371 256621 299372
rect 255451 298756 255517 298757
rect 255451 298692 255452 298756
rect 255516 298692 255517 298756
rect 255451 298691 255517 298692
rect 255267 298620 255333 298621
rect 255267 298556 255268 298620
rect 255332 298556 255333 298620
rect 255267 298555 255333 298556
rect 254531 298212 254597 298213
rect 254531 298148 254532 298212
rect 254596 298148 254597 298212
rect 254531 298147 254597 298148
rect 254163 294268 254229 294269
rect 254163 294204 254164 294268
rect 254228 294204 254229 294268
rect 254163 294203 254229 294204
rect 253611 292772 253677 292773
rect 253611 292708 253612 292772
rect 253676 292708 253677 292772
rect 253611 292707 253677 292708
rect 252510 248370 252754 248430
rect 252694 244290 252754 248370
rect 252694 244230 253122 244290
rect 252875 243676 252941 243677
rect 252875 243612 252876 243676
rect 252940 243612 252941 243676
rect 252875 243611 252941 243612
rect 252878 242450 252938 243611
rect 252510 242390 252938 242450
rect 252510 239461 252570 242390
rect 252507 239460 252573 239461
rect 252507 239396 252508 239460
rect 252572 239396 252573 239460
rect 252507 239395 252573 239396
rect 253062 234630 253122 244230
rect 252510 234570 253122 234630
rect 251219 194036 251285 194037
rect 251219 193972 251220 194036
rect 251284 193972 251285 194036
rect 251219 193971 251285 193972
rect 247723 181388 247789 181389
rect 247723 181324 247724 181388
rect 247788 181324 247789 181388
rect 247723 181323 247789 181324
rect 246954 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 247574 176614
rect 246954 176294 247574 176378
rect 246954 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 247574 176294
rect 244411 147116 244477 147117
rect 244411 147052 244412 147116
rect 244476 147052 244477 147116
rect 244411 147051 244477 147052
rect 243234 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 243854 136894
rect 243234 136574 243854 136658
rect 243234 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 243854 136574
rect 240731 111892 240797 111893
rect 240731 111828 240732 111892
rect 240796 111828 240797 111892
rect 240731 111827 240797 111828
rect 239514 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 240134 97174
rect 239514 96854 240134 96938
rect 239514 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 240134 96854
rect 239514 61174 240134 96618
rect 239514 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 240134 61174
rect 239514 60854 240134 60938
rect 239514 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 240134 60854
rect 239514 25174 240134 60618
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 100894 243854 136338
rect 243234 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 243854 100894
rect 243234 100574 243854 100658
rect 243234 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 243854 100574
rect 243234 64894 243854 100338
rect 243234 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 243854 64894
rect 243234 64574 243854 64658
rect 243234 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 243854 64574
rect 243234 28894 243854 64338
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 140614 247574 176058
rect 252510 166293 252570 234570
rect 253794 219454 254414 239592
rect 254534 231165 254594 298147
rect 256558 294541 256618 299371
rect 256555 294540 256621 294541
rect 256555 294476 256556 294540
rect 256620 294476 256621 294540
rect 256555 294475 256621 294476
rect 256742 290733 256802 300187
rect 257514 295174 258134 330618
rect 258395 318340 258461 318341
rect 258395 318276 258396 318340
rect 258460 318276 258461 318340
rect 258395 318275 258461 318276
rect 258398 316050 258458 318275
rect 260054 318069 260114 699755
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 550894 261854 586338
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 514894 261854 550338
rect 261234 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 261854 514894
rect 261234 514574 261854 514658
rect 261234 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 261854 514574
rect 261234 478894 261854 514338
rect 261234 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 261854 478894
rect 261234 478574 261854 478658
rect 261234 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 261854 478574
rect 261234 442894 261854 478338
rect 261234 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 261854 442894
rect 261234 442574 261854 442658
rect 261234 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 261854 442574
rect 261234 406894 261854 442338
rect 261234 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 261854 406894
rect 261234 406574 261854 406658
rect 261234 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 261854 406574
rect 261234 370894 261854 406338
rect 261234 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 261854 370894
rect 261234 370574 261854 370658
rect 261234 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 261854 370574
rect 261234 334894 261854 370338
rect 261234 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 261854 334894
rect 261234 334574 261854 334658
rect 261234 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 261854 334574
rect 260051 318068 260117 318069
rect 260051 318004 260052 318068
rect 260116 318004 260117 318068
rect 260051 318003 260117 318004
rect 260054 316050 260114 318003
rect 257514 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 258134 295174
rect 257514 294854 258134 294938
rect 257514 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 258134 294854
rect 256739 290732 256805 290733
rect 256739 290668 256740 290732
rect 256804 290668 256805 290732
rect 256739 290667 256805 290668
rect 255451 261900 255517 261901
rect 255451 261836 255452 261900
rect 255516 261836 255517 261900
rect 255451 261835 255517 261836
rect 255267 260812 255333 260813
rect 255267 260748 255268 260812
rect 255332 260748 255333 260812
rect 255267 260747 255333 260748
rect 254715 253468 254781 253469
rect 254715 253404 254716 253468
rect 254780 253404 254781 253468
rect 254715 253403 254781 253404
rect 254718 240141 254778 253403
rect 254715 240140 254781 240141
rect 254715 240076 254716 240140
rect 254780 240076 254781 240140
rect 254715 240075 254781 240076
rect 254531 231164 254597 231165
rect 254531 231100 254532 231164
rect 254596 231100 254597 231164
rect 254531 231099 254597 231100
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 255270 213349 255330 260747
rect 255454 221509 255514 261835
rect 256739 260540 256805 260541
rect 256739 260476 256740 260540
rect 256804 260476 256805 260540
rect 256739 260475 256805 260476
rect 256742 239597 256802 260475
rect 257514 259174 258134 294618
rect 257514 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 258134 259174
rect 257514 258854 258134 258938
rect 257514 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 258134 258854
rect 256739 239596 256805 239597
rect 256739 239532 256740 239596
rect 256804 239532 256805 239596
rect 256739 239531 256805 239532
rect 257514 223174 258134 258618
rect 258214 315990 258458 316050
rect 259502 315990 260114 316050
rect 258214 258090 258274 315990
rect 258395 314940 258461 314941
rect 258395 314876 258396 314940
rect 258460 314876 258461 314940
rect 258395 314875 258461 314876
rect 258398 265301 258458 314875
rect 259502 267477 259562 315990
rect 261234 298894 261854 334338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 268331 702540 268397 702541
rect 268331 702476 268332 702540
rect 268396 702476 268397 702540
rect 268331 702475 268397 702476
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 554614 265574 590058
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 518614 265574 554058
rect 264954 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 265574 518614
rect 264954 518294 265574 518378
rect 264954 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 265574 518294
rect 264954 482614 265574 518058
rect 264954 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 265574 482614
rect 264954 482294 265574 482378
rect 264954 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 265574 482294
rect 264954 446614 265574 482058
rect 264954 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 265574 446614
rect 264954 446294 265574 446378
rect 264954 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 265574 446294
rect 264954 410614 265574 446058
rect 264954 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 265574 410614
rect 264954 410294 265574 410378
rect 264954 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 265574 410294
rect 264954 374614 265574 410058
rect 264954 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 265574 374614
rect 264954 374294 265574 374378
rect 264954 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 265574 374294
rect 264954 338614 265574 374058
rect 264954 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 265574 338614
rect 264954 338294 265574 338378
rect 264954 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 265574 338294
rect 262259 319428 262325 319429
rect 262259 319364 262260 319428
rect 262324 319364 262325 319428
rect 262259 319363 262325 319364
rect 261234 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 261854 298894
rect 261234 298574 261854 298658
rect 261234 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 261854 298574
rect 259499 267476 259565 267477
rect 259499 267412 259500 267476
rect 259564 267412 259565 267476
rect 259499 267411 259565 267412
rect 258395 265300 258461 265301
rect 258395 265236 258396 265300
rect 258460 265236 258461 265300
rect 258395 265235 258461 265236
rect 261234 262894 261854 298338
rect 261234 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 261854 262894
rect 261234 262574 261854 262658
rect 261234 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 261854 262574
rect 258214 258030 258458 258090
rect 258398 254829 258458 258030
rect 259499 257412 259565 257413
rect 259499 257348 259500 257412
rect 259564 257348 259565 257412
rect 259499 257347 259565 257348
rect 258395 254828 258461 254829
rect 258395 254764 258396 254828
rect 258460 254764 258461 254828
rect 258395 254763 258461 254764
rect 258395 247076 258461 247077
rect 258395 247012 258396 247076
rect 258460 247012 258461 247076
rect 258395 247011 258461 247012
rect 258398 240821 258458 247011
rect 258395 240820 258461 240821
rect 258395 240756 258396 240820
rect 258460 240756 258461 240820
rect 258395 240755 258461 240756
rect 259502 226269 259562 257347
rect 259683 248436 259749 248437
rect 259683 248372 259684 248436
rect 259748 248372 259749 248436
rect 259683 248371 259749 248372
rect 259686 244221 259746 248371
rect 259683 244220 259749 244221
rect 259683 244156 259684 244220
rect 259748 244156 259749 244220
rect 259683 244155 259749 244156
rect 259686 238781 259746 244155
rect 259683 238780 259749 238781
rect 259683 238716 259684 238780
rect 259748 238716 259749 238780
rect 259683 238715 259749 238716
rect 261234 226894 261854 262338
rect 262262 259861 262322 319363
rect 264954 302614 265574 338058
rect 264954 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 265574 302614
rect 264954 302294 265574 302378
rect 264954 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 265574 302294
rect 264954 266614 265574 302058
rect 264954 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 265574 266614
rect 264954 266294 265574 266378
rect 264954 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 265574 266294
rect 262259 259860 262325 259861
rect 262259 259796 262260 259860
rect 262324 259796 262325 259860
rect 262259 259795 262325 259796
rect 263547 258636 263613 258637
rect 263547 258572 263548 258636
rect 263612 258572 263613 258636
rect 263547 258571 263613 258572
rect 262259 258228 262325 258229
rect 262259 258164 262260 258228
rect 262324 258164 262325 258228
rect 262259 258163 262325 258164
rect 262262 238101 262322 258163
rect 262259 238100 262325 238101
rect 262259 238036 262260 238100
rect 262324 238036 262325 238100
rect 262259 238035 262325 238036
rect 261234 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 261854 226894
rect 261234 226574 261854 226658
rect 261234 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 261854 226574
rect 259499 226268 259565 226269
rect 259499 226204 259500 226268
rect 259564 226204 259565 226268
rect 259499 226203 259565 226204
rect 257514 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 258134 223174
rect 257514 222854 258134 222938
rect 257514 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 258134 222854
rect 255451 221508 255517 221509
rect 255451 221444 255452 221508
rect 255516 221444 255517 221508
rect 255451 221443 255517 221444
rect 255267 213348 255333 213349
rect 255267 213284 255268 213348
rect 255332 213284 255333 213348
rect 255267 213283 255333 213284
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 252507 166292 252573 166293
rect 252507 166228 252508 166292
rect 252572 166228 252573 166292
rect 252507 166227 252573 166228
rect 246954 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 247574 140614
rect 246954 140294 247574 140378
rect 246954 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 247574 140294
rect 246954 104614 247574 140058
rect 246954 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 247574 104614
rect 246954 104294 247574 104378
rect 246954 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 247574 104294
rect 246954 68614 247574 104058
rect 246954 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 247574 68614
rect 246954 68294 247574 68378
rect 246954 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 247574 68294
rect 246954 32614 247574 68058
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 187174 258134 222618
rect 257514 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 258134 187174
rect 257514 186854 258134 186938
rect 257514 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 258134 186854
rect 257514 151174 258134 186618
rect 257514 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 258134 151174
rect 257514 150854 258134 150938
rect 257514 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 258134 150854
rect 257514 115174 258134 150618
rect 257514 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 258134 115174
rect 257514 114854 258134 114938
rect 257514 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 258134 114854
rect 257514 79174 258134 114618
rect 257514 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 258134 79174
rect 257514 78854 258134 78938
rect 257514 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 258134 78854
rect 257514 43174 258134 78618
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 190894 261854 226338
rect 263550 220829 263610 258571
rect 264954 230614 265574 266058
rect 268334 265437 268394 702475
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 268331 265436 268397 265437
rect 268331 265372 268332 265436
rect 268396 265372 268397 265436
rect 268331 265371 268397 265372
rect 267779 257276 267845 257277
rect 267779 257212 267780 257276
rect 267844 257212 267845 257276
rect 267779 257211 267845 257212
rect 266307 254012 266373 254013
rect 266307 253948 266308 254012
rect 266372 253948 266373 254012
rect 266307 253947 266373 253948
rect 266310 235245 266370 253947
rect 266307 235244 266373 235245
rect 266307 235180 266308 235244
rect 266372 235180 266373 235244
rect 266307 235179 266373 235180
rect 267782 234429 267842 257211
rect 269067 255644 269133 255645
rect 269067 255580 269068 255644
rect 269132 255580 269133 255644
rect 269067 255579 269133 255580
rect 269070 235925 269130 255579
rect 271794 237454 272414 272898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 601174 276134 636618
rect 275514 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 276134 601174
rect 275514 600854 276134 600938
rect 275514 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 276134 600854
rect 275514 565174 276134 600618
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 529174 276134 564618
rect 275514 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 276134 529174
rect 275514 528854 276134 528938
rect 275514 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 276134 528854
rect 275514 493174 276134 528618
rect 275514 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 276134 493174
rect 275514 492854 276134 492938
rect 275514 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 276134 492854
rect 275514 457174 276134 492618
rect 275514 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 276134 457174
rect 275514 456854 276134 456938
rect 275514 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 276134 456854
rect 275514 421174 276134 456618
rect 275514 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 276134 421174
rect 275514 420854 276134 420938
rect 275514 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 276134 420854
rect 275514 385174 276134 420618
rect 275514 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 276134 385174
rect 275514 384854 276134 384938
rect 275514 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 276134 384854
rect 275514 349174 276134 384618
rect 275514 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 276134 349174
rect 275514 348854 276134 348938
rect 275514 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 276134 348854
rect 275514 313174 276134 348618
rect 275514 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 276134 313174
rect 275514 312854 276134 312938
rect 275514 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 276134 312854
rect 275514 277174 276134 312618
rect 275514 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 276134 277174
rect 275514 276854 276134 276938
rect 275514 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 276134 276854
rect 273299 254012 273365 254013
rect 273299 253948 273300 254012
rect 273364 253948 273365 254012
rect 273299 253947 273365 253948
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 269067 235924 269133 235925
rect 269067 235860 269068 235924
rect 269132 235860 269133 235924
rect 269067 235859 269133 235860
rect 267779 234428 267845 234429
rect 267779 234364 267780 234428
rect 267844 234364 267845 234428
rect 267779 234363 267845 234364
rect 264954 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 265574 230614
rect 264954 230294 265574 230378
rect 264954 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 265574 230294
rect 263547 220828 263613 220829
rect 263547 220764 263548 220828
rect 263612 220764 263613 220828
rect 263547 220763 263613 220764
rect 261234 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 261854 190894
rect 261234 190574 261854 190658
rect 261234 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 261854 190574
rect 261234 154894 261854 190338
rect 261234 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 261854 154894
rect 261234 154574 261854 154658
rect 261234 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 261854 154574
rect 261234 118894 261854 154338
rect 261234 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 261854 118894
rect 261234 118574 261854 118658
rect 261234 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 261854 118574
rect 261234 82894 261854 118338
rect 261234 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 261854 82894
rect 261234 82574 261854 82658
rect 261234 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 261854 82574
rect 261234 46894 261854 82338
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 194614 265574 230058
rect 264954 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 265574 194614
rect 264954 194294 265574 194378
rect 264954 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 265574 194294
rect 264954 158614 265574 194058
rect 264954 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 265574 158614
rect 264954 158294 265574 158378
rect 264954 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 265574 158294
rect 264954 122614 265574 158058
rect 264954 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 265574 122614
rect 264954 122294 265574 122378
rect 264954 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 265574 122294
rect 264954 86614 265574 122058
rect 264954 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 265574 86614
rect 264954 86294 265574 86378
rect 264954 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 265574 86294
rect 264954 50614 265574 86058
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 201454 272414 236898
rect 273302 226133 273362 253947
rect 275514 241174 276134 276618
rect 275514 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 276134 241174
rect 275514 240854 276134 240938
rect 275514 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 276134 240854
rect 273299 226132 273365 226133
rect 273299 226068 273300 226132
rect 273364 226068 273365 226132
rect 273299 226067 273365 226068
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 205174 276134 240618
rect 275514 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 276134 205174
rect 275514 204854 276134 204938
rect 275514 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 276134 204854
rect 275514 169174 276134 204618
rect 275514 168938 275546 169174
rect 275782 168938 275866 169174
rect 276102 168938 276134 169174
rect 275514 168854 276134 168938
rect 275514 168618 275546 168854
rect 275782 168618 275866 168854
rect 276102 168618 276134 168854
rect 275514 133174 276134 168618
rect 275514 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 276134 133174
rect 275514 132854 276134 132938
rect 275514 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 276134 132854
rect 275514 97174 276134 132618
rect 275514 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 276134 97174
rect 275514 96854 276134 96938
rect 275514 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 276134 96854
rect 275514 61174 276134 96618
rect 275514 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 276134 61174
rect 275514 60854 276134 60938
rect 275514 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 276134 60854
rect 275514 25174 276134 60618
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 604894 279854 640338
rect 279234 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 279854 604894
rect 279234 604574 279854 604658
rect 279234 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 279854 604574
rect 279234 568894 279854 604338
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 279234 532894 279854 568338
rect 279234 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 279854 532894
rect 279234 532574 279854 532658
rect 279234 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 279854 532574
rect 279234 496894 279854 532338
rect 279234 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 279854 496894
rect 279234 496574 279854 496658
rect 279234 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 279854 496574
rect 279234 460894 279854 496338
rect 279234 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 279854 460894
rect 279234 460574 279854 460658
rect 279234 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 279854 460574
rect 279234 424894 279854 460338
rect 279234 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 279854 424894
rect 279234 424574 279854 424658
rect 279234 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 279854 424574
rect 279234 388894 279854 424338
rect 279234 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 279854 388894
rect 279234 388574 279854 388658
rect 279234 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 279854 388574
rect 279234 352894 279854 388338
rect 279234 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 279854 352894
rect 279234 352574 279854 352658
rect 279234 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 279854 352574
rect 279234 316894 279854 352338
rect 279234 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 279854 316894
rect 279234 316574 279854 316658
rect 279234 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 279854 316574
rect 279234 280894 279854 316338
rect 279234 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 279854 280894
rect 279234 280574 279854 280658
rect 279234 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 279854 280574
rect 279234 244894 279854 280338
rect 279234 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 279854 244894
rect 279234 244574 279854 244658
rect 279234 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 279854 244574
rect 279234 208894 279854 244338
rect 279234 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 279854 208894
rect 279234 208574 279854 208658
rect 279234 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 279854 208574
rect 279234 172894 279854 208338
rect 279234 172658 279266 172894
rect 279502 172658 279586 172894
rect 279822 172658 279854 172894
rect 279234 172574 279854 172658
rect 279234 172338 279266 172574
rect 279502 172338 279586 172574
rect 279822 172338 279854 172574
rect 279234 136894 279854 172338
rect 279234 136658 279266 136894
rect 279502 136658 279586 136894
rect 279822 136658 279854 136894
rect 279234 136574 279854 136658
rect 279234 136338 279266 136574
rect 279502 136338 279586 136574
rect 279822 136338 279854 136574
rect 279234 100894 279854 136338
rect 279234 100658 279266 100894
rect 279502 100658 279586 100894
rect 279822 100658 279854 100894
rect 279234 100574 279854 100658
rect 279234 100338 279266 100574
rect 279502 100338 279586 100574
rect 279822 100338 279854 100574
rect 279234 64894 279854 100338
rect 279234 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 279854 64894
rect 279234 64574 279854 64658
rect 279234 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 279854 64574
rect 279234 28894 279854 64338
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 608614 283574 644058
rect 282954 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 283574 608614
rect 282954 608294 283574 608378
rect 282954 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 283574 608294
rect 282954 572614 283574 608058
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 536614 283574 572058
rect 282954 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 283574 536614
rect 282954 536294 283574 536378
rect 282954 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 283574 536294
rect 282954 500614 283574 536058
rect 282954 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 283574 500614
rect 282954 500294 283574 500378
rect 282954 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 283574 500294
rect 282954 464614 283574 500058
rect 282954 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 283574 464614
rect 282954 464294 283574 464378
rect 282954 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 283574 464294
rect 282954 428614 283574 464058
rect 282954 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 283574 428614
rect 282954 428294 283574 428378
rect 282954 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 283574 428294
rect 282954 392614 283574 428058
rect 282954 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 283574 392614
rect 282954 392294 283574 392378
rect 282954 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 283574 392294
rect 282954 356614 283574 392058
rect 282954 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 283574 356614
rect 282954 356294 283574 356378
rect 282954 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 283574 356294
rect 282954 320614 283574 356058
rect 282954 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 283574 320614
rect 282954 320294 283574 320378
rect 282954 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 283574 320294
rect 282954 284614 283574 320058
rect 282954 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 283574 284614
rect 282954 284294 283574 284378
rect 282954 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 283574 284294
rect 282954 248614 283574 284058
rect 282954 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 283574 248614
rect 282954 248294 283574 248378
rect 282954 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 283574 248294
rect 282954 212614 283574 248058
rect 282954 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 283574 212614
rect 282954 212294 283574 212378
rect 282954 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 283574 212294
rect 282954 176614 283574 212058
rect 282954 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 283574 176614
rect 282954 176294 283574 176378
rect 282954 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 283574 176294
rect 282954 140614 283574 176058
rect 282954 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 283574 140614
rect 282954 140294 283574 140378
rect 282954 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 283574 140294
rect 282954 104614 283574 140058
rect 282954 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 283574 104614
rect 282954 104294 283574 104378
rect 282954 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 283574 104294
rect 282954 68614 283574 104058
rect 282954 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 283574 68614
rect 282954 68294 283574 68378
rect 282954 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 283574 68294
rect 282954 32614 283574 68058
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 511174 294134 546618
rect 293514 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 294134 511174
rect 293514 510854 294134 510938
rect 293514 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 294134 510854
rect 293514 475174 294134 510618
rect 293514 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 294134 475174
rect 293514 474854 294134 474938
rect 293514 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 294134 474854
rect 293514 439174 294134 474618
rect 293514 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 294134 439174
rect 293514 438854 294134 438938
rect 293514 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 294134 438854
rect 293514 403174 294134 438618
rect 293514 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 294134 403174
rect 293514 402854 294134 402938
rect 293514 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 294134 402854
rect 293514 367174 294134 402618
rect 293514 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 294134 367174
rect 293514 366854 294134 366938
rect 293514 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 294134 366854
rect 293514 331174 294134 366618
rect 293514 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 294134 331174
rect 293514 330854 294134 330938
rect 293514 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 294134 330854
rect 293514 295174 294134 330618
rect 293514 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 294134 295174
rect 293514 294854 294134 294938
rect 293514 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 294134 294854
rect 293514 259174 294134 294618
rect 293514 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 294134 259174
rect 293514 258854 294134 258938
rect 293514 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 294134 258854
rect 293514 223174 294134 258618
rect 293514 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 294134 223174
rect 293514 222854 294134 222938
rect 293514 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 294134 222854
rect 293514 187174 294134 222618
rect 293514 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 294134 187174
rect 293514 186854 294134 186938
rect 293514 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 294134 186854
rect 293514 151174 294134 186618
rect 293514 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 294134 151174
rect 293514 150854 294134 150938
rect 293514 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 294134 150854
rect 293514 115174 294134 150618
rect 293514 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 294134 115174
rect 293514 114854 294134 114938
rect 293514 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 294134 114854
rect 293514 79174 294134 114618
rect 293514 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 294134 79174
rect 293514 78854 294134 78938
rect 293514 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 294134 78854
rect 293514 43174 294134 78618
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 514894 297854 550338
rect 297234 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 297854 514894
rect 297234 514574 297854 514658
rect 297234 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 297854 514574
rect 297234 478894 297854 514338
rect 297234 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 297854 478894
rect 297234 478574 297854 478658
rect 297234 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 297854 478574
rect 297234 442894 297854 478338
rect 297234 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 297854 442894
rect 297234 442574 297854 442658
rect 297234 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 297854 442574
rect 297234 406894 297854 442338
rect 297234 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 297854 406894
rect 297234 406574 297854 406658
rect 297234 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 297854 406574
rect 297234 370894 297854 406338
rect 297234 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 297854 370894
rect 297234 370574 297854 370658
rect 297234 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 297854 370574
rect 297234 334894 297854 370338
rect 297234 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 297854 334894
rect 297234 334574 297854 334658
rect 297234 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 297854 334574
rect 297234 298894 297854 334338
rect 297234 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 297854 298894
rect 297234 298574 297854 298658
rect 297234 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 297854 298574
rect 297234 262894 297854 298338
rect 297234 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 297854 262894
rect 297234 262574 297854 262658
rect 297234 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 297854 262574
rect 297234 226894 297854 262338
rect 297234 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 297854 226894
rect 297234 226574 297854 226658
rect 297234 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 297854 226574
rect 297234 190894 297854 226338
rect 297234 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 297854 190894
rect 297234 190574 297854 190658
rect 297234 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 297854 190574
rect 297234 154894 297854 190338
rect 297234 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 297854 154894
rect 297234 154574 297854 154658
rect 297234 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 297854 154574
rect 297234 118894 297854 154338
rect 297234 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 297854 118894
rect 297234 118574 297854 118658
rect 297234 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 297854 118574
rect 297234 82894 297854 118338
rect 297234 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 297854 82894
rect 297234 82574 297854 82658
rect 297234 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 297854 82574
rect 297234 46894 297854 82338
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 518614 301574 554058
rect 300954 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 301574 518614
rect 300954 518294 301574 518378
rect 300954 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 301574 518294
rect 300954 482614 301574 518058
rect 300954 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 301574 482614
rect 300954 482294 301574 482378
rect 300954 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 301574 482294
rect 300954 446614 301574 482058
rect 300954 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 301574 446614
rect 300954 446294 301574 446378
rect 300954 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 301574 446294
rect 300954 410614 301574 446058
rect 300954 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 301574 410614
rect 300954 410294 301574 410378
rect 300954 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 301574 410294
rect 300954 374614 301574 410058
rect 300954 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 301574 374614
rect 300954 374294 301574 374378
rect 300954 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 301574 374294
rect 300954 338614 301574 374058
rect 300954 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 301574 338614
rect 300954 338294 301574 338378
rect 300954 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 301574 338294
rect 300954 302614 301574 338058
rect 300954 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 301574 302614
rect 300954 302294 301574 302378
rect 300954 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 301574 302294
rect 300954 266614 301574 302058
rect 300954 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 301574 266614
rect 300954 266294 301574 266378
rect 300954 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 301574 266294
rect 300954 230614 301574 266058
rect 300954 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 301574 230614
rect 300954 230294 301574 230378
rect 300954 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 301574 230294
rect 300954 194614 301574 230058
rect 300954 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 301574 194614
rect 300954 194294 301574 194378
rect 300954 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 301574 194294
rect 300954 158614 301574 194058
rect 300954 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 301574 158614
rect 300954 158294 301574 158378
rect 300954 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 301574 158294
rect 300954 122614 301574 158058
rect 300954 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 301574 122614
rect 300954 122294 301574 122378
rect 300954 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 301574 122294
rect 300954 86614 301574 122058
rect 300954 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 301574 86614
rect 300954 86294 301574 86378
rect 300954 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 301574 86294
rect 300954 50614 301574 86058
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 529174 312134 564618
rect 311514 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 312134 529174
rect 311514 528854 312134 528938
rect 311514 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 312134 528854
rect 311514 493174 312134 528618
rect 311514 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 312134 493174
rect 311514 492854 312134 492938
rect 311514 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 312134 492854
rect 311514 457174 312134 492618
rect 311514 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 312134 457174
rect 311514 456854 312134 456938
rect 311514 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 312134 456854
rect 311514 421174 312134 456618
rect 311514 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 312134 421174
rect 311514 420854 312134 420938
rect 311514 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 312134 420854
rect 311514 385174 312134 420618
rect 311514 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 312134 385174
rect 311514 384854 312134 384938
rect 311514 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 312134 384854
rect 311514 349174 312134 384618
rect 311514 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 312134 349174
rect 311514 348854 312134 348938
rect 311514 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 312134 348854
rect 311514 313174 312134 348618
rect 311514 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 312134 313174
rect 311514 312854 312134 312938
rect 311514 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 312134 312854
rect 311514 277174 312134 312618
rect 311514 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 312134 277174
rect 311514 276854 312134 276938
rect 311514 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 312134 276854
rect 311514 241174 312134 276618
rect 311514 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 312134 241174
rect 311514 240854 312134 240938
rect 311514 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 312134 240854
rect 311514 205174 312134 240618
rect 311514 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 312134 205174
rect 311514 204854 312134 204938
rect 311514 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 312134 204854
rect 311514 169174 312134 204618
rect 311514 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 312134 169174
rect 311514 168854 312134 168938
rect 311514 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 312134 168854
rect 311514 133174 312134 168618
rect 311514 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 312134 133174
rect 311514 132854 312134 132938
rect 311514 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 312134 132854
rect 311514 97174 312134 132618
rect 311514 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 312134 97174
rect 311514 96854 312134 96938
rect 311514 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 312134 96854
rect 311514 61174 312134 96618
rect 311514 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 312134 61174
rect 311514 60854 312134 60938
rect 311514 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 312134 60854
rect 311514 25174 312134 60618
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 532894 315854 568338
rect 315234 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 315854 532894
rect 315234 532574 315854 532658
rect 315234 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 315854 532574
rect 315234 496894 315854 532338
rect 315234 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 315854 496894
rect 315234 496574 315854 496658
rect 315234 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 315854 496574
rect 315234 460894 315854 496338
rect 315234 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 315854 460894
rect 315234 460574 315854 460658
rect 315234 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 315854 460574
rect 315234 424894 315854 460338
rect 315234 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 315854 424894
rect 315234 424574 315854 424658
rect 315234 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 315854 424574
rect 315234 388894 315854 424338
rect 315234 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 315854 388894
rect 315234 388574 315854 388658
rect 315234 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 315854 388574
rect 315234 352894 315854 388338
rect 315234 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 315854 352894
rect 315234 352574 315854 352658
rect 315234 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 315854 352574
rect 315234 316894 315854 352338
rect 315234 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 315854 316894
rect 315234 316574 315854 316658
rect 315234 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 315854 316574
rect 315234 280894 315854 316338
rect 315234 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 315854 280894
rect 315234 280574 315854 280658
rect 315234 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 315854 280574
rect 315234 244894 315854 280338
rect 315234 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 315854 244894
rect 315234 244574 315854 244658
rect 315234 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 315854 244574
rect 315234 208894 315854 244338
rect 315234 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 315854 208894
rect 315234 208574 315854 208658
rect 315234 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 315854 208574
rect 315234 172894 315854 208338
rect 315234 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 315854 172894
rect 315234 172574 315854 172658
rect 315234 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 315854 172574
rect 315234 136894 315854 172338
rect 315234 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 315854 136894
rect 315234 136574 315854 136658
rect 315234 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 315854 136574
rect 315234 100894 315854 136338
rect 315234 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 315854 100894
rect 315234 100574 315854 100658
rect 315234 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 315854 100574
rect 315234 64894 315854 100338
rect 315234 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 315854 64894
rect 315234 64574 315854 64658
rect 315234 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 315854 64574
rect 315234 28894 315854 64338
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 536614 319574 572058
rect 318954 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 319574 536614
rect 318954 536294 319574 536378
rect 318954 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 319574 536294
rect 318954 500614 319574 536058
rect 318954 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 319574 500614
rect 318954 500294 319574 500378
rect 318954 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 319574 500294
rect 318954 464614 319574 500058
rect 318954 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 319574 464614
rect 318954 464294 319574 464378
rect 318954 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 319574 464294
rect 318954 428614 319574 464058
rect 318954 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 319574 428614
rect 318954 428294 319574 428378
rect 318954 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 319574 428294
rect 318954 392614 319574 428058
rect 318954 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 319574 392614
rect 318954 392294 319574 392378
rect 318954 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 319574 392294
rect 318954 356614 319574 392058
rect 318954 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 319574 356614
rect 318954 356294 319574 356378
rect 318954 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 319574 356294
rect 318954 320614 319574 356058
rect 318954 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 319574 320614
rect 318954 320294 319574 320378
rect 318954 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 319574 320294
rect 318954 284614 319574 320058
rect 318954 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 319574 284614
rect 318954 284294 319574 284378
rect 318954 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 319574 284294
rect 318954 248614 319574 284058
rect 318954 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 319574 248614
rect 318954 248294 319574 248378
rect 318954 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 319574 248294
rect 318954 212614 319574 248058
rect 318954 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 319574 212614
rect 318954 212294 319574 212378
rect 318954 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 319574 212294
rect 318954 176614 319574 212058
rect 318954 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 319574 176614
rect 318954 176294 319574 176378
rect 318954 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 319574 176294
rect 318954 140614 319574 176058
rect 318954 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 319574 140614
rect 318954 140294 319574 140378
rect 318954 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 319574 140294
rect 318954 104614 319574 140058
rect 318954 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 319574 104614
rect 318954 104294 319574 104378
rect 318954 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 319574 104294
rect 318954 68614 319574 104058
rect 318954 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 319574 68614
rect 318954 68294 319574 68378
rect 318954 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 319574 68294
rect 318954 32614 319574 68058
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547174 330134 582618
rect 329514 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 330134 547174
rect 329514 546854 330134 546938
rect 329514 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 330134 546854
rect 329514 511174 330134 546618
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 475174 330134 510618
rect 329514 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 330134 475174
rect 329514 474854 330134 474938
rect 329514 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 330134 474854
rect 329514 439174 330134 474618
rect 329514 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 330134 439174
rect 329514 438854 330134 438938
rect 329514 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 330134 438854
rect 329514 403174 330134 438618
rect 329514 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 330134 403174
rect 329514 402854 330134 402938
rect 329514 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 330134 402854
rect 329514 367174 330134 402618
rect 329514 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 330134 367174
rect 329514 366854 330134 366938
rect 329514 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 330134 366854
rect 329514 331174 330134 366618
rect 329514 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 330134 331174
rect 329514 330854 330134 330938
rect 329514 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 330134 330854
rect 329514 295174 330134 330618
rect 329514 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 330134 295174
rect 329514 294854 330134 294938
rect 329514 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 330134 294854
rect 329514 259174 330134 294618
rect 329514 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 330134 259174
rect 329514 258854 330134 258938
rect 329514 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 330134 258854
rect 329514 223174 330134 258618
rect 329514 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 330134 223174
rect 329514 222854 330134 222938
rect 329514 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 330134 222854
rect 329514 187174 330134 222618
rect 329514 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 330134 187174
rect 329514 186854 330134 186938
rect 329514 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 330134 186854
rect 329514 151174 330134 186618
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 115174 330134 150618
rect 329514 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 330134 115174
rect 329514 114854 330134 114938
rect 329514 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 330134 114854
rect 329514 79174 330134 114618
rect 329514 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 330134 79174
rect 329514 78854 330134 78938
rect 329514 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 330134 78854
rect 329514 43174 330134 78618
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 550894 333854 586338
rect 333234 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 333854 550894
rect 333234 550574 333854 550658
rect 333234 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 333854 550574
rect 333234 514894 333854 550338
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 478894 333854 514338
rect 333234 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 333854 478894
rect 333234 478574 333854 478658
rect 333234 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 333854 478574
rect 333234 442894 333854 478338
rect 333234 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 333854 442894
rect 333234 442574 333854 442658
rect 333234 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 333854 442574
rect 333234 406894 333854 442338
rect 333234 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 333854 406894
rect 333234 406574 333854 406658
rect 333234 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 333854 406574
rect 333234 370894 333854 406338
rect 333234 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 333854 370894
rect 333234 370574 333854 370658
rect 333234 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 333854 370574
rect 333234 334894 333854 370338
rect 333234 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 333854 334894
rect 333234 334574 333854 334658
rect 333234 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 333854 334574
rect 333234 298894 333854 334338
rect 333234 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 333854 298894
rect 333234 298574 333854 298658
rect 333234 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 333854 298574
rect 333234 262894 333854 298338
rect 333234 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 333854 262894
rect 333234 262574 333854 262658
rect 333234 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 333854 262574
rect 333234 226894 333854 262338
rect 333234 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 333854 226894
rect 333234 226574 333854 226658
rect 333234 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 333854 226574
rect 333234 190894 333854 226338
rect 333234 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 333854 190894
rect 333234 190574 333854 190658
rect 333234 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 333854 190574
rect 333234 154894 333854 190338
rect 333234 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 333854 154894
rect 333234 154574 333854 154658
rect 333234 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 333854 154574
rect 333234 118894 333854 154338
rect 333234 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 333854 118894
rect 333234 118574 333854 118658
rect 333234 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 333854 118574
rect 333234 82894 333854 118338
rect 333234 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 333854 82894
rect 333234 82574 333854 82658
rect 333234 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 333854 82574
rect 333234 46894 333854 82338
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 336954 518614 337574 554058
rect 336954 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 337574 518614
rect 336954 518294 337574 518378
rect 336954 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 337574 518294
rect 336954 482614 337574 518058
rect 336954 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 337574 482614
rect 336954 482294 337574 482378
rect 336954 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 337574 482294
rect 336954 446614 337574 482058
rect 336954 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 337574 446614
rect 336954 446294 337574 446378
rect 336954 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 337574 446294
rect 336954 410614 337574 446058
rect 336954 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 337574 410614
rect 336954 410294 337574 410378
rect 336954 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 337574 410294
rect 336954 374614 337574 410058
rect 336954 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 337574 374614
rect 336954 374294 337574 374378
rect 336954 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 337574 374294
rect 336954 338614 337574 374058
rect 336954 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 337574 338614
rect 336954 338294 337574 338378
rect 336954 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 337574 338294
rect 336954 302614 337574 338058
rect 336954 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 337574 302614
rect 336954 302294 337574 302378
rect 336954 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 337574 302294
rect 336954 266614 337574 302058
rect 336954 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 337574 266614
rect 336954 266294 337574 266378
rect 336954 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 337574 266294
rect 336954 230614 337574 266058
rect 336954 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 337574 230614
rect 336954 230294 337574 230378
rect 336954 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 337574 230294
rect 336954 194614 337574 230058
rect 336954 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 337574 194614
rect 336954 194294 337574 194378
rect 336954 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 337574 194294
rect 336954 158614 337574 194058
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 336954 122614 337574 158058
rect 336954 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 337574 122614
rect 336954 122294 337574 122378
rect 336954 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 337574 122294
rect 336954 86614 337574 122058
rect 336954 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 337574 86614
rect 336954 86294 337574 86378
rect 336954 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 337574 86294
rect 336954 50614 337574 86058
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 565174 348134 600618
rect 347514 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 348134 565174
rect 347514 564854 348134 564938
rect 347514 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 348134 564854
rect 347514 529174 348134 564618
rect 347514 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 348134 529174
rect 347514 528854 348134 528938
rect 347514 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 348134 528854
rect 347514 493174 348134 528618
rect 347514 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 348134 493174
rect 347514 492854 348134 492938
rect 347514 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 348134 492854
rect 347514 457174 348134 492618
rect 347514 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 348134 457174
rect 347514 456854 348134 456938
rect 347514 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 348134 456854
rect 347514 421174 348134 456618
rect 347514 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 348134 421174
rect 347514 420854 348134 420938
rect 347514 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 348134 420854
rect 347514 385174 348134 420618
rect 347514 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 348134 385174
rect 347514 384854 348134 384938
rect 347514 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 348134 384854
rect 347514 349174 348134 384618
rect 347514 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 348134 349174
rect 347514 348854 348134 348938
rect 347514 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 348134 348854
rect 347514 313174 348134 348618
rect 347514 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 348134 313174
rect 347514 312854 348134 312938
rect 347514 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 348134 312854
rect 347514 277174 348134 312618
rect 347514 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 348134 277174
rect 347514 276854 348134 276938
rect 347514 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 348134 276854
rect 347514 241174 348134 276618
rect 347514 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 348134 241174
rect 347514 240854 348134 240938
rect 347514 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 348134 240854
rect 347514 205174 348134 240618
rect 347514 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 348134 205174
rect 347514 204854 348134 204938
rect 347514 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 348134 204854
rect 347514 169174 348134 204618
rect 347514 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 348134 169174
rect 347514 168854 348134 168938
rect 347514 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 348134 168854
rect 347514 133174 348134 168618
rect 347514 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 348134 133174
rect 347514 132854 348134 132938
rect 347514 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 348134 132854
rect 347514 97174 348134 132618
rect 347514 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 348134 97174
rect 347514 96854 348134 96938
rect 347514 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 348134 96854
rect 347514 61174 348134 96618
rect 347514 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 348134 61174
rect 347514 60854 348134 60938
rect 347514 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 348134 60854
rect 347514 25174 348134 60618
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 568894 351854 604338
rect 351234 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 351854 568894
rect 351234 568574 351854 568658
rect 351234 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 351854 568574
rect 351234 532894 351854 568338
rect 351234 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 351854 532894
rect 351234 532574 351854 532658
rect 351234 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 351854 532574
rect 351234 496894 351854 532338
rect 351234 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 351854 496894
rect 351234 496574 351854 496658
rect 351234 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 351854 496574
rect 351234 460894 351854 496338
rect 351234 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 351854 460894
rect 351234 460574 351854 460658
rect 351234 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 351854 460574
rect 351234 424894 351854 460338
rect 351234 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 351854 424894
rect 351234 424574 351854 424658
rect 351234 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 351854 424574
rect 351234 388894 351854 424338
rect 351234 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 351854 388894
rect 351234 388574 351854 388658
rect 351234 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 351854 388574
rect 351234 352894 351854 388338
rect 351234 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 351854 352894
rect 351234 352574 351854 352658
rect 351234 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 351854 352574
rect 351234 316894 351854 352338
rect 351234 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 351854 316894
rect 351234 316574 351854 316658
rect 351234 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 351854 316574
rect 351234 280894 351854 316338
rect 351234 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 351854 280894
rect 351234 280574 351854 280658
rect 351234 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 351854 280574
rect 351234 244894 351854 280338
rect 351234 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 351854 244894
rect 351234 244574 351854 244658
rect 351234 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 351854 244574
rect 351234 208894 351854 244338
rect 351234 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 351854 208894
rect 351234 208574 351854 208658
rect 351234 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 351854 208574
rect 351234 172894 351854 208338
rect 351234 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 351854 172894
rect 351234 172574 351854 172658
rect 351234 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 351854 172574
rect 351234 136894 351854 172338
rect 351234 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 351854 136894
rect 351234 136574 351854 136658
rect 351234 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 351854 136574
rect 351234 100894 351854 136338
rect 351234 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 351854 100894
rect 351234 100574 351854 100658
rect 351234 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 351854 100574
rect 351234 64894 351854 100338
rect 351234 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 351854 64894
rect 351234 64574 351854 64658
rect 351234 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 351854 64574
rect 351234 28894 351854 64338
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 354954 536614 355574 572058
rect 354954 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 355574 536614
rect 354954 536294 355574 536378
rect 354954 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 355574 536294
rect 354954 500614 355574 536058
rect 354954 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 355574 500614
rect 354954 500294 355574 500378
rect 354954 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 355574 500294
rect 354954 464614 355574 500058
rect 354954 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 355574 464614
rect 354954 464294 355574 464378
rect 354954 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 355574 464294
rect 354954 428614 355574 464058
rect 354954 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 355574 428614
rect 354954 428294 355574 428378
rect 354954 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 355574 428294
rect 354954 392614 355574 428058
rect 354954 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 355574 392614
rect 354954 392294 355574 392378
rect 354954 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 355574 392294
rect 354954 356614 355574 392058
rect 354954 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 355574 356614
rect 354954 356294 355574 356378
rect 354954 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 355574 356294
rect 354954 320614 355574 356058
rect 354954 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 355574 320614
rect 354954 320294 355574 320378
rect 354954 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 355574 320294
rect 354954 284614 355574 320058
rect 354954 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 355574 284614
rect 354954 284294 355574 284378
rect 354954 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 355574 284294
rect 354954 248614 355574 284058
rect 354954 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 355574 248614
rect 354954 248294 355574 248378
rect 354954 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 355574 248294
rect 354954 212614 355574 248058
rect 354954 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 355574 212614
rect 354954 212294 355574 212378
rect 354954 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 355574 212294
rect 354954 176614 355574 212058
rect 354954 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 355574 176614
rect 354954 176294 355574 176378
rect 354954 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 355574 176294
rect 354954 140614 355574 176058
rect 354954 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 355574 140614
rect 354954 140294 355574 140378
rect 354954 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 355574 140294
rect 354954 104614 355574 140058
rect 354954 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 355574 104614
rect 354954 104294 355574 104378
rect 354954 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 355574 104294
rect 354954 68614 355574 104058
rect 354954 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 355574 68614
rect 354954 68294 355574 68378
rect 354954 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 355574 68294
rect 354954 32614 355574 68058
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 365514 367174 366134 402618
rect 365514 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 366134 367174
rect 365514 366854 366134 366938
rect 365514 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 366134 366854
rect 365514 331174 366134 366618
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 295174 366134 330618
rect 365514 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 366134 295174
rect 365514 294854 366134 294938
rect 365514 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 366134 294854
rect 365514 259174 366134 294618
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 223174 366134 258618
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 370894 369854 406338
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 369234 334894 369854 370338
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 369234 298894 369854 334338
rect 369234 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 369854 298894
rect 369234 298574 369854 298658
rect 369234 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 369854 298574
rect 369234 262894 369854 298338
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 226894 369854 262338
rect 369234 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 369854 226894
rect 369234 226574 369854 226658
rect 369234 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 369854 226574
rect 369234 190894 369854 226338
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 154894 369854 190338
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 338614 373574 374058
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 230614 373574 266058
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 565174 384134 600618
rect 383514 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 384134 565174
rect 383514 564854 384134 564938
rect 383514 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 384134 564854
rect 383514 529174 384134 564618
rect 383514 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 384134 529174
rect 383514 528854 384134 528938
rect 383514 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 384134 528854
rect 383514 493174 384134 528618
rect 383514 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 384134 493174
rect 383514 492854 384134 492938
rect 383514 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 384134 492854
rect 383514 457174 384134 492618
rect 383514 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 384134 457174
rect 383514 456854 384134 456938
rect 383514 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 384134 456854
rect 383514 421174 384134 456618
rect 383514 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 384134 421174
rect 383514 420854 384134 420938
rect 383514 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 384134 420854
rect 383514 385174 384134 420618
rect 383514 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 384134 385174
rect 383514 384854 384134 384938
rect 383514 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 384134 384854
rect 383514 349174 384134 384618
rect 383514 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 384134 349174
rect 383514 348854 384134 348938
rect 383514 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 384134 348854
rect 383514 313174 384134 348618
rect 383514 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 384134 313174
rect 383514 312854 384134 312938
rect 383514 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 384134 312854
rect 383514 277174 384134 312618
rect 383514 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 384134 277174
rect 383514 276854 384134 276938
rect 383514 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 384134 276854
rect 383514 241174 384134 276618
rect 383514 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 384134 241174
rect 383514 240854 384134 240938
rect 383514 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 384134 240854
rect 383514 205174 384134 240618
rect 383514 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 384134 205174
rect 383514 204854 384134 204938
rect 383514 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 384134 204854
rect 383514 169174 384134 204618
rect 383514 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 384134 169174
rect 383514 168854 384134 168938
rect 383514 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 384134 168854
rect 383514 133174 384134 168618
rect 383514 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 384134 133174
rect 383514 132854 384134 132938
rect 383514 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 384134 132854
rect 383514 97174 384134 132618
rect 383514 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 384134 97174
rect 383514 96854 384134 96938
rect 383514 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 384134 96854
rect 383514 61174 384134 96618
rect 383514 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 384134 61174
rect 383514 60854 384134 60938
rect 383514 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 384134 60854
rect 383514 25174 384134 60618
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 568894 387854 604338
rect 387234 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 387854 568894
rect 387234 568574 387854 568658
rect 387234 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 387854 568574
rect 387234 532894 387854 568338
rect 387234 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 387854 532894
rect 387234 532574 387854 532658
rect 387234 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 387854 532574
rect 387234 496894 387854 532338
rect 387234 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 387854 496894
rect 387234 496574 387854 496658
rect 387234 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 387854 496574
rect 387234 460894 387854 496338
rect 387234 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 387854 460894
rect 387234 460574 387854 460658
rect 387234 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 387854 460574
rect 387234 424894 387854 460338
rect 387234 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 387854 424894
rect 387234 424574 387854 424658
rect 387234 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 387854 424574
rect 387234 388894 387854 424338
rect 387234 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 387854 388894
rect 387234 388574 387854 388658
rect 387234 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 387854 388574
rect 387234 352894 387854 388338
rect 387234 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 387854 352894
rect 387234 352574 387854 352658
rect 387234 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 387854 352574
rect 387234 316894 387854 352338
rect 387234 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 387854 316894
rect 387234 316574 387854 316658
rect 387234 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 387854 316574
rect 387234 280894 387854 316338
rect 387234 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 387854 280894
rect 387234 280574 387854 280658
rect 387234 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 387854 280574
rect 387234 244894 387854 280338
rect 387234 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 387854 244894
rect 387234 244574 387854 244658
rect 387234 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 387854 244574
rect 387234 208894 387854 244338
rect 387234 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 387854 208894
rect 387234 208574 387854 208658
rect 387234 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 387854 208574
rect 387234 172894 387854 208338
rect 387234 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 387854 172894
rect 387234 172574 387854 172658
rect 387234 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 387854 172574
rect 387234 136894 387854 172338
rect 387234 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 387854 136894
rect 387234 136574 387854 136658
rect 387234 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 387854 136574
rect 387234 100894 387854 136338
rect 387234 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 387854 100894
rect 387234 100574 387854 100658
rect 387234 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 387854 100574
rect 387234 64894 387854 100338
rect 387234 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 387854 64894
rect 387234 64574 387854 64658
rect 387234 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 387854 64574
rect 387234 28894 387854 64338
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 390954 536614 391574 572058
rect 390954 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 391574 536614
rect 390954 536294 391574 536378
rect 390954 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 391574 536294
rect 390954 500614 391574 536058
rect 390954 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 391574 500614
rect 390954 500294 391574 500378
rect 390954 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 391574 500294
rect 390954 464614 391574 500058
rect 390954 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 391574 464614
rect 390954 464294 391574 464378
rect 390954 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 391574 464294
rect 390954 428614 391574 464058
rect 390954 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 391574 428614
rect 390954 428294 391574 428378
rect 390954 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 391574 428294
rect 390954 392614 391574 428058
rect 390954 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 391574 392614
rect 390954 392294 391574 392378
rect 390954 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 391574 392294
rect 390954 356614 391574 392058
rect 390954 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 391574 356614
rect 390954 356294 391574 356378
rect 390954 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 391574 356294
rect 390954 320614 391574 356058
rect 390954 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 391574 320614
rect 390954 320294 391574 320378
rect 390954 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 391574 320294
rect 390954 284614 391574 320058
rect 390954 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 391574 284614
rect 390954 284294 391574 284378
rect 390954 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 391574 284294
rect 390954 248614 391574 284058
rect 390954 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 391574 248614
rect 390954 248294 391574 248378
rect 390954 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 391574 248294
rect 390954 212614 391574 248058
rect 390954 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 391574 212614
rect 390954 212294 391574 212378
rect 390954 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 391574 212294
rect 390954 176614 391574 212058
rect 390954 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 391574 176614
rect 390954 176294 391574 176378
rect 390954 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 391574 176294
rect 390954 140614 391574 176058
rect 390954 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 391574 140614
rect 390954 140294 391574 140378
rect 390954 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 391574 140294
rect 390954 104614 391574 140058
rect 390954 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 391574 104614
rect 390954 104294 391574 104378
rect 390954 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 391574 104294
rect 390954 68614 391574 104058
rect 390954 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 391574 68614
rect 390954 68294 391574 68378
rect 390954 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 391574 68294
rect 390954 32614 391574 68058
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 439174 402134 474618
rect 401514 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 402134 439174
rect 401514 438854 402134 438938
rect 401514 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 402134 438854
rect 401514 403174 402134 438618
rect 401514 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 402134 403174
rect 401514 402854 402134 402938
rect 401514 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 402134 402854
rect 401514 367174 402134 402618
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 331174 402134 366618
rect 401514 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 402134 331174
rect 401514 330854 402134 330938
rect 401514 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 402134 330854
rect 401514 295174 402134 330618
rect 401514 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 402134 295174
rect 401514 294854 402134 294938
rect 401514 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 402134 294854
rect 401514 259174 402134 294618
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 223174 402134 258618
rect 401514 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 402134 223174
rect 401514 222854 402134 222938
rect 401514 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 402134 222854
rect 401514 187174 402134 222618
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 151174 402134 186618
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 79174 402134 114618
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 442894 405854 478338
rect 405234 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 405854 442894
rect 405234 442574 405854 442658
rect 405234 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 405854 442574
rect 405234 406894 405854 442338
rect 405234 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 405854 406894
rect 405234 406574 405854 406658
rect 405234 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 405854 406574
rect 405234 370894 405854 406338
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 334894 405854 370338
rect 405234 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 405854 334894
rect 405234 334574 405854 334658
rect 405234 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 405854 334574
rect 405234 298894 405854 334338
rect 405234 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 405854 298894
rect 405234 298574 405854 298658
rect 405234 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 405854 298574
rect 405234 262894 405854 298338
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 226894 405854 262338
rect 405234 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 405854 226894
rect 405234 226574 405854 226658
rect 405234 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 405854 226574
rect 405234 190894 405854 226338
rect 405234 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 405854 190894
rect 405234 190574 405854 190658
rect 405234 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 405854 190574
rect 405234 154894 405854 190338
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 118894 405854 154338
rect 405234 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 405854 118894
rect 405234 118574 405854 118658
rect 405234 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 405854 118574
rect 405234 82894 405854 118338
rect 405234 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 405854 82894
rect 405234 82574 405854 82658
rect 405234 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 405854 82574
rect 405234 46894 405854 82338
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 446614 409574 482058
rect 408954 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 409574 446614
rect 408954 446294 409574 446378
rect 408954 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 409574 446294
rect 408954 410614 409574 446058
rect 408954 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 409574 410614
rect 408954 410294 409574 410378
rect 408954 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 409574 410294
rect 408954 374614 409574 410058
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 408954 338614 409574 374058
rect 408954 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 409574 338614
rect 408954 338294 409574 338378
rect 408954 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 409574 338294
rect 408954 302614 409574 338058
rect 408954 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 409574 302614
rect 408954 302294 409574 302378
rect 408954 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 409574 302294
rect 408954 266614 409574 302058
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 230614 409574 266058
rect 408954 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 409574 230614
rect 408954 230294 409574 230378
rect 408954 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 409574 230294
rect 408954 194614 409574 230058
rect 408954 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 409574 194614
rect 408954 194294 409574 194378
rect 408954 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 409574 194294
rect 408954 158614 409574 194058
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 122614 409574 158058
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 408954 86614 409574 122058
rect 408954 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 409574 86614
rect 408954 86294 409574 86378
rect 408954 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 409574 86294
rect 408954 50614 409574 86058
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 565174 420134 600618
rect 419514 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 420134 565174
rect 419514 564854 420134 564938
rect 419514 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 420134 564854
rect 419514 529174 420134 564618
rect 419514 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 420134 529174
rect 419514 528854 420134 528938
rect 419514 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 420134 528854
rect 419514 493174 420134 528618
rect 419514 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 420134 493174
rect 419514 492854 420134 492938
rect 419514 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 420134 492854
rect 419514 457174 420134 492618
rect 419514 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 420134 457174
rect 419514 456854 420134 456938
rect 419514 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 420134 456854
rect 419514 421174 420134 456618
rect 419514 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 420134 421174
rect 419514 420854 420134 420938
rect 419514 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 420134 420854
rect 419514 385174 420134 420618
rect 419514 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 420134 385174
rect 419514 384854 420134 384938
rect 419514 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 420134 384854
rect 419514 349174 420134 384618
rect 419514 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 420134 349174
rect 419514 348854 420134 348938
rect 419514 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 420134 348854
rect 419514 313174 420134 348618
rect 419514 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 420134 313174
rect 419514 312854 420134 312938
rect 419514 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 420134 312854
rect 419514 277174 420134 312618
rect 419514 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 420134 277174
rect 419514 276854 420134 276938
rect 419514 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 420134 276854
rect 419514 241174 420134 276618
rect 419514 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 420134 241174
rect 419514 240854 420134 240938
rect 419514 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 420134 240854
rect 419514 205174 420134 240618
rect 419514 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 420134 205174
rect 419514 204854 420134 204938
rect 419514 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 420134 204854
rect 419514 169174 420134 204618
rect 419514 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 420134 169174
rect 419514 168854 420134 168938
rect 419514 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 420134 168854
rect 419514 133174 420134 168618
rect 419514 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 420134 133174
rect 419514 132854 420134 132938
rect 419514 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 420134 132854
rect 419514 97174 420134 132618
rect 419514 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 420134 97174
rect 419514 96854 420134 96938
rect 419514 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 420134 96854
rect 419514 61174 420134 96618
rect 419514 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 420134 61174
rect 419514 60854 420134 60938
rect 419514 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 420134 60854
rect 419514 25174 420134 60618
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 568894 423854 604338
rect 423234 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 423854 568894
rect 423234 568574 423854 568658
rect 423234 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 423854 568574
rect 423234 532894 423854 568338
rect 423234 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 423854 532894
rect 423234 532574 423854 532658
rect 423234 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 423854 532574
rect 423234 496894 423854 532338
rect 423234 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 423854 496894
rect 423234 496574 423854 496658
rect 423234 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 423854 496574
rect 423234 460894 423854 496338
rect 423234 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 423854 460894
rect 423234 460574 423854 460658
rect 423234 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 423854 460574
rect 423234 424894 423854 460338
rect 423234 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 423854 424894
rect 423234 424574 423854 424658
rect 423234 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 423854 424574
rect 423234 388894 423854 424338
rect 423234 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 423854 388894
rect 423234 388574 423854 388658
rect 423234 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 423854 388574
rect 423234 352894 423854 388338
rect 423234 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 423854 352894
rect 423234 352574 423854 352658
rect 423234 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 423854 352574
rect 423234 316894 423854 352338
rect 423234 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 423854 316894
rect 423234 316574 423854 316658
rect 423234 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 423854 316574
rect 423234 280894 423854 316338
rect 423234 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 423854 280894
rect 423234 280574 423854 280658
rect 423234 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 423854 280574
rect 423234 244894 423854 280338
rect 423234 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 423854 244894
rect 423234 244574 423854 244658
rect 423234 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 423854 244574
rect 423234 208894 423854 244338
rect 423234 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 423854 208894
rect 423234 208574 423854 208658
rect 423234 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 423854 208574
rect 423234 172894 423854 208338
rect 423234 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 423854 172894
rect 423234 172574 423854 172658
rect 423234 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 423854 172574
rect 423234 136894 423854 172338
rect 423234 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 423854 136894
rect 423234 136574 423854 136658
rect 423234 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 423854 136574
rect 423234 100894 423854 136338
rect 423234 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 423854 100894
rect 423234 100574 423854 100658
rect 423234 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 423854 100574
rect 423234 64894 423854 100338
rect 423234 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 423854 64894
rect 423234 64574 423854 64658
rect 423234 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 423854 64574
rect 423234 28894 423854 64338
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 572614 427574 608058
rect 426954 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 427574 572614
rect 426954 572294 427574 572378
rect 426954 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 427574 572294
rect 426954 536614 427574 572058
rect 426954 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 427574 536614
rect 426954 536294 427574 536378
rect 426954 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 427574 536294
rect 426954 500614 427574 536058
rect 426954 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 427574 500614
rect 426954 500294 427574 500378
rect 426954 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 427574 500294
rect 426954 464614 427574 500058
rect 426954 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 427574 464614
rect 426954 464294 427574 464378
rect 426954 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 427574 464294
rect 426954 428614 427574 464058
rect 426954 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 427574 428614
rect 426954 428294 427574 428378
rect 426954 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 427574 428294
rect 426954 392614 427574 428058
rect 426954 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 427574 392614
rect 426954 392294 427574 392378
rect 426954 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 427574 392294
rect 426954 356614 427574 392058
rect 426954 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 427574 356614
rect 426954 356294 427574 356378
rect 426954 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 427574 356294
rect 426954 320614 427574 356058
rect 426954 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 427574 320614
rect 426954 320294 427574 320378
rect 426954 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 427574 320294
rect 426954 284614 427574 320058
rect 426954 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 427574 284614
rect 426954 284294 427574 284378
rect 426954 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 427574 284294
rect 426954 248614 427574 284058
rect 426954 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 427574 248614
rect 426954 248294 427574 248378
rect 426954 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 427574 248294
rect 426954 212614 427574 248058
rect 426954 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 427574 212614
rect 426954 212294 427574 212378
rect 426954 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 427574 212294
rect 426954 176614 427574 212058
rect 426954 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 427574 176614
rect 426954 176294 427574 176378
rect 426954 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 427574 176294
rect 426954 140614 427574 176058
rect 426954 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 427574 140614
rect 426954 140294 427574 140378
rect 426954 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 427574 140294
rect 426954 104614 427574 140058
rect 426954 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 427574 104614
rect 426954 104294 427574 104378
rect 426954 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 427574 104294
rect 426954 68614 427574 104058
rect 426954 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 427574 68614
rect 426954 68294 427574 68378
rect 426954 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 427574 68294
rect 426954 32614 427574 68058
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 439174 438134 474618
rect 437514 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 438134 439174
rect 437514 438854 438134 438938
rect 437514 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 438134 438854
rect 437514 403174 438134 438618
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 437514 367174 438134 402618
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 331174 438134 366618
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 295174 438134 330618
rect 437514 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 438134 295174
rect 437514 294854 438134 294938
rect 437514 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 438134 294854
rect 437514 259174 438134 294618
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 223174 438134 258618
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 187174 438134 222618
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 151174 438134 186618
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 437514 115174 438134 150618
rect 437514 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 438134 115174
rect 437514 114854 438134 114938
rect 437514 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 438134 114854
rect 437514 79174 438134 114618
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 442894 441854 478338
rect 441234 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 441854 442894
rect 441234 442574 441854 442658
rect 441234 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 441854 442574
rect 441234 406894 441854 442338
rect 441234 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 441854 406894
rect 441234 406574 441854 406658
rect 441234 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 441854 406574
rect 441234 370894 441854 406338
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 334894 441854 370338
rect 441234 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 441854 334894
rect 441234 334574 441854 334658
rect 441234 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 441854 334574
rect 441234 298894 441854 334338
rect 441234 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 441854 298894
rect 441234 298574 441854 298658
rect 441234 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 441854 298574
rect 441234 262894 441854 298338
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 226894 441854 262338
rect 441234 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 441854 226894
rect 441234 226574 441854 226658
rect 441234 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 441854 226574
rect 441234 190894 441854 226338
rect 441234 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 441854 190894
rect 441234 190574 441854 190658
rect 441234 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 441854 190574
rect 441234 154894 441854 190338
rect 441234 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 441854 154894
rect 441234 154574 441854 154658
rect 441234 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 441854 154574
rect 441234 118894 441854 154338
rect 441234 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 441854 118894
rect 441234 118574 441854 118658
rect 441234 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 441854 118574
rect 441234 82894 441854 118338
rect 441234 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 441854 82894
rect 441234 82574 441854 82658
rect 441234 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 441854 82574
rect 441234 46894 441854 82338
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 444954 410614 445574 446058
rect 444954 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 445574 410614
rect 444954 410294 445574 410378
rect 444954 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 445574 410294
rect 444954 374614 445574 410058
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 444954 338614 445574 374058
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 444954 302614 445574 338058
rect 444954 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 445574 302614
rect 444954 302294 445574 302378
rect 444954 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 445574 302294
rect 444954 266614 445574 302058
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 230614 445574 266058
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 444954 158614 445574 194058
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 444954 122614 445574 158058
rect 444954 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 445574 122614
rect 444954 122294 445574 122378
rect 444954 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 445574 122294
rect 444954 86614 445574 122058
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 444954 50614 445574 86058
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 529174 456134 564618
rect 455514 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 456134 529174
rect 455514 528854 456134 528938
rect 455514 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 456134 528854
rect 455514 493174 456134 528618
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 455514 457174 456134 492618
rect 455514 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 456134 457174
rect 455514 456854 456134 456938
rect 455514 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 456134 456854
rect 455514 421174 456134 456618
rect 455514 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 456134 421174
rect 455514 420854 456134 420938
rect 455514 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 456134 420854
rect 455514 385174 456134 420618
rect 455514 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 456134 385174
rect 455514 384854 456134 384938
rect 455514 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 456134 384854
rect 455514 349174 456134 384618
rect 455514 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 456134 349174
rect 455514 348854 456134 348938
rect 455514 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 456134 348854
rect 455514 313174 456134 348618
rect 455514 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 456134 313174
rect 455514 312854 456134 312938
rect 455514 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 456134 312854
rect 455514 277174 456134 312618
rect 455514 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 456134 277174
rect 455514 276854 456134 276938
rect 455514 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 456134 276854
rect 455514 241174 456134 276618
rect 455514 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 456134 241174
rect 455514 240854 456134 240938
rect 455514 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 456134 240854
rect 455514 205174 456134 240618
rect 455514 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 456134 205174
rect 455514 204854 456134 204938
rect 455514 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 456134 204854
rect 455514 169174 456134 204618
rect 455514 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 456134 169174
rect 455514 168854 456134 168938
rect 455514 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 456134 168854
rect 455514 133174 456134 168618
rect 455514 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 456134 133174
rect 455514 132854 456134 132938
rect 455514 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 456134 132854
rect 455514 97174 456134 132618
rect 455514 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 456134 97174
rect 455514 96854 456134 96938
rect 455514 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 456134 96854
rect 455514 61174 456134 96618
rect 455514 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 456134 61174
rect 455514 60854 456134 60938
rect 455514 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 456134 60854
rect 455514 25174 456134 60618
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 568894 459854 604338
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 532894 459854 568338
rect 459234 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 459854 532894
rect 459234 532574 459854 532658
rect 459234 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 459854 532574
rect 459234 496894 459854 532338
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 460894 459854 496338
rect 459234 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 459854 460894
rect 459234 460574 459854 460658
rect 459234 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 459854 460574
rect 459234 424894 459854 460338
rect 459234 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 459854 424894
rect 459234 424574 459854 424658
rect 459234 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 459854 424574
rect 459234 388894 459854 424338
rect 459234 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 459854 388894
rect 459234 388574 459854 388658
rect 459234 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 459854 388574
rect 459234 352894 459854 388338
rect 459234 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 459854 352894
rect 459234 352574 459854 352658
rect 459234 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 459854 352574
rect 459234 316894 459854 352338
rect 459234 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 459854 316894
rect 459234 316574 459854 316658
rect 459234 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 459854 316574
rect 459234 280894 459854 316338
rect 459234 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 459854 280894
rect 459234 280574 459854 280658
rect 459234 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 459854 280574
rect 459234 244894 459854 280338
rect 459234 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 459854 244894
rect 459234 244574 459854 244658
rect 459234 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 459854 244574
rect 459234 208894 459854 244338
rect 459234 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 459854 208894
rect 459234 208574 459854 208658
rect 459234 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 459854 208574
rect 459234 172894 459854 208338
rect 459234 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 459854 172894
rect 459234 172574 459854 172658
rect 459234 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 459854 172574
rect 459234 136894 459854 172338
rect 459234 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 459854 136894
rect 459234 136574 459854 136658
rect 459234 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 459854 136574
rect 459234 100894 459854 136338
rect 459234 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 459854 100894
rect 459234 100574 459854 100658
rect 459234 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 459854 100574
rect 459234 64894 459854 100338
rect 459234 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 459854 64894
rect 459234 64574 459854 64658
rect 459234 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 459854 64574
rect 459234 28894 459854 64338
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 572614 463574 608058
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 536614 463574 572058
rect 462954 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 463574 536614
rect 462954 536294 463574 536378
rect 462954 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 463574 536294
rect 462954 500614 463574 536058
rect 462954 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 463574 500614
rect 462954 500294 463574 500378
rect 462954 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 463574 500294
rect 462954 464614 463574 500058
rect 462954 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 463574 464614
rect 462954 464294 463574 464378
rect 462954 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 463574 464294
rect 462954 428614 463574 464058
rect 462954 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 463574 428614
rect 462954 428294 463574 428378
rect 462954 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 463574 428294
rect 462954 392614 463574 428058
rect 462954 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 463574 392614
rect 462954 392294 463574 392378
rect 462954 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 463574 392294
rect 462954 356614 463574 392058
rect 462954 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 463574 356614
rect 462954 356294 463574 356378
rect 462954 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 463574 356294
rect 462954 320614 463574 356058
rect 462954 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 463574 320614
rect 462954 320294 463574 320378
rect 462954 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 463574 320294
rect 462954 284614 463574 320058
rect 462954 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 463574 284614
rect 462954 284294 463574 284378
rect 462954 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 463574 284294
rect 462954 248614 463574 284058
rect 462954 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 463574 248614
rect 462954 248294 463574 248378
rect 462954 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 463574 248294
rect 462954 212614 463574 248058
rect 462954 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 463574 212614
rect 462954 212294 463574 212378
rect 462954 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 463574 212294
rect 462954 176614 463574 212058
rect 462954 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 463574 176614
rect 462954 176294 463574 176378
rect 462954 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 463574 176294
rect 462954 140614 463574 176058
rect 462954 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 463574 140614
rect 462954 140294 463574 140378
rect 462954 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 463574 140294
rect 462954 104614 463574 140058
rect 462954 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 463574 104614
rect 462954 104294 463574 104378
rect 462954 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 463574 104294
rect 462954 68614 463574 104058
rect 462954 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 463574 68614
rect 462954 68294 463574 68378
rect 462954 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 463574 68294
rect 462954 32614 463574 68058
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 439174 474134 474618
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 473514 403174 474134 438618
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 473514 367174 474134 402618
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 331174 474134 366618
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 473514 295174 474134 330618
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 473514 259174 474134 294618
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 223174 474134 258618
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 406894 477854 442338
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 477234 370894 477854 406338
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 334894 477854 370338
rect 477234 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 477854 334894
rect 477234 334574 477854 334658
rect 477234 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 477854 334574
rect 477234 298894 477854 334338
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 226894 477854 262338
rect 477234 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 477854 226894
rect 477234 226574 477854 226658
rect 477234 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 477854 226574
rect 477234 190894 477854 226338
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 446614 481574 482058
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 480954 410614 481574 446058
rect 480954 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 481574 410614
rect 480954 410294 481574 410378
rect 480954 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 481574 410294
rect 480954 374614 481574 410058
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 480954 338614 481574 374058
rect 480954 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 481574 338614
rect 480954 338294 481574 338378
rect 480954 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 481574 338294
rect 480954 302614 481574 338058
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 480954 266614 481574 302058
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 230614 481574 266058
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 480954 194614 481574 230058
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 601174 492134 636618
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 565174 492134 600618
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 491514 457174 492134 492618
rect 491514 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 492134 457174
rect 491514 456854 492134 456938
rect 491514 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 492134 456854
rect 491514 421174 492134 456618
rect 491514 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 492134 421174
rect 491514 420854 492134 420938
rect 491514 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 492134 420854
rect 491514 385174 492134 420618
rect 491514 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 492134 385174
rect 491514 384854 492134 384938
rect 491514 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 492134 384854
rect 491514 349174 492134 384618
rect 491514 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 492134 349174
rect 491514 348854 492134 348938
rect 491514 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 492134 348854
rect 491514 313174 492134 348618
rect 491514 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 492134 313174
rect 491514 312854 492134 312938
rect 491514 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 492134 312854
rect 491514 277174 492134 312618
rect 491514 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 492134 277174
rect 491514 276854 492134 276938
rect 491514 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 492134 276854
rect 491514 241174 492134 276618
rect 491514 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 492134 241174
rect 491514 240854 492134 240938
rect 491514 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 492134 240854
rect 491514 205174 492134 240618
rect 491514 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 492134 205174
rect 491514 204854 492134 204938
rect 491514 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 492134 204854
rect 491514 169174 492134 204618
rect 491514 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 492134 169174
rect 491514 168854 492134 168938
rect 491514 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 492134 168854
rect 491514 133174 492134 168618
rect 491514 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 492134 133174
rect 491514 132854 492134 132938
rect 491514 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 492134 132854
rect 491514 97174 492134 132618
rect 491514 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 492134 97174
rect 491514 96854 492134 96938
rect 491514 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 492134 96854
rect 491514 61174 492134 96618
rect 491514 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 492134 61174
rect 491514 60854 492134 60938
rect 491514 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 492134 60854
rect 491514 25174 492134 60618
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 604894 495854 640338
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 568894 495854 604338
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 532894 495854 568338
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 460894 495854 496338
rect 495234 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 495854 460894
rect 495234 460574 495854 460658
rect 495234 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 495854 460574
rect 495234 424894 495854 460338
rect 495234 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 495854 424894
rect 495234 424574 495854 424658
rect 495234 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 495854 424574
rect 495234 388894 495854 424338
rect 495234 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 495854 388894
rect 495234 388574 495854 388658
rect 495234 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 495854 388574
rect 495234 352894 495854 388338
rect 495234 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 495854 352894
rect 495234 352574 495854 352658
rect 495234 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 495854 352574
rect 495234 316894 495854 352338
rect 495234 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 495854 316894
rect 495234 316574 495854 316658
rect 495234 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 495854 316574
rect 495234 280894 495854 316338
rect 495234 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 495854 280894
rect 495234 280574 495854 280658
rect 495234 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 495854 280574
rect 495234 244894 495854 280338
rect 495234 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 495854 244894
rect 495234 244574 495854 244658
rect 495234 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 495854 244574
rect 495234 208894 495854 244338
rect 495234 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 495854 208894
rect 495234 208574 495854 208658
rect 495234 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 495854 208574
rect 495234 172894 495854 208338
rect 495234 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 495854 172894
rect 495234 172574 495854 172658
rect 495234 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 495854 172574
rect 495234 136894 495854 172338
rect 495234 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 495854 136894
rect 495234 136574 495854 136658
rect 495234 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 495854 136574
rect 495234 100894 495854 136338
rect 495234 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 495854 100894
rect 495234 100574 495854 100658
rect 495234 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 495854 100574
rect 495234 64894 495854 100338
rect 495234 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 495854 64894
rect 495234 64574 495854 64658
rect 495234 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 495854 64574
rect 495234 28894 495854 64338
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 608614 499574 644058
rect 498954 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 499574 608614
rect 498954 608294 499574 608378
rect 498954 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 499574 608294
rect 498954 572614 499574 608058
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 536614 499574 572058
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498954 464614 499574 500058
rect 498954 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 499574 464614
rect 498954 464294 499574 464378
rect 498954 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 499574 464294
rect 498954 428614 499574 464058
rect 498954 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 499574 428614
rect 498954 428294 499574 428378
rect 498954 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 499574 428294
rect 498954 392614 499574 428058
rect 498954 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 499574 392614
rect 498954 392294 499574 392378
rect 498954 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 499574 392294
rect 498954 356614 499574 392058
rect 498954 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 499574 356614
rect 498954 356294 499574 356378
rect 498954 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 499574 356294
rect 498954 320614 499574 356058
rect 498954 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 499574 320614
rect 498954 320294 499574 320378
rect 498954 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 499574 320294
rect 498954 284614 499574 320058
rect 498954 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 499574 284614
rect 498954 284294 499574 284378
rect 498954 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 499574 284294
rect 498954 248614 499574 284058
rect 498954 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 499574 248614
rect 498954 248294 499574 248378
rect 498954 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 499574 248294
rect 498954 212614 499574 248058
rect 498954 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 499574 212614
rect 498954 212294 499574 212378
rect 498954 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 499574 212294
rect 498954 176614 499574 212058
rect 498954 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 499574 176614
rect 498954 176294 499574 176378
rect 498954 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 499574 176294
rect 498954 140614 499574 176058
rect 498954 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 499574 140614
rect 498954 140294 499574 140378
rect 498954 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 499574 140294
rect 498954 104614 499574 140058
rect 498954 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 499574 104614
rect 498954 104294 499574 104378
rect 498954 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 499574 104294
rect 498954 68614 499574 104058
rect 498954 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 499574 68614
rect 498954 68294 499574 68378
rect 498954 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 499574 68294
rect 498954 32614 499574 68058
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509514 295174 510134 330618
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 513234 298894 513854 334338
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 513234 262894 513854 298338
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 516954 302614 517574 338058
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 516954 266614 517574 302058
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 59546 456938 59782 457174
rect 59866 456938 60102 457174
rect 59546 456618 59782 456854
rect 59866 456618 60102 456854
rect 59546 420938 59782 421174
rect 59866 420938 60102 421174
rect 59546 420618 59782 420854
rect 59866 420618 60102 420854
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 59546 384938 59782 385174
rect 59866 384938 60102 385174
rect 59546 384618 59782 384854
rect 59866 384618 60102 384854
rect 59546 348938 59782 349174
rect 59866 348938 60102 349174
rect 59546 348618 59782 348854
rect 59866 348618 60102 348854
rect 59546 312938 59782 313174
rect 59866 312938 60102 313174
rect 59546 312618 59782 312854
rect 59866 312618 60102 312854
rect 59546 276938 59782 277174
rect 59866 276938 60102 277174
rect 59546 276618 59782 276854
rect 59866 276618 60102 276854
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 63266 460658 63502 460894
rect 63586 460658 63822 460894
rect 63266 460338 63502 460574
rect 63586 460338 63822 460574
rect 66986 536378 67222 536614
rect 67306 536378 67542 536614
rect 66986 536058 67222 536294
rect 67306 536058 67542 536294
rect 66986 500378 67222 500614
rect 67306 500378 67542 500614
rect 66986 500058 67222 500294
rect 67306 500058 67542 500294
rect 66986 464378 67222 464614
rect 67306 464378 67542 464614
rect 66986 464058 67222 464294
rect 67306 464058 67542 464294
rect 63266 424658 63502 424894
rect 63586 424658 63822 424894
rect 63266 424338 63502 424574
rect 63586 424338 63822 424574
rect 63266 388658 63502 388894
rect 63586 388658 63822 388894
rect 63266 388338 63502 388574
rect 63586 388338 63822 388574
rect 63266 352658 63502 352894
rect 63586 352658 63822 352894
rect 63266 352338 63502 352574
rect 63586 352338 63822 352574
rect 63266 316658 63502 316894
rect 63586 316658 63822 316894
rect 63266 316338 63502 316574
rect 63586 316338 63822 316574
rect 63266 280658 63502 280894
rect 63586 280658 63822 280894
rect 63266 280338 63502 280574
rect 63586 280338 63822 280574
rect 59546 240938 59782 241174
rect 59866 240938 60102 241174
rect 59546 240618 59782 240854
rect 59866 240618 60102 240854
rect 63266 244658 63502 244894
rect 63586 244658 63822 244894
rect 63266 244338 63502 244574
rect 63586 244338 63822 244574
rect 59546 204938 59782 205174
rect 59866 204938 60102 205174
rect 59546 204618 59782 204854
rect 59866 204618 60102 204854
rect 59546 168938 59782 169174
rect 59866 168938 60102 169174
rect 59546 168618 59782 168854
rect 59866 168618 60102 168854
rect 59546 132938 59782 133174
rect 59866 132938 60102 133174
rect 59546 132618 59782 132854
rect 59866 132618 60102 132854
rect 59546 96938 59782 97174
rect 59866 96938 60102 97174
rect 59546 96618 59782 96854
rect 59866 96618 60102 96854
rect 59546 60938 59782 61174
rect 59866 60938 60102 61174
rect 59546 60618 59782 60854
rect 59866 60618 60102 60854
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 208658 63502 208894
rect 63586 208658 63822 208894
rect 63266 208338 63502 208574
rect 63586 208338 63822 208574
rect 63266 172658 63502 172894
rect 63586 172658 63822 172894
rect 63266 172338 63502 172574
rect 63586 172338 63822 172574
rect 63266 136658 63502 136894
rect 63586 136658 63822 136894
rect 63266 136338 63502 136574
rect 63586 136338 63822 136574
rect 63266 100658 63502 100894
rect 63586 100658 63822 100894
rect 63266 100338 63502 100574
rect 63586 100338 63822 100574
rect 63266 64658 63502 64894
rect 63586 64658 63822 64894
rect 63266 64338 63502 64574
rect 63586 64338 63822 64574
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 73721 543218 73957 543454
rect 73721 542898 73957 543134
rect 66986 356378 67222 356614
rect 67306 356378 67542 356614
rect 66986 356058 67222 356294
rect 67306 356058 67542 356294
rect 66986 320378 67222 320614
rect 67306 320378 67542 320614
rect 66986 320058 67222 320294
rect 67306 320058 67542 320294
rect 66986 212378 67222 212614
rect 67306 212378 67542 212614
rect 66986 212058 67222 212294
rect 67306 212058 67542 212294
rect 66986 176378 67222 176614
rect 67306 176378 67542 176614
rect 66986 176058 67222 176294
rect 67306 176058 67542 176294
rect 66986 140378 67222 140614
rect 67306 140378 67542 140614
rect 66986 140058 67222 140294
rect 67306 140058 67542 140294
rect 73020 399218 73256 399454
rect 73020 398898 73256 399134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 81266 586658 81502 586894
rect 81586 586658 81822 586894
rect 81266 586338 81502 586574
rect 81586 586338 81822 586574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 84986 590378 85222 590614
rect 85306 590378 85542 590614
rect 84986 590058 85222 590294
rect 85306 590058 85542 590294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 77686 561218 77922 561454
rect 77686 560898 77922 561134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 81651 543218 81887 543454
rect 81651 542898 81887 543134
rect 77546 438938 77782 439174
rect 77866 438938 78102 439174
rect 77546 438618 77782 438854
rect 77866 438618 78102 438854
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 85617 561218 85853 561454
rect 85617 560898 85853 561134
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 81266 442658 81502 442894
rect 81586 442658 81822 442894
rect 81266 442338 81502 442574
rect 81586 442338 81822 442574
rect 77546 366938 77782 367174
rect 77866 366938 78102 367174
rect 77546 366618 77782 366854
rect 77866 366618 78102 366854
rect 77546 330938 77782 331174
rect 77866 330938 78102 331174
rect 77546 330618 77782 330854
rect 77866 330618 78102 330854
rect 84986 446378 85222 446614
rect 85306 446378 85542 446614
rect 84986 446058 85222 446294
rect 85306 446058 85542 446294
rect 89582 543218 89818 543454
rect 89582 542898 89818 543134
rect 99266 568658 99502 568894
rect 99586 568658 99822 568894
rect 99266 568338 99502 568574
rect 99586 568338 99822 568574
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 81266 370658 81502 370894
rect 81586 370658 81822 370894
rect 81266 370338 81502 370574
rect 81586 370338 81822 370574
rect 81266 334658 81502 334894
rect 81586 334658 81822 334894
rect 81266 334338 81502 334574
rect 81586 334338 81822 334574
rect 77546 294938 77782 295174
rect 77866 294938 78102 295174
rect 77546 294618 77782 294854
rect 77866 294618 78102 294854
rect 81266 298658 81502 298894
rect 81586 298658 81822 298894
rect 81266 298338 81502 298574
rect 81586 298338 81822 298574
rect 84986 374378 85222 374614
rect 85306 374378 85542 374614
rect 84986 374058 85222 374294
rect 85306 374058 85542 374294
rect 84986 338378 85222 338614
rect 85306 338378 85542 338614
rect 84986 338058 85222 338294
rect 85306 338058 85542 338294
rect 84986 302378 85222 302614
rect 85306 302378 85542 302614
rect 84986 302058 85222 302294
rect 85306 302058 85542 302294
rect 79019 273218 79255 273454
rect 79019 272898 79255 273134
rect 74387 255218 74623 255454
rect 74387 254898 74623 255134
rect 83651 255218 83887 255454
rect 83651 254898 83887 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 77546 222938 77782 223174
rect 77866 222938 78102 223174
rect 77546 222618 77782 222854
rect 77866 222618 78102 222854
rect 77546 186938 77782 187174
rect 77866 186938 78102 187174
rect 77546 186618 77782 186854
rect 77866 186618 78102 186854
rect 77546 150938 77782 151174
rect 77866 150938 78102 151174
rect 77546 150618 77782 150854
rect 77866 150618 78102 150854
rect 88380 417218 88616 417454
rect 88380 416898 88616 417134
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 102986 572378 103222 572614
rect 103306 572378 103542 572614
rect 102986 572058 103222 572294
rect 103306 572058 103542 572294
rect 99266 532658 99502 532894
rect 99586 532658 99822 532894
rect 99266 532338 99502 532574
rect 99586 532338 99822 532574
rect 95546 528938 95782 529174
rect 95866 528938 96102 529174
rect 95546 528618 95782 528854
rect 95866 528618 96102 528854
rect 95546 492938 95782 493174
rect 95866 492938 96102 493174
rect 95546 492618 95782 492854
rect 95866 492618 96102 492854
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 81266 226658 81502 226894
rect 81586 226658 81822 226894
rect 81266 226338 81502 226574
rect 81586 226338 81822 226574
rect 84986 230378 85222 230614
rect 85306 230378 85542 230614
rect 84986 230058 85222 230294
rect 85306 230058 85542 230294
rect 81266 190658 81502 190894
rect 81586 190658 81822 190894
rect 81266 190338 81502 190574
rect 81586 190338 81822 190574
rect 81266 154658 81502 154894
rect 81586 154658 81822 154894
rect 81266 154338 81502 154574
rect 81586 154338 81822 154574
rect 84986 194378 85222 194614
rect 85306 194378 85542 194614
rect 84986 194058 85222 194294
rect 85306 194058 85542 194294
rect 95546 456938 95782 457174
rect 95866 456938 96102 457174
rect 95546 456618 95782 456854
rect 95866 456618 96102 456854
rect 99266 496658 99502 496894
rect 99586 496658 99822 496894
rect 99266 496338 99502 496574
rect 99586 496338 99822 496574
rect 99266 460658 99502 460894
rect 99586 460658 99822 460894
rect 99266 460338 99502 460574
rect 99586 460338 99822 460574
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 88283 273218 88519 273454
rect 88283 272898 88519 273134
rect 84986 158378 85222 158614
rect 85306 158378 85542 158614
rect 84986 158058 85222 158294
rect 85306 158058 85542 158294
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 95546 384938 95782 385174
rect 95866 384938 96102 385174
rect 95546 384618 95782 384854
rect 95866 384618 96102 384854
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 92915 255218 93151 255454
rect 92915 254898 93151 255134
rect 95546 348938 95782 349174
rect 95866 348938 96102 349174
rect 95546 348618 95782 348854
rect 95866 348618 96102 348854
rect 95546 312938 95782 313174
rect 95866 312938 96102 313174
rect 95546 312618 95782 312854
rect 95866 312618 96102 312854
rect 99266 352658 99502 352894
rect 99586 352658 99822 352894
rect 99266 352338 99502 352574
rect 99586 352338 99822 352574
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 102986 536378 103222 536614
rect 103306 536378 103542 536614
rect 102986 536058 103222 536294
rect 103306 536058 103542 536294
rect 102986 500378 103222 500614
rect 103306 500378 103542 500614
rect 102986 500058 103222 500294
rect 103306 500058 103542 500294
rect 102986 464378 103222 464614
rect 103306 464378 103542 464614
rect 102986 464058 103222 464294
rect 103306 464058 103542 464294
rect 103740 399218 103976 399454
rect 103740 398898 103976 399134
rect 102986 356378 103222 356614
rect 103306 356378 103542 356614
rect 102986 356058 103222 356294
rect 103306 356058 103542 356294
rect 99266 316658 99502 316894
rect 99586 316658 99822 316894
rect 99266 316338 99502 316574
rect 99586 316338 99822 316574
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 102986 320378 103222 320614
rect 103306 320378 103542 320614
rect 102986 320058 103222 320294
rect 103306 320058 103542 320294
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 77686 129218 77922 129454
rect 77686 128898 77922 129134
rect 85617 129218 85853 129454
rect 85617 128898 85853 129134
rect 73721 111218 73957 111454
rect 73721 110898 73957 111134
rect 81651 111218 81887 111454
rect 81651 110898 81887 111134
rect 89582 111218 89818 111454
rect 89582 110898 89818 111134
rect 102986 284378 103222 284614
rect 103306 284378 103542 284614
rect 102986 284058 103222 284294
rect 103306 284058 103542 284294
rect 102986 248378 103222 248614
rect 103306 248378 103542 248614
rect 102986 248058 103222 248294
rect 103306 248058 103542 248294
rect 95546 204938 95782 205174
rect 95866 204938 96102 205174
rect 95546 204618 95782 204854
rect 95866 204618 96102 204854
rect 95546 168938 95782 169174
rect 95866 168938 96102 169174
rect 95546 168618 95782 168854
rect 95866 168618 96102 168854
rect 99266 208658 99502 208894
rect 99586 208658 99822 208894
rect 99266 208338 99502 208574
rect 99586 208338 99822 208574
rect 99266 172658 99502 172894
rect 99586 172658 99822 172894
rect 99266 172338 99502 172574
rect 99586 172338 99822 172574
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 113546 438938 113782 439174
rect 113866 438938 114102 439174
rect 113546 438618 113782 438854
rect 113866 438618 114102 438854
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 117266 442658 117502 442894
rect 117586 442658 117822 442894
rect 117266 442338 117502 442574
rect 117586 442338 117822 442574
rect 113546 366938 113782 367174
rect 113866 366938 114102 367174
rect 113546 366618 113782 366854
rect 113866 366618 114102 366854
rect 113546 330938 113782 331174
rect 113866 330938 114102 331174
rect 113546 330618 113782 330854
rect 113866 330618 114102 330854
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 113546 294938 113782 295174
rect 113866 294938 114102 295174
rect 113546 294618 113782 294854
rect 113866 294618 114102 294854
rect 117266 406658 117502 406894
rect 117586 406658 117822 406894
rect 117266 406338 117502 406574
rect 117586 406338 117822 406574
rect 117266 370658 117502 370894
rect 117586 370658 117822 370894
rect 117266 370338 117502 370574
rect 117586 370338 117822 370574
rect 117266 334658 117502 334894
rect 117586 334658 117822 334894
rect 117266 334338 117502 334574
rect 117586 334338 117822 334574
rect 117266 298658 117502 298894
rect 117586 298658 117822 298894
rect 117266 298338 117502 298574
rect 117586 298338 117822 298574
rect 113546 258938 113782 259174
rect 113866 258938 114102 259174
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 102986 212378 103222 212614
rect 103306 212378 103542 212614
rect 102986 212058 103222 212294
rect 103306 212058 103542 212294
rect 113546 258618 113782 258854
rect 113866 258618 114102 258854
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 102986 176378 103222 176614
rect 103306 176378 103542 176614
rect 102986 176058 103222 176294
rect 103306 176058 103542 176294
rect 99266 136658 99502 136894
rect 99586 136658 99822 136894
rect 99266 136338 99502 136574
rect 99586 136338 99822 136574
rect 99266 100658 99502 100894
rect 99586 100658 99822 100894
rect 99266 100338 99502 100574
rect 99586 100338 99822 100574
rect 66986 68378 67222 68614
rect 67306 68378 67542 68614
rect 66986 68058 67222 68294
rect 67306 68058 67542 68294
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 78938 77782 79174
rect 77866 78938 78102 79174
rect 77546 78618 77782 78854
rect 77866 78618 78102 78854
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 82658 81502 82894
rect 81586 82658 81822 82894
rect 81266 82338 81502 82574
rect 81586 82338 81822 82574
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 86378 85222 86614
rect 85306 86378 85542 86614
rect 84986 86058 85222 86294
rect 85306 86058 85542 86294
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 60938 95782 61174
rect 95866 60938 96102 61174
rect 95546 60618 95782 60854
rect 95866 60618 96102 60854
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 102986 140378 103222 140614
rect 103306 140378 103542 140614
rect 102986 140058 103222 140294
rect 103306 140058 103542 140294
rect 102986 104378 103222 104614
rect 103306 104378 103542 104614
rect 102986 104058 103222 104294
rect 103306 104058 103542 104294
rect 99266 64658 99502 64894
rect 99586 64658 99822 64894
rect 99266 64338 99502 64574
rect 99586 64338 99822 64574
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 102986 68378 103222 68614
rect 103306 68378 103542 68614
rect 102986 68058 103222 68294
rect 103306 68058 103542 68294
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 222938 113782 223174
rect 113866 222938 114102 223174
rect 113546 222618 113782 222854
rect 113866 222618 114102 222854
rect 113546 186938 113782 187174
rect 113866 186938 114102 187174
rect 113546 186618 113782 186854
rect 113866 186618 114102 186854
rect 113546 150938 113782 151174
rect 113866 150938 114102 151174
rect 113546 150618 113782 150854
rect 113866 150618 114102 150854
rect 113546 114938 113782 115174
rect 113866 114938 114102 115174
rect 113546 114618 113782 114854
rect 113866 114618 114102 114854
rect 113546 78938 113782 79174
rect 113866 78938 114102 79174
rect 113546 78618 113782 78854
rect 113866 78618 114102 78854
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 262658 117502 262894
rect 117586 262658 117822 262894
rect 117266 262338 117502 262574
rect 117586 262338 117822 262574
rect 117266 226658 117502 226894
rect 117586 226658 117822 226894
rect 117266 226338 117502 226574
rect 117586 226338 117822 226574
rect 117266 190658 117502 190894
rect 117586 190658 117822 190894
rect 117266 190338 117502 190574
rect 117586 190338 117822 190574
rect 117266 154658 117502 154894
rect 117586 154658 117822 154894
rect 117266 154338 117502 154574
rect 117586 154338 117822 154574
rect 117266 118658 117502 118894
rect 117586 118658 117822 118894
rect 117266 118338 117502 118574
rect 117586 118338 117822 118574
rect 117266 82658 117502 82894
rect 117586 82658 117822 82894
rect 117266 82338 117502 82574
rect 117586 82338 117822 82574
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 120986 446378 121222 446614
rect 121306 446378 121542 446614
rect 120986 446058 121222 446294
rect 121306 446058 121542 446294
rect 120986 410378 121222 410614
rect 121306 410378 121542 410614
rect 120986 410058 121222 410294
rect 121306 410058 121542 410294
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 120986 374378 121222 374614
rect 121306 374378 121542 374614
rect 120986 374058 121222 374294
rect 121306 374058 121542 374294
rect 120986 338378 121222 338614
rect 121306 338378 121542 338614
rect 120986 338058 121222 338294
rect 121306 338058 121542 338294
rect 120986 302378 121222 302614
rect 121306 302378 121542 302614
rect 120986 302058 121222 302294
rect 121306 302058 121542 302294
rect 120986 266378 121222 266614
rect 121306 266378 121542 266614
rect 120986 266058 121222 266294
rect 121306 266058 121542 266294
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 120986 230378 121222 230614
rect 121306 230378 121542 230614
rect 120986 230058 121222 230294
rect 121306 230058 121542 230294
rect 120986 194378 121222 194614
rect 121306 194378 121542 194614
rect 120986 194058 121222 194294
rect 121306 194058 121542 194294
rect 120986 158378 121222 158614
rect 121306 158378 121542 158614
rect 120986 158058 121222 158294
rect 121306 158058 121542 158294
rect 120986 122378 121222 122614
rect 121306 122378 121542 122614
rect 120986 122058 121222 122294
rect 121306 122058 121542 122294
rect 120986 86378 121222 86614
rect 121306 86378 121542 86614
rect 120986 86058 121222 86294
rect 121306 86058 121542 86294
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 127826 165218 128062 165454
rect 128146 165218 128382 165454
rect 127826 164898 128062 165134
rect 128146 164898 128382 165134
rect 127826 129218 128062 129454
rect 128146 129218 128382 129454
rect 127826 128898 128062 129134
rect 128146 128898 128382 129134
rect 127826 93218 128062 93454
rect 128146 93218 128382 93454
rect 127826 92898 128062 93134
rect 128146 92898 128382 93134
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 131546 528938 131782 529174
rect 131866 528938 132102 529174
rect 131546 528618 131782 528854
rect 131866 528618 132102 528854
rect 131546 492938 131782 493174
rect 131866 492938 132102 493174
rect 131546 492618 131782 492854
rect 131866 492618 132102 492854
rect 131546 456938 131782 457174
rect 131866 456938 132102 457174
rect 131546 456618 131782 456854
rect 131866 456618 132102 456854
rect 131546 420938 131782 421174
rect 131866 420938 132102 421174
rect 131546 420618 131782 420854
rect 131866 420618 132102 420854
rect 131546 384938 131782 385174
rect 131866 384938 132102 385174
rect 131546 384618 131782 384854
rect 131866 384618 132102 384854
rect 131546 348938 131782 349174
rect 131866 348938 132102 349174
rect 131546 348618 131782 348854
rect 131866 348618 132102 348854
rect 131546 312938 131782 313174
rect 131866 312938 132102 313174
rect 131546 312618 131782 312854
rect 131866 312618 132102 312854
rect 131546 276938 131782 277174
rect 131866 276938 132102 277174
rect 131546 276618 131782 276854
rect 131866 276618 132102 276854
rect 131546 240938 131782 241174
rect 131866 240938 132102 241174
rect 131546 240618 131782 240854
rect 131866 240618 132102 240854
rect 131546 204938 131782 205174
rect 131866 204938 132102 205174
rect 131546 204618 131782 204854
rect 131866 204618 132102 204854
rect 131546 168938 131782 169174
rect 131866 168938 132102 169174
rect 131546 168618 131782 168854
rect 131866 168618 132102 168854
rect 131546 132938 131782 133174
rect 131866 132938 132102 133174
rect 131546 132618 131782 132854
rect 131866 132618 132102 132854
rect 131546 96938 131782 97174
rect 131866 96938 132102 97174
rect 131546 96618 131782 96854
rect 131866 96618 132102 96854
rect 131546 60938 131782 61174
rect 131866 60938 132102 61174
rect 131546 60618 131782 60854
rect 131866 60618 132102 60854
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 135266 532658 135502 532894
rect 135586 532658 135822 532894
rect 135266 532338 135502 532574
rect 135586 532338 135822 532574
rect 135266 496658 135502 496894
rect 135586 496658 135822 496894
rect 135266 496338 135502 496574
rect 135586 496338 135822 496574
rect 135266 460658 135502 460894
rect 135586 460658 135822 460894
rect 135266 460338 135502 460574
rect 135586 460338 135822 460574
rect 135266 424658 135502 424894
rect 135586 424658 135822 424894
rect 135266 424338 135502 424574
rect 135586 424338 135822 424574
rect 135266 388658 135502 388894
rect 135586 388658 135822 388894
rect 135266 388338 135502 388574
rect 135586 388338 135822 388574
rect 135266 352658 135502 352894
rect 135586 352658 135822 352894
rect 135266 352338 135502 352574
rect 135586 352338 135822 352574
rect 135266 316658 135502 316894
rect 135586 316658 135822 316894
rect 135266 316338 135502 316574
rect 135586 316338 135822 316574
rect 135266 280658 135502 280894
rect 135586 280658 135822 280894
rect 135266 280338 135502 280574
rect 135586 280338 135822 280574
rect 135266 244658 135502 244894
rect 135586 244658 135822 244894
rect 135266 244338 135502 244574
rect 135586 244338 135822 244574
rect 135266 208658 135502 208894
rect 135586 208658 135822 208894
rect 135266 208338 135502 208574
rect 135586 208338 135822 208574
rect 135266 172658 135502 172894
rect 135586 172658 135822 172894
rect 135266 172338 135502 172574
rect 135586 172338 135822 172574
rect 135266 136658 135502 136894
rect 135586 136658 135822 136894
rect 135266 136338 135502 136574
rect 135586 136338 135822 136574
rect 135266 100658 135502 100894
rect 135586 100658 135822 100894
rect 135266 100338 135502 100574
rect 135586 100338 135822 100574
rect 135266 64658 135502 64894
rect 135586 64658 135822 64894
rect 135266 64338 135502 64574
rect 135586 64338 135822 64574
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 138986 536378 139222 536614
rect 139306 536378 139542 536614
rect 138986 536058 139222 536294
rect 139306 536058 139542 536294
rect 138986 500378 139222 500614
rect 139306 500378 139542 500614
rect 138986 500058 139222 500294
rect 139306 500058 139542 500294
rect 138986 464378 139222 464614
rect 139306 464378 139542 464614
rect 138986 464058 139222 464294
rect 139306 464058 139542 464294
rect 138986 428378 139222 428614
rect 139306 428378 139542 428614
rect 138986 428058 139222 428294
rect 139306 428058 139542 428294
rect 138986 392378 139222 392614
rect 139306 392378 139542 392614
rect 138986 392058 139222 392294
rect 139306 392058 139542 392294
rect 138986 356378 139222 356614
rect 139306 356378 139542 356614
rect 138986 356058 139222 356294
rect 139306 356058 139542 356294
rect 138986 320378 139222 320614
rect 139306 320378 139542 320614
rect 138986 320058 139222 320294
rect 139306 320058 139542 320294
rect 138986 284378 139222 284614
rect 139306 284378 139542 284614
rect 138986 284058 139222 284294
rect 139306 284058 139542 284294
rect 138986 248378 139222 248614
rect 139306 248378 139542 248614
rect 138986 248058 139222 248294
rect 139306 248058 139542 248294
rect 138986 212378 139222 212614
rect 139306 212378 139542 212614
rect 138986 212058 139222 212294
rect 139306 212058 139542 212294
rect 138986 176378 139222 176614
rect 139306 176378 139542 176614
rect 138986 176058 139222 176294
rect 139306 176058 139542 176294
rect 138986 140378 139222 140614
rect 139306 140378 139542 140614
rect 138986 140058 139222 140294
rect 139306 140058 139542 140294
rect 138986 104378 139222 104614
rect 139306 104378 139542 104614
rect 138986 104058 139222 104294
rect 139306 104058 139542 104294
rect 138986 68378 139222 68614
rect 139306 68378 139542 68614
rect 138986 68058 139222 68294
rect 139306 68058 139542 68294
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 149546 438938 149782 439174
rect 149866 438938 150102 439174
rect 149546 438618 149782 438854
rect 149866 438618 150102 438854
rect 149546 402938 149782 403174
rect 149866 402938 150102 403174
rect 149546 402618 149782 402854
rect 149866 402618 150102 402854
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 149546 330938 149782 331174
rect 149866 330938 150102 331174
rect 149546 330618 149782 330854
rect 149866 330618 150102 330854
rect 149546 294938 149782 295174
rect 149866 294938 150102 295174
rect 149546 294618 149782 294854
rect 149866 294618 150102 294854
rect 149546 258938 149782 259174
rect 149866 258938 150102 259174
rect 149546 258618 149782 258854
rect 149866 258618 150102 258854
rect 149546 222938 149782 223174
rect 149866 222938 150102 223174
rect 149546 222618 149782 222854
rect 149866 222618 150102 222854
rect 149546 186938 149782 187174
rect 149866 186938 150102 187174
rect 149546 186618 149782 186854
rect 149866 186618 150102 186854
rect 149546 150938 149782 151174
rect 149866 150938 150102 151174
rect 149546 150618 149782 150854
rect 149866 150618 150102 150854
rect 149546 114938 149782 115174
rect 149866 114938 150102 115174
rect 149546 114618 149782 114854
rect 149866 114618 150102 114854
rect 149546 78938 149782 79174
rect 149866 78938 150102 79174
rect 149546 78618 149782 78854
rect 149866 78618 150102 78854
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 153266 514658 153502 514894
rect 153586 514658 153822 514894
rect 153266 514338 153502 514574
rect 153586 514338 153822 514574
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 153266 442658 153502 442894
rect 153586 442658 153822 442894
rect 153266 442338 153502 442574
rect 153586 442338 153822 442574
rect 153266 406658 153502 406894
rect 153586 406658 153822 406894
rect 153266 406338 153502 406574
rect 153586 406338 153822 406574
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 153266 334658 153502 334894
rect 153586 334658 153822 334894
rect 153266 334338 153502 334574
rect 153586 334338 153822 334574
rect 153266 298658 153502 298894
rect 153586 298658 153822 298894
rect 153266 298338 153502 298574
rect 153586 298338 153822 298574
rect 153266 262658 153502 262894
rect 153586 262658 153822 262894
rect 153266 262338 153502 262574
rect 153586 262338 153822 262574
rect 153266 226658 153502 226894
rect 153586 226658 153822 226894
rect 153266 226338 153502 226574
rect 153586 226338 153822 226574
rect 153266 190658 153502 190894
rect 153586 190658 153822 190894
rect 153266 190338 153502 190574
rect 153586 190338 153822 190574
rect 153266 154658 153502 154894
rect 153586 154658 153822 154894
rect 153266 154338 153502 154574
rect 153586 154338 153822 154574
rect 153266 118658 153502 118894
rect 153586 118658 153822 118894
rect 153266 118338 153502 118574
rect 153586 118338 153822 118574
rect 153266 82658 153502 82894
rect 153586 82658 153822 82894
rect 153266 82338 153502 82574
rect 153586 82338 153822 82574
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 156986 518378 157222 518614
rect 157306 518378 157542 518614
rect 156986 518058 157222 518294
rect 157306 518058 157542 518294
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 156986 446378 157222 446614
rect 157306 446378 157542 446614
rect 156986 446058 157222 446294
rect 157306 446058 157542 446294
rect 156986 410378 157222 410614
rect 157306 410378 157542 410614
rect 156986 410058 157222 410294
rect 157306 410058 157542 410294
rect 156986 374378 157222 374614
rect 157306 374378 157542 374614
rect 156986 374058 157222 374294
rect 157306 374058 157542 374294
rect 156986 338378 157222 338614
rect 157306 338378 157542 338614
rect 156986 338058 157222 338294
rect 157306 338058 157542 338294
rect 156986 302378 157222 302614
rect 157306 302378 157542 302614
rect 156986 302058 157222 302294
rect 157306 302058 157542 302294
rect 156986 266378 157222 266614
rect 157306 266378 157542 266614
rect 156986 266058 157222 266294
rect 157306 266058 157542 266294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 156986 230378 157222 230614
rect 157306 230378 157542 230614
rect 156986 230058 157222 230294
rect 157306 230058 157542 230294
rect 156986 194378 157222 194614
rect 157306 194378 157542 194614
rect 156986 194058 157222 194294
rect 157306 194058 157542 194294
rect 156986 158378 157222 158614
rect 157306 158378 157542 158614
rect 156986 158058 157222 158294
rect 157306 158058 157542 158294
rect 156986 122378 157222 122614
rect 157306 122378 157542 122614
rect 156986 122058 157222 122294
rect 157306 122058 157542 122294
rect 156986 86378 157222 86614
rect 157306 86378 157542 86614
rect 156986 86058 157222 86294
rect 157306 86058 157542 86294
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 163826 165218 164062 165454
rect 164146 165218 164382 165454
rect 163826 164898 164062 165134
rect 164146 164898 164382 165134
rect 163826 129218 164062 129454
rect 164146 129218 164382 129454
rect 163826 128898 164062 129134
rect 164146 128898 164382 129134
rect 163826 93218 164062 93454
rect 164146 93218 164382 93454
rect 163826 92898 164062 93134
rect 164146 92898 164382 93134
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 167546 528938 167782 529174
rect 167866 528938 168102 529174
rect 167546 528618 167782 528854
rect 167866 528618 168102 528854
rect 167546 492938 167782 493174
rect 167866 492938 168102 493174
rect 167546 492618 167782 492854
rect 167866 492618 168102 492854
rect 167546 456938 167782 457174
rect 167866 456938 168102 457174
rect 167546 456618 167782 456854
rect 167866 456618 168102 456854
rect 167546 420938 167782 421174
rect 167866 420938 168102 421174
rect 167546 420618 167782 420854
rect 167866 420618 168102 420854
rect 167546 384938 167782 385174
rect 167866 384938 168102 385174
rect 167546 384618 167782 384854
rect 167866 384618 168102 384854
rect 167546 348938 167782 349174
rect 167866 348938 168102 349174
rect 167546 348618 167782 348854
rect 167866 348618 168102 348854
rect 167546 312938 167782 313174
rect 167866 312938 168102 313174
rect 167546 312618 167782 312854
rect 167866 312618 168102 312854
rect 167546 276938 167782 277174
rect 167866 276938 168102 277174
rect 167546 276618 167782 276854
rect 167866 276618 168102 276854
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 171266 532658 171502 532894
rect 171586 532658 171822 532894
rect 171266 532338 171502 532574
rect 171586 532338 171822 532574
rect 171266 496658 171502 496894
rect 171586 496658 171822 496894
rect 171266 496338 171502 496574
rect 171586 496338 171822 496574
rect 171266 460658 171502 460894
rect 171586 460658 171822 460894
rect 171266 460338 171502 460574
rect 171586 460338 171822 460574
rect 171266 424658 171502 424894
rect 171586 424658 171822 424894
rect 171266 424338 171502 424574
rect 171586 424338 171822 424574
rect 171266 388658 171502 388894
rect 171586 388658 171822 388894
rect 171266 388338 171502 388574
rect 171586 388338 171822 388574
rect 171266 352658 171502 352894
rect 171586 352658 171822 352894
rect 171266 352338 171502 352574
rect 171586 352338 171822 352574
rect 171266 316658 171502 316894
rect 171586 316658 171822 316894
rect 171266 316338 171502 316574
rect 171586 316338 171822 316574
rect 171266 280658 171502 280894
rect 171586 280658 171822 280894
rect 171266 280338 171502 280574
rect 171586 280338 171822 280574
rect 171266 244658 171502 244894
rect 171586 244658 171822 244894
rect 171266 244338 171502 244574
rect 171586 244338 171822 244574
rect 167546 240938 167782 241174
rect 167866 240938 168102 241174
rect 167546 240618 167782 240854
rect 167866 240618 168102 240854
rect 167546 204938 167782 205174
rect 167866 204938 168102 205174
rect 167546 204618 167782 204854
rect 167866 204618 168102 204854
rect 167546 168938 167782 169174
rect 167866 168938 168102 169174
rect 167546 168618 167782 168854
rect 167866 168618 168102 168854
rect 167546 132938 167782 133174
rect 167866 132938 168102 133174
rect 167546 132618 167782 132854
rect 167866 132618 168102 132854
rect 167546 96938 167782 97174
rect 167866 96938 168102 97174
rect 167546 96618 167782 96854
rect 167866 96618 168102 96854
rect 167546 60938 167782 61174
rect 167866 60938 168102 61174
rect 167546 60618 167782 60854
rect 167866 60618 168102 60854
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 171266 208658 171502 208894
rect 171586 208658 171822 208894
rect 171266 208338 171502 208574
rect 171586 208338 171822 208574
rect 171266 172658 171502 172894
rect 171586 172658 171822 172894
rect 171266 172338 171502 172574
rect 171586 172338 171822 172574
rect 171266 136658 171502 136894
rect 171586 136658 171822 136894
rect 171266 136338 171502 136574
rect 171586 136338 171822 136574
rect 171266 100658 171502 100894
rect 171586 100658 171822 100894
rect 171266 100338 171502 100574
rect 171586 100338 171822 100574
rect 171266 64658 171502 64894
rect 171586 64658 171822 64894
rect 171266 64338 171502 64574
rect 171586 64338 171822 64574
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 174986 536378 175222 536614
rect 175306 536378 175542 536614
rect 174986 536058 175222 536294
rect 175306 536058 175542 536294
rect 174986 500378 175222 500614
rect 175306 500378 175542 500614
rect 174986 500058 175222 500294
rect 175306 500058 175542 500294
rect 174986 464378 175222 464614
rect 175306 464378 175542 464614
rect 174986 464058 175222 464294
rect 175306 464058 175542 464294
rect 174986 428378 175222 428614
rect 175306 428378 175542 428614
rect 174986 428058 175222 428294
rect 175306 428058 175542 428294
rect 174986 392378 175222 392614
rect 175306 392378 175542 392614
rect 174986 392058 175222 392294
rect 175306 392058 175542 392294
rect 174986 356378 175222 356614
rect 175306 356378 175542 356614
rect 174986 356058 175222 356294
rect 175306 356058 175542 356294
rect 174986 320378 175222 320614
rect 175306 320378 175542 320614
rect 174986 320058 175222 320294
rect 175306 320058 175542 320294
rect 174986 284378 175222 284614
rect 175306 284378 175542 284614
rect 174986 284058 175222 284294
rect 175306 284058 175542 284294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 174986 248378 175222 248614
rect 175306 248378 175542 248614
rect 174986 248058 175222 248294
rect 175306 248058 175542 248294
rect 174986 212378 175222 212614
rect 175306 212378 175542 212614
rect 174986 212058 175222 212294
rect 175306 212058 175542 212294
rect 174986 176378 175222 176614
rect 175306 176378 175542 176614
rect 174986 176058 175222 176294
rect 175306 176058 175542 176294
rect 174986 140378 175222 140614
rect 175306 140378 175542 140614
rect 174986 140058 175222 140294
rect 175306 140058 175542 140294
rect 174986 104378 175222 104614
rect 175306 104378 175542 104614
rect 174986 104058 175222 104294
rect 175306 104058 175542 104294
rect 174986 68378 175222 68614
rect 175306 68378 175542 68614
rect 174986 68058 175222 68294
rect 175306 68058 175542 68294
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 185546 438938 185782 439174
rect 185866 438938 186102 439174
rect 185546 438618 185782 438854
rect 185866 438618 186102 438854
rect 185546 402938 185782 403174
rect 185866 402938 186102 403174
rect 185546 402618 185782 402854
rect 185866 402618 186102 402854
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 185546 330938 185782 331174
rect 185866 330938 186102 331174
rect 185546 330618 185782 330854
rect 185866 330618 186102 330854
rect 185546 294938 185782 295174
rect 185866 294938 186102 295174
rect 185546 294618 185782 294854
rect 185866 294618 186102 294854
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 189266 442658 189502 442894
rect 189586 442658 189822 442894
rect 189266 442338 189502 442574
rect 189586 442338 189822 442574
rect 189266 406658 189502 406894
rect 189586 406658 189822 406894
rect 189266 406338 189502 406574
rect 189586 406338 189822 406574
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 189266 334658 189502 334894
rect 189586 334658 189822 334894
rect 189266 334338 189502 334574
rect 189586 334338 189822 334574
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 192986 518378 193222 518614
rect 193306 518378 193542 518614
rect 192986 518058 193222 518294
rect 193306 518058 193542 518294
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 192986 446378 193222 446614
rect 193306 446378 193542 446614
rect 192986 446058 193222 446294
rect 193306 446058 193542 446294
rect 192986 410378 193222 410614
rect 193306 410378 193542 410614
rect 192986 410058 193222 410294
rect 193306 410058 193542 410294
rect 192986 374378 193222 374614
rect 193306 374378 193542 374614
rect 192986 374058 193222 374294
rect 193306 374058 193542 374294
rect 192986 338378 193222 338614
rect 193306 338378 193542 338614
rect 192986 338058 193222 338294
rect 193306 338058 193542 338294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 203546 528938 203782 529174
rect 203866 528938 204102 529174
rect 203546 528618 203782 528854
rect 203866 528618 204102 528854
rect 203546 492938 203782 493174
rect 203866 492938 204102 493174
rect 203546 492618 203782 492854
rect 203866 492618 204102 492854
rect 203546 456938 203782 457174
rect 203866 456938 204102 457174
rect 203546 456618 203782 456854
rect 203866 456618 204102 456854
rect 203546 420938 203782 421174
rect 203866 420938 204102 421174
rect 203546 420618 203782 420854
rect 203866 420618 204102 420854
rect 203546 384938 203782 385174
rect 203866 384938 204102 385174
rect 203546 384618 203782 384854
rect 203866 384618 204102 384854
rect 203546 348938 203782 349174
rect 203866 348938 204102 349174
rect 203546 348618 203782 348854
rect 203866 348618 204102 348854
rect 203546 312938 203782 313174
rect 203866 312938 204102 313174
rect 203546 312618 203782 312854
rect 203866 312618 204102 312854
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 189266 298658 189502 298894
rect 189586 298658 189822 298894
rect 189266 298338 189502 298574
rect 189586 298338 189822 298574
rect 189266 262658 189502 262894
rect 189586 262658 189822 262894
rect 189266 262338 189502 262574
rect 189586 262338 189822 262574
rect 185546 222938 185782 223174
rect 185866 222938 186102 223174
rect 185546 222618 185782 222854
rect 185866 222618 186102 222854
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 189266 226658 189502 226894
rect 189586 226658 189822 226894
rect 189266 226338 189502 226574
rect 189586 226338 189822 226574
rect 185546 186938 185782 187174
rect 185866 186938 186102 187174
rect 185546 186618 185782 186854
rect 185866 186618 186102 186854
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 185546 114938 185782 115174
rect 185866 114938 186102 115174
rect 185546 114618 185782 114854
rect 185866 114618 186102 114854
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 189266 190658 189502 190894
rect 189586 190658 189822 190894
rect 189266 190338 189502 190574
rect 189586 190338 189822 190574
rect 189266 154658 189502 154894
rect 189586 154658 189822 154894
rect 189266 154338 189502 154574
rect 189586 154338 189822 154574
rect 189266 118658 189502 118894
rect 189586 118658 189822 118894
rect 189266 118338 189502 118574
rect 189586 118338 189822 118574
rect 185546 78938 185782 79174
rect 185866 78938 186102 79174
rect 185546 78618 185782 78854
rect 185866 78618 186102 78854
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 192986 230378 193222 230614
rect 193306 230378 193542 230614
rect 192986 230058 193222 230294
rect 193306 230058 193542 230294
rect 192986 194378 193222 194614
rect 193306 194378 193542 194614
rect 192986 194058 193222 194294
rect 193306 194058 193542 194294
rect 192986 158378 193222 158614
rect 193306 158378 193542 158614
rect 192986 158058 193222 158294
rect 193306 158058 193542 158294
rect 189266 82658 189502 82894
rect 189586 82658 189822 82894
rect 189266 82338 189502 82574
rect 189586 82338 189822 82574
rect 197818 291218 198054 291454
rect 197818 290898 198054 291134
rect 197818 255218 198054 255454
rect 197818 254898 198054 255134
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 207266 532658 207502 532894
rect 207586 532658 207822 532894
rect 207266 532338 207502 532574
rect 207586 532338 207822 532574
rect 207266 496658 207502 496894
rect 207586 496658 207822 496894
rect 207266 496338 207502 496574
rect 207586 496338 207822 496574
rect 207266 460658 207502 460894
rect 207586 460658 207822 460894
rect 207266 460338 207502 460574
rect 207586 460338 207822 460574
rect 207266 424658 207502 424894
rect 207586 424658 207822 424894
rect 207266 424338 207502 424574
rect 207586 424338 207822 424574
rect 207266 388658 207502 388894
rect 207586 388658 207822 388894
rect 207266 388338 207502 388574
rect 207586 388338 207822 388574
rect 207266 352658 207502 352894
rect 207586 352658 207822 352894
rect 207266 352338 207502 352574
rect 207586 352338 207822 352574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 210986 536378 211222 536614
rect 211306 536378 211542 536614
rect 210986 536058 211222 536294
rect 211306 536058 211542 536294
rect 210986 500378 211222 500614
rect 211306 500378 211542 500614
rect 210986 500058 211222 500294
rect 211306 500058 211542 500294
rect 210986 464378 211222 464614
rect 211306 464378 211542 464614
rect 210986 464058 211222 464294
rect 211306 464058 211542 464294
rect 210986 428378 211222 428614
rect 211306 428378 211542 428614
rect 210986 428058 211222 428294
rect 211306 428058 211542 428294
rect 210986 392378 211222 392614
rect 211306 392378 211542 392614
rect 210986 392058 211222 392294
rect 211306 392058 211542 392294
rect 210986 356378 211222 356614
rect 211306 356378 211542 356614
rect 210986 356058 211222 356294
rect 211306 356058 211542 356294
rect 210986 320378 211222 320614
rect 211306 320378 211542 320614
rect 207266 316658 207502 316894
rect 207586 316658 207822 316894
rect 207266 316338 207502 316574
rect 207586 316338 207822 316574
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 192986 86378 193222 86614
rect 193306 86378 193542 86614
rect 192986 86058 193222 86294
rect 193306 86058 193542 86294
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 199430 111218 199666 111454
rect 199430 110898 199666 111134
rect 203546 204938 203782 205174
rect 203866 204938 204102 205174
rect 203546 204618 203782 204854
rect 203866 204618 204102 204854
rect 207266 208658 207502 208894
rect 207586 208658 207822 208894
rect 207266 208338 207502 208574
rect 207586 208338 207822 208574
rect 203546 168938 203782 169174
rect 203866 168938 204102 169174
rect 203546 168618 203782 168854
rect 203866 168618 204102 168854
rect 204306 129218 204542 129454
rect 204306 128898 204542 129134
rect 210986 320058 211222 320294
rect 211306 320058 211542 320294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 221546 510938 221782 511174
rect 221866 510938 222102 511174
rect 221546 510618 221782 510854
rect 221866 510618 222102 510854
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 221546 438938 221782 439174
rect 221866 438938 222102 439174
rect 221546 438618 221782 438854
rect 221866 438618 222102 438854
rect 221546 402938 221782 403174
rect 221866 402938 222102 403174
rect 221546 402618 221782 402854
rect 221866 402618 222102 402854
rect 221546 366938 221782 367174
rect 221866 366938 222102 367174
rect 221546 366618 221782 366854
rect 221866 366618 222102 366854
rect 221546 330938 221782 331174
rect 221866 330938 222102 331174
rect 221546 330618 221782 330854
rect 221866 330618 222102 330854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 225266 514658 225502 514894
rect 225586 514658 225822 514894
rect 225266 514338 225502 514574
rect 225586 514338 225822 514574
rect 225266 478658 225502 478894
rect 225586 478658 225822 478894
rect 225266 478338 225502 478574
rect 225586 478338 225822 478574
rect 225266 442658 225502 442894
rect 225586 442658 225822 442894
rect 225266 442338 225502 442574
rect 225586 442338 225822 442574
rect 225266 406658 225502 406894
rect 225586 406658 225822 406894
rect 225266 406338 225502 406574
rect 225586 406338 225822 406574
rect 225266 370658 225502 370894
rect 225586 370658 225822 370894
rect 225266 370338 225502 370574
rect 225586 370338 225822 370574
rect 225266 334658 225502 334894
rect 225586 334658 225822 334894
rect 225266 334338 225502 334574
rect 225586 334338 225822 334574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 228986 518378 229222 518614
rect 229306 518378 229542 518614
rect 228986 518058 229222 518294
rect 229306 518058 229542 518294
rect 228986 482378 229222 482614
rect 229306 482378 229542 482614
rect 228986 482058 229222 482294
rect 229306 482058 229542 482294
rect 228986 446378 229222 446614
rect 229306 446378 229542 446614
rect 228986 446058 229222 446294
rect 229306 446058 229542 446294
rect 228986 410378 229222 410614
rect 229306 410378 229542 410614
rect 228986 410058 229222 410294
rect 229306 410058 229542 410294
rect 228986 374378 229222 374614
rect 229306 374378 229542 374614
rect 228986 374058 229222 374294
rect 229306 374058 229542 374294
rect 228986 338378 229222 338614
rect 229306 338378 229542 338614
rect 228986 338058 229222 338294
rect 229306 338058 229542 338294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 239546 600938 239782 601174
rect 239866 600938 240102 601174
rect 239546 600618 239782 600854
rect 239866 600618 240102 600854
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 239546 528938 239782 529174
rect 239866 528938 240102 529174
rect 239546 528618 239782 528854
rect 239866 528618 240102 528854
rect 239546 492938 239782 493174
rect 239866 492938 240102 493174
rect 239546 492618 239782 492854
rect 239866 492618 240102 492854
rect 239546 456938 239782 457174
rect 239866 456938 240102 457174
rect 239546 456618 239782 456854
rect 239866 456618 240102 456854
rect 239546 420938 239782 421174
rect 239866 420938 240102 421174
rect 239546 420618 239782 420854
rect 239866 420618 240102 420854
rect 239546 384938 239782 385174
rect 239866 384938 240102 385174
rect 239546 384618 239782 384854
rect 239866 384618 240102 384854
rect 239546 348938 239782 349174
rect 239866 348938 240102 349174
rect 239546 348618 239782 348854
rect 239866 348618 240102 348854
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 243266 604658 243502 604894
rect 243586 604658 243822 604894
rect 243266 604338 243502 604574
rect 243586 604338 243822 604574
rect 243266 568658 243502 568894
rect 243586 568658 243822 568894
rect 243266 568338 243502 568574
rect 243586 568338 243822 568574
rect 243266 532658 243502 532894
rect 243586 532658 243822 532894
rect 243266 532338 243502 532574
rect 243586 532338 243822 532574
rect 243266 496658 243502 496894
rect 243586 496658 243822 496894
rect 243266 496338 243502 496574
rect 243586 496338 243822 496574
rect 243266 460658 243502 460894
rect 243586 460658 243822 460894
rect 243266 460338 243502 460574
rect 243586 460338 243822 460574
rect 243266 424658 243502 424894
rect 243586 424658 243822 424894
rect 243266 424338 243502 424574
rect 243586 424338 243822 424574
rect 243266 388658 243502 388894
rect 243586 388658 243822 388894
rect 243266 388338 243502 388574
rect 243586 388338 243822 388574
rect 243266 352658 243502 352894
rect 243586 352658 243822 352894
rect 243266 352338 243502 352574
rect 243586 352338 243822 352574
rect 239546 312938 239782 313174
rect 239866 312938 240102 313174
rect 239546 312618 239782 312854
rect 239866 312618 240102 312854
rect 207266 172658 207502 172894
rect 207586 172658 207822 172894
rect 207266 172338 207502 172574
rect 207586 172338 207822 172574
rect 209182 111218 209418 111454
rect 209182 110898 209418 111134
rect 210986 212378 211222 212614
rect 211306 212378 211542 212614
rect 210986 212058 211222 212294
rect 211306 212058 211542 212294
rect 210986 176378 211222 176614
rect 211306 176378 211542 176614
rect 210986 176058 211222 176294
rect 211306 176058 211542 176294
rect 213178 273218 213414 273454
rect 213178 272898 213414 273134
rect 214058 129218 214294 129454
rect 214058 128898 214294 129134
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 221546 222938 221782 223174
rect 221866 222938 222102 223174
rect 221546 222618 221782 222854
rect 221866 222618 222102 222854
rect 221546 186938 221782 187174
rect 221866 186938 222102 187174
rect 221546 186618 221782 186854
rect 221866 186618 222102 186854
rect 221546 150938 221782 151174
rect 221866 150938 222102 151174
rect 221546 150618 221782 150854
rect 221866 150618 222102 150854
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 225266 226658 225502 226894
rect 225586 226658 225822 226894
rect 225266 226338 225502 226574
rect 225586 226338 225822 226574
rect 228538 291218 228774 291454
rect 228538 290898 228774 291134
rect 228538 255218 228774 255454
rect 228538 254898 228774 255134
rect 225266 190658 225502 190894
rect 225586 190658 225822 190894
rect 225266 190338 225502 190574
rect 225586 190338 225822 190574
rect 225266 154658 225502 154894
rect 225586 154658 225822 154894
rect 225266 154338 225502 154574
rect 225586 154338 225822 154574
rect 218934 111218 219170 111454
rect 218934 110898 219170 111134
rect 228986 230378 229222 230614
rect 229306 230378 229542 230614
rect 228986 230058 229222 230294
rect 229306 230058 229542 230294
rect 228986 194378 229222 194614
rect 229306 194378 229542 194614
rect 228986 194058 229222 194294
rect 229306 194058 229542 194294
rect 228986 158378 229222 158614
rect 229306 158378 229542 158614
rect 228986 158058 229222 158294
rect 229306 158058 229542 158294
rect 228986 122378 229222 122614
rect 229306 122378 229542 122614
rect 228986 122058 229222 122294
rect 229306 122058 229542 122294
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 60938 203782 61174
rect 203866 60938 204102 61174
rect 203546 60618 203782 60854
rect 203866 60618 204102 60854
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 64658 207502 64894
rect 207586 64658 207822 64894
rect 207266 64338 207502 64574
rect 207586 64338 207822 64574
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 210986 68378 211222 68614
rect 211306 68378 211542 68614
rect 210986 68058 211222 68294
rect 211306 68058 211542 68294
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 228986 86378 229222 86614
rect 229306 86378 229542 86614
rect 228986 86058 229222 86294
rect 229306 86058 229542 86294
rect 225266 82658 225502 82894
rect 225586 82658 225822 82894
rect 225266 82338 225502 82574
rect 225586 82338 225822 82574
rect 221546 78938 221782 79174
rect 221866 78938 222102 79174
rect 221546 78618 221782 78854
rect 221866 78618 222102 78854
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 243266 316658 243502 316894
rect 243586 316658 243822 316894
rect 243266 316338 243502 316574
rect 243586 316338 243822 316574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 246986 608378 247222 608614
rect 247306 608378 247542 608614
rect 246986 608058 247222 608294
rect 247306 608058 247542 608294
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 246986 536378 247222 536614
rect 247306 536378 247542 536614
rect 246986 536058 247222 536294
rect 247306 536058 247542 536294
rect 246986 500378 247222 500614
rect 247306 500378 247542 500614
rect 246986 500058 247222 500294
rect 247306 500058 247542 500294
rect 246986 464378 247222 464614
rect 247306 464378 247542 464614
rect 246986 464058 247222 464294
rect 247306 464058 247542 464294
rect 246986 428378 247222 428614
rect 247306 428378 247542 428614
rect 246986 428058 247222 428294
rect 247306 428058 247542 428294
rect 246986 392378 247222 392614
rect 247306 392378 247542 392614
rect 246986 392058 247222 392294
rect 247306 392058 247542 392294
rect 246986 356378 247222 356614
rect 247306 356378 247542 356614
rect 246986 356058 247222 356294
rect 247306 356058 247542 356294
rect 246986 320378 247222 320614
rect 247306 320378 247542 320614
rect 246986 320058 247222 320294
rect 247306 320058 247542 320294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 239546 204938 239782 205174
rect 239866 204938 240102 205174
rect 239546 204618 239782 204854
rect 239866 204618 240102 204854
rect 239546 168938 239782 169174
rect 239866 168938 240102 169174
rect 239546 168618 239782 168854
rect 239866 168618 240102 168854
rect 239546 132938 239782 133174
rect 239866 132938 240102 133174
rect 239546 132618 239782 132854
rect 239866 132618 240102 132854
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 243898 273218 244134 273454
rect 243898 272898 244134 273134
rect 243266 208658 243502 208894
rect 243586 208658 243822 208894
rect 243266 208338 243502 208574
rect 243586 208338 243822 208574
rect 243266 172658 243502 172894
rect 243586 172658 243822 172894
rect 243266 172338 243502 172574
rect 243586 172338 243822 172574
rect 246986 212378 247222 212614
rect 247306 212378 247542 212614
rect 246986 212058 247222 212294
rect 247306 212058 247542 212294
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 257546 510938 257782 511174
rect 257866 510938 258102 511174
rect 257546 510618 257782 510854
rect 257866 510618 258102 510854
rect 257546 474938 257782 475174
rect 257866 474938 258102 475174
rect 257546 474618 257782 474854
rect 257866 474618 258102 474854
rect 257546 438938 257782 439174
rect 257866 438938 258102 439174
rect 257546 438618 257782 438854
rect 257866 438618 258102 438854
rect 257546 402938 257782 403174
rect 257866 402938 258102 403174
rect 257546 402618 257782 402854
rect 257866 402618 258102 402854
rect 257546 366938 257782 367174
rect 257866 366938 258102 367174
rect 257546 366618 257782 366854
rect 257866 366618 258102 366854
rect 257546 330938 257782 331174
rect 257866 330938 258102 331174
rect 257546 330618 257782 330854
rect 257866 330618 258102 330854
rect 246986 176378 247222 176614
rect 247306 176378 247542 176614
rect 246986 176058 247222 176294
rect 247306 176058 247542 176294
rect 243266 136658 243502 136894
rect 243586 136658 243822 136894
rect 243266 136338 243502 136574
rect 243586 136338 243822 136574
rect 239546 96938 239782 97174
rect 239866 96938 240102 97174
rect 239546 96618 239782 96854
rect 239866 96618 240102 96854
rect 239546 60938 239782 61174
rect 239866 60938 240102 61174
rect 239546 60618 239782 60854
rect 239866 60618 240102 60854
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 100658 243502 100894
rect 243586 100658 243822 100894
rect 243266 100338 243502 100574
rect 243586 100338 243822 100574
rect 243266 64658 243502 64894
rect 243586 64658 243822 64894
rect 243266 64338 243502 64574
rect 243586 64338 243822 64574
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 261266 514658 261502 514894
rect 261586 514658 261822 514894
rect 261266 514338 261502 514574
rect 261586 514338 261822 514574
rect 261266 478658 261502 478894
rect 261586 478658 261822 478894
rect 261266 478338 261502 478574
rect 261586 478338 261822 478574
rect 261266 442658 261502 442894
rect 261586 442658 261822 442894
rect 261266 442338 261502 442574
rect 261586 442338 261822 442574
rect 261266 406658 261502 406894
rect 261586 406658 261822 406894
rect 261266 406338 261502 406574
rect 261586 406338 261822 406574
rect 261266 370658 261502 370894
rect 261586 370658 261822 370894
rect 261266 370338 261502 370574
rect 261586 370338 261822 370574
rect 261266 334658 261502 334894
rect 261586 334658 261822 334894
rect 261266 334338 261502 334574
rect 261586 334338 261822 334574
rect 257546 294938 257782 295174
rect 257866 294938 258102 295174
rect 257546 294618 257782 294854
rect 257866 294618 258102 294854
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 257546 258938 257782 259174
rect 257866 258938 258102 259174
rect 257546 258618 257782 258854
rect 257866 258618 258102 258854
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 264986 518378 265222 518614
rect 265306 518378 265542 518614
rect 264986 518058 265222 518294
rect 265306 518058 265542 518294
rect 264986 482378 265222 482614
rect 265306 482378 265542 482614
rect 264986 482058 265222 482294
rect 265306 482058 265542 482294
rect 264986 446378 265222 446614
rect 265306 446378 265542 446614
rect 264986 446058 265222 446294
rect 265306 446058 265542 446294
rect 264986 410378 265222 410614
rect 265306 410378 265542 410614
rect 264986 410058 265222 410294
rect 265306 410058 265542 410294
rect 264986 374378 265222 374614
rect 265306 374378 265542 374614
rect 264986 374058 265222 374294
rect 265306 374058 265542 374294
rect 264986 338378 265222 338614
rect 265306 338378 265542 338614
rect 264986 338058 265222 338294
rect 265306 338058 265542 338294
rect 261266 298658 261502 298894
rect 261586 298658 261822 298894
rect 261266 298338 261502 298574
rect 261586 298338 261822 298574
rect 261266 262658 261502 262894
rect 261586 262658 261822 262894
rect 261266 262338 261502 262574
rect 261586 262338 261822 262574
rect 264986 302378 265222 302614
rect 265306 302378 265542 302614
rect 264986 302058 265222 302294
rect 265306 302058 265542 302294
rect 264986 266378 265222 266614
rect 265306 266378 265542 266614
rect 264986 266058 265222 266294
rect 265306 266058 265542 266294
rect 261266 226658 261502 226894
rect 261586 226658 261822 226894
rect 261266 226338 261502 226574
rect 261586 226338 261822 226574
rect 257546 222938 257782 223174
rect 257866 222938 258102 223174
rect 257546 222618 257782 222854
rect 257866 222618 258102 222854
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 246986 140378 247222 140614
rect 247306 140378 247542 140614
rect 246986 140058 247222 140294
rect 247306 140058 247542 140294
rect 246986 104378 247222 104614
rect 247306 104378 247542 104614
rect 246986 104058 247222 104294
rect 247306 104058 247542 104294
rect 246986 68378 247222 68614
rect 247306 68378 247542 68614
rect 246986 68058 247222 68294
rect 247306 68058 247542 68294
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 186938 257782 187174
rect 257866 186938 258102 187174
rect 257546 186618 257782 186854
rect 257866 186618 258102 186854
rect 257546 150938 257782 151174
rect 257866 150938 258102 151174
rect 257546 150618 257782 150854
rect 257866 150618 258102 150854
rect 257546 114938 257782 115174
rect 257866 114938 258102 115174
rect 257546 114618 257782 114854
rect 257866 114618 258102 114854
rect 257546 78938 257782 79174
rect 257866 78938 258102 79174
rect 257546 78618 257782 78854
rect 257866 78618 258102 78854
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 275546 600938 275782 601174
rect 275866 600938 276102 601174
rect 275546 600618 275782 600854
rect 275866 600618 276102 600854
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 275546 528938 275782 529174
rect 275866 528938 276102 529174
rect 275546 528618 275782 528854
rect 275866 528618 276102 528854
rect 275546 492938 275782 493174
rect 275866 492938 276102 493174
rect 275546 492618 275782 492854
rect 275866 492618 276102 492854
rect 275546 456938 275782 457174
rect 275866 456938 276102 457174
rect 275546 456618 275782 456854
rect 275866 456618 276102 456854
rect 275546 420938 275782 421174
rect 275866 420938 276102 421174
rect 275546 420618 275782 420854
rect 275866 420618 276102 420854
rect 275546 384938 275782 385174
rect 275866 384938 276102 385174
rect 275546 384618 275782 384854
rect 275866 384618 276102 384854
rect 275546 348938 275782 349174
rect 275866 348938 276102 349174
rect 275546 348618 275782 348854
rect 275866 348618 276102 348854
rect 275546 312938 275782 313174
rect 275866 312938 276102 313174
rect 275546 312618 275782 312854
rect 275866 312618 276102 312854
rect 275546 276938 275782 277174
rect 275866 276938 276102 277174
rect 275546 276618 275782 276854
rect 275866 276618 276102 276854
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 264986 230378 265222 230614
rect 265306 230378 265542 230614
rect 264986 230058 265222 230294
rect 265306 230058 265542 230294
rect 261266 190658 261502 190894
rect 261586 190658 261822 190894
rect 261266 190338 261502 190574
rect 261586 190338 261822 190574
rect 261266 154658 261502 154894
rect 261586 154658 261822 154894
rect 261266 154338 261502 154574
rect 261586 154338 261822 154574
rect 261266 118658 261502 118894
rect 261586 118658 261822 118894
rect 261266 118338 261502 118574
rect 261586 118338 261822 118574
rect 261266 82658 261502 82894
rect 261586 82658 261822 82894
rect 261266 82338 261502 82574
rect 261586 82338 261822 82574
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 194378 265222 194614
rect 265306 194378 265542 194614
rect 264986 194058 265222 194294
rect 265306 194058 265542 194294
rect 264986 158378 265222 158614
rect 265306 158378 265542 158614
rect 264986 158058 265222 158294
rect 265306 158058 265542 158294
rect 264986 122378 265222 122614
rect 265306 122378 265542 122614
rect 264986 122058 265222 122294
rect 265306 122058 265542 122294
rect 264986 86378 265222 86614
rect 265306 86378 265542 86614
rect 264986 86058 265222 86294
rect 265306 86058 265542 86294
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 275546 240938 275782 241174
rect 275866 240938 276102 241174
rect 275546 240618 275782 240854
rect 275866 240618 276102 240854
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 204938 275782 205174
rect 275866 204938 276102 205174
rect 275546 204618 275782 204854
rect 275866 204618 276102 204854
rect 275546 168938 275782 169174
rect 275866 168938 276102 169174
rect 275546 168618 275782 168854
rect 275866 168618 276102 168854
rect 275546 132938 275782 133174
rect 275866 132938 276102 133174
rect 275546 132618 275782 132854
rect 275866 132618 276102 132854
rect 275546 96938 275782 97174
rect 275866 96938 276102 97174
rect 275546 96618 275782 96854
rect 275866 96618 276102 96854
rect 275546 60938 275782 61174
rect 275866 60938 276102 61174
rect 275546 60618 275782 60854
rect 275866 60618 276102 60854
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 279266 604658 279502 604894
rect 279586 604658 279822 604894
rect 279266 604338 279502 604574
rect 279586 604338 279822 604574
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 279266 532658 279502 532894
rect 279586 532658 279822 532894
rect 279266 532338 279502 532574
rect 279586 532338 279822 532574
rect 279266 496658 279502 496894
rect 279586 496658 279822 496894
rect 279266 496338 279502 496574
rect 279586 496338 279822 496574
rect 279266 460658 279502 460894
rect 279586 460658 279822 460894
rect 279266 460338 279502 460574
rect 279586 460338 279822 460574
rect 279266 424658 279502 424894
rect 279586 424658 279822 424894
rect 279266 424338 279502 424574
rect 279586 424338 279822 424574
rect 279266 388658 279502 388894
rect 279586 388658 279822 388894
rect 279266 388338 279502 388574
rect 279586 388338 279822 388574
rect 279266 352658 279502 352894
rect 279586 352658 279822 352894
rect 279266 352338 279502 352574
rect 279586 352338 279822 352574
rect 279266 316658 279502 316894
rect 279586 316658 279822 316894
rect 279266 316338 279502 316574
rect 279586 316338 279822 316574
rect 279266 280658 279502 280894
rect 279586 280658 279822 280894
rect 279266 280338 279502 280574
rect 279586 280338 279822 280574
rect 279266 244658 279502 244894
rect 279586 244658 279822 244894
rect 279266 244338 279502 244574
rect 279586 244338 279822 244574
rect 279266 208658 279502 208894
rect 279586 208658 279822 208894
rect 279266 208338 279502 208574
rect 279586 208338 279822 208574
rect 279266 172658 279502 172894
rect 279586 172658 279822 172894
rect 279266 172338 279502 172574
rect 279586 172338 279822 172574
rect 279266 136658 279502 136894
rect 279586 136658 279822 136894
rect 279266 136338 279502 136574
rect 279586 136338 279822 136574
rect 279266 100658 279502 100894
rect 279586 100658 279822 100894
rect 279266 100338 279502 100574
rect 279586 100338 279822 100574
rect 279266 64658 279502 64894
rect 279586 64658 279822 64894
rect 279266 64338 279502 64574
rect 279586 64338 279822 64574
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 282986 608378 283222 608614
rect 283306 608378 283542 608614
rect 282986 608058 283222 608294
rect 283306 608058 283542 608294
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 282986 536378 283222 536614
rect 283306 536378 283542 536614
rect 282986 536058 283222 536294
rect 283306 536058 283542 536294
rect 282986 500378 283222 500614
rect 283306 500378 283542 500614
rect 282986 500058 283222 500294
rect 283306 500058 283542 500294
rect 282986 464378 283222 464614
rect 283306 464378 283542 464614
rect 282986 464058 283222 464294
rect 283306 464058 283542 464294
rect 282986 428378 283222 428614
rect 283306 428378 283542 428614
rect 282986 428058 283222 428294
rect 283306 428058 283542 428294
rect 282986 392378 283222 392614
rect 283306 392378 283542 392614
rect 282986 392058 283222 392294
rect 283306 392058 283542 392294
rect 282986 356378 283222 356614
rect 283306 356378 283542 356614
rect 282986 356058 283222 356294
rect 283306 356058 283542 356294
rect 282986 320378 283222 320614
rect 283306 320378 283542 320614
rect 282986 320058 283222 320294
rect 283306 320058 283542 320294
rect 282986 284378 283222 284614
rect 283306 284378 283542 284614
rect 282986 284058 283222 284294
rect 283306 284058 283542 284294
rect 282986 248378 283222 248614
rect 283306 248378 283542 248614
rect 282986 248058 283222 248294
rect 283306 248058 283542 248294
rect 282986 212378 283222 212614
rect 283306 212378 283542 212614
rect 282986 212058 283222 212294
rect 283306 212058 283542 212294
rect 282986 176378 283222 176614
rect 283306 176378 283542 176614
rect 282986 176058 283222 176294
rect 283306 176058 283542 176294
rect 282986 140378 283222 140614
rect 283306 140378 283542 140614
rect 282986 140058 283222 140294
rect 283306 140058 283542 140294
rect 282986 104378 283222 104614
rect 283306 104378 283542 104614
rect 282986 104058 283222 104294
rect 283306 104058 283542 104294
rect 282986 68378 283222 68614
rect 283306 68378 283542 68614
rect 282986 68058 283222 68294
rect 283306 68058 283542 68294
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 293546 510938 293782 511174
rect 293866 510938 294102 511174
rect 293546 510618 293782 510854
rect 293866 510618 294102 510854
rect 293546 474938 293782 475174
rect 293866 474938 294102 475174
rect 293546 474618 293782 474854
rect 293866 474618 294102 474854
rect 293546 438938 293782 439174
rect 293866 438938 294102 439174
rect 293546 438618 293782 438854
rect 293866 438618 294102 438854
rect 293546 402938 293782 403174
rect 293866 402938 294102 403174
rect 293546 402618 293782 402854
rect 293866 402618 294102 402854
rect 293546 366938 293782 367174
rect 293866 366938 294102 367174
rect 293546 366618 293782 366854
rect 293866 366618 294102 366854
rect 293546 330938 293782 331174
rect 293866 330938 294102 331174
rect 293546 330618 293782 330854
rect 293866 330618 294102 330854
rect 293546 294938 293782 295174
rect 293866 294938 294102 295174
rect 293546 294618 293782 294854
rect 293866 294618 294102 294854
rect 293546 258938 293782 259174
rect 293866 258938 294102 259174
rect 293546 258618 293782 258854
rect 293866 258618 294102 258854
rect 293546 222938 293782 223174
rect 293866 222938 294102 223174
rect 293546 222618 293782 222854
rect 293866 222618 294102 222854
rect 293546 186938 293782 187174
rect 293866 186938 294102 187174
rect 293546 186618 293782 186854
rect 293866 186618 294102 186854
rect 293546 150938 293782 151174
rect 293866 150938 294102 151174
rect 293546 150618 293782 150854
rect 293866 150618 294102 150854
rect 293546 114938 293782 115174
rect 293866 114938 294102 115174
rect 293546 114618 293782 114854
rect 293866 114618 294102 114854
rect 293546 78938 293782 79174
rect 293866 78938 294102 79174
rect 293546 78618 293782 78854
rect 293866 78618 294102 78854
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 297266 514658 297502 514894
rect 297586 514658 297822 514894
rect 297266 514338 297502 514574
rect 297586 514338 297822 514574
rect 297266 478658 297502 478894
rect 297586 478658 297822 478894
rect 297266 478338 297502 478574
rect 297586 478338 297822 478574
rect 297266 442658 297502 442894
rect 297586 442658 297822 442894
rect 297266 442338 297502 442574
rect 297586 442338 297822 442574
rect 297266 406658 297502 406894
rect 297586 406658 297822 406894
rect 297266 406338 297502 406574
rect 297586 406338 297822 406574
rect 297266 370658 297502 370894
rect 297586 370658 297822 370894
rect 297266 370338 297502 370574
rect 297586 370338 297822 370574
rect 297266 334658 297502 334894
rect 297586 334658 297822 334894
rect 297266 334338 297502 334574
rect 297586 334338 297822 334574
rect 297266 298658 297502 298894
rect 297586 298658 297822 298894
rect 297266 298338 297502 298574
rect 297586 298338 297822 298574
rect 297266 262658 297502 262894
rect 297586 262658 297822 262894
rect 297266 262338 297502 262574
rect 297586 262338 297822 262574
rect 297266 226658 297502 226894
rect 297586 226658 297822 226894
rect 297266 226338 297502 226574
rect 297586 226338 297822 226574
rect 297266 190658 297502 190894
rect 297586 190658 297822 190894
rect 297266 190338 297502 190574
rect 297586 190338 297822 190574
rect 297266 154658 297502 154894
rect 297586 154658 297822 154894
rect 297266 154338 297502 154574
rect 297586 154338 297822 154574
rect 297266 118658 297502 118894
rect 297586 118658 297822 118894
rect 297266 118338 297502 118574
rect 297586 118338 297822 118574
rect 297266 82658 297502 82894
rect 297586 82658 297822 82894
rect 297266 82338 297502 82574
rect 297586 82338 297822 82574
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 300986 518378 301222 518614
rect 301306 518378 301542 518614
rect 300986 518058 301222 518294
rect 301306 518058 301542 518294
rect 300986 482378 301222 482614
rect 301306 482378 301542 482614
rect 300986 482058 301222 482294
rect 301306 482058 301542 482294
rect 300986 446378 301222 446614
rect 301306 446378 301542 446614
rect 300986 446058 301222 446294
rect 301306 446058 301542 446294
rect 300986 410378 301222 410614
rect 301306 410378 301542 410614
rect 300986 410058 301222 410294
rect 301306 410058 301542 410294
rect 300986 374378 301222 374614
rect 301306 374378 301542 374614
rect 300986 374058 301222 374294
rect 301306 374058 301542 374294
rect 300986 338378 301222 338614
rect 301306 338378 301542 338614
rect 300986 338058 301222 338294
rect 301306 338058 301542 338294
rect 300986 302378 301222 302614
rect 301306 302378 301542 302614
rect 300986 302058 301222 302294
rect 301306 302058 301542 302294
rect 300986 266378 301222 266614
rect 301306 266378 301542 266614
rect 300986 266058 301222 266294
rect 301306 266058 301542 266294
rect 300986 230378 301222 230614
rect 301306 230378 301542 230614
rect 300986 230058 301222 230294
rect 301306 230058 301542 230294
rect 300986 194378 301222 194614
rect 301306 194378 301542 194614
rect 300986 194058 301222 194294
rect 301306 194058 301542 194294
rect 300986 158378 301222 158614
rect 301306 158378 301542 158614
rect 300986 158058 301222 158294
rect 301306 158058 301542 158294
rect 300986 122378 301222 122614
rect 301306 122378 301542 122614
rect 300986 122058 301222 122294
rect 301306 122058 301542 122294
rect 300986 86378 301222 86614
rect 301306 86378 301542 86614
rect 300986 86058 301222 86294
rect 301306 86058 301542 86294
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 311546 528938 311782 529174
rect 311866 528938 312102 529174
rect 311546 528618 311782 528854
rect 311866 528618 312102 528854
rect 311546 492938 311782 493174
rect 311866 492938 312102 493174
rect 311546 492618 311782 492854
rect 311866 492618 312102 492854
rect 311546 456938 311782 457174
rect 311866 456938 312102 457174
rect 311546 456618 311782 456854
rect 311866 456618 312102 456854
rect 311546 420938 311782 421174
rect 311866 420938 312102 421174
rect 311546 420618 311782 420854
rect 311866 420618 312102 420854
rect 311546 384938 311782 385174
rect 311866 384938 312102 385174
rect 311546 384618 311782 384854
rect 311866 384618 312102 384854
rect 311546 348938 311782 349174
rect 311866 348938 312102 349174
rect 311546 348618 311782 348854
rect 311866 348618 312102 348854
rect 311546 312938 311782 313174
rect 311866 312938 312102 313174
rect 311546 312618 311782 312854
rect 311866 312618 312102 312854
rect 311546 276938 311782 277174
rect 311866 276938 312102 277174
rect 311546 276618 311782 276854
rect 311866 276618 312102 276854
rect 311546 240938 311782 241174
rect 311866 240938 312102 241174
rect 311546 240618 311782 240854
rect 311866 240618 312102 240854
rect 311546 204938 311782 205174
rect 311866 204938 312102 205174
rect 311546 204618 311782 204854
rect 311866 204618 312102 204854
rect 311546 168938 311782 169174
rect 311866 168938 312102 169174
rect 311546 168618 311782 168854
rect 311866 168618 312102 168854
rect 311546 132938 311782 133174
rect 311866 132938 312102 133174
rect 311546 132618 311782 132854
rect 311866 132618 312102 132854
rect 311546 96938 311782 97174
rect 311866 96938 312102 97174
rect 311546 96618 311782 96854
rect 311866 96618 312102 96854
rect 311546 60938 311782 61174
rect 311866 60938 312102 61174
rect 311546 60618 311782 60854
rect 311866 60618 312102 60854
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 315266 532658 315502 532894
rect 315586 532658 315822 532894
rect 315266 532338 315502 532574
rect 315586 532338 315822 532574
rect 315266 496658 315502 496894
rect 315586 496658 315822 496894
rect 315266 496338 315502 496574
rect 315586 496338 315822 496574
rect 315266 460658 315502 460894
rect 315586 460658 315822 460894
rect 315266 460338 315502 460574
rect 315586 460338 315822 460574
rect 315266 424658 315502 424894
rect 315586 424658 315822 424894
rect 315266 424338 315502 424574
rect 315586 424338 315822 424574
rect 315266 388658 315502 388894
rect 315586 388658 315822 388894
rect 315266 388338 315502 388574
rect 315586 388338 315822 388574
rect 315266 352658 315502 352894
rect 315586 352658 315822 352894
rect 315266 352338 315502 352574
rect 315586 352338 315822 352574
rect 315266 316658 315502 316894
rect 315586 316658 315822 316894
rect 315266 316338 315502 316574
rect 315586 316338 315822 316574
rect 315266 280658 315502 280894
rect 315586 280658 315822 280894
rect 315266 280338 315502 280574
rect 315586 280338 315822 280574
rect 315266 244658 315502 244894
rect 315586 244658 315822 244894
rect 315266 244338 315502 244574
rect 315586 244338 315822 244574
rect 315266 208658 315502 208894
rect 315586 208658 315822 208894
rect 315266 208338 315502 208574
rect 315586 208338 315822 208574
rect 315266 172658 315502 172894
rect 315586 172658 315822 172894
rect 315266 172338 315502 172574
rect 315586 172338 315822 172574
rect 315266 136658 315502 136894
rect 315586 136658 315822 136894
rect 315266 136338 315502 136574
rect 315586 136338 315822 136574
rect 315266 100658 315502 100894
rect 315586 100658 315822 100894
rect 315266 100338 315502 100574
rect 315586 100338 315822 100574
rect 315266 64658 315502 64894
rect 315586 64658 315822 64894
rect 315266 64338 315502 64574
rect 315586 64338 315822 64574
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 318986 536378 319222 536614
rect 319306 536378 319542 536614
rect 318986 536058 319222 536294
rect 319306 536058 319542 536294
rect 318986 500378 319222 500614
rect 319306 500378 319542 500614
rect 318986 500058 319222 500294
rect 319306 500058 319542 500294
rect 318986 464378 319222 464614
rect 319306 464378 319542 464614
rect 318986 464058 319222 464294
rect 319306 464058 319542 464294
rect 318986 428378 319222 428614
rect 319306 428378 319542 428614
rect 318986 428058 319222 428294
rect 319306 428058 319542 428294
rect 318986 392378 319222 392614
rect 319306 392378 319542 392614
rect 318986 392058 319222 392294
rect 319306 392058 319542 392294
rect 318986 356378 319222 356614
rect 319306 356378 319542 356614
rect 318986 356058 319222 356294
rect 319306 356058 319542 356294
rect 318986 320378 319222 320614
rect 319306 320378 319542 320614
rect 318986 320058 319222 320294
rect 319306 320058 319542 320294
rect 318986 284378 319222 284614
rect 319306 284378 319542 284614
rect 318986 284058 319222 284294
rect 319306 284058 319542 284294
rect 318986 248378 319222 248614
rect 319306 248378 319542 248614
rect 318986 248058 319222 248294
rect 319306 248058 319542 248294
rect 318986 212378 319222 212614
rect 319306 212378 319542 212614
rect 318986 212058 319222 212294
rect 319306 212058 319542 212294
rect 318986 176378 319222 176614
rect 319306 176378 319542 176614
rect 318986 176058 319222 176294
rect 319306 176058 319542 176294
rect 318986 140378 319222 140614
rect 319306 140378 319542 140614
rect 318986 140058 319222 140294
rect 319306 140058 319542 140294
rect 318986 104378 319222 104614
rect 319306 104378 319542 104614
rect 318986 104058 319222 104294
rect 319306 104058 319542 104294
rect 318986 68378 319222 68614
rect 319306 68378 319542 68614
rect 318986 68058 319222 68294
rect 319306 68058 319542 68294
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 329546 546938 329782 547174
rect 329866 546938 330102 547174
rect 329546 546618 329782 546854
rect 329866 546618 330102 546854
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 329546 474938 329782 475174
rect 329866 474938 330102 475174
rect 329546 474618 329782 474854
rect 329866 474618 330102 474854
rect 329546 438938 329782 439174
rect 329866 438938 330102 439174
rect 329546 438618 329782 438854
rect 329866 438618 330102 438854
rect 329546 402938 329782 403174
rect 329866 402938 330102 403174
rect 329546 402618 329782 402854
rect 329866 402618 330102 402854
rect 329546 366938 329782 367174
rect 329866 366938 330102 367174
rect 329546 366618 329782 366854
rect 329866 366618 330102 366854
rect 329546 330938 329782 331174
rect 329866 330938 330102 331174
rect 329546 330618 329782 330854
rect 329866 330618 330102 330854
rect 329546 294938 329782 295174
rect 329866 294938 330102 295174
rect 329546 294618 329782 294854
rect 329866 294618 330102 294854
rect 329546 258938 329782 259174
rect 329866 258938 330102 259174
rect 329546 258618 329782 258854
rect 329866 258618 330102 258854
rect 329546 222938 329782 223174
rect 329866 222938 330102 223174
rect 329546 222618 329782 222854
rect 329866 222618 330102 222854
rect 329546 186938 329782 187174
rect 329866 186938 330102 187174
rect 329546 186618 329782 186854
rect 329866 186618 330102 186854
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 329546 114938 329782 115174
rect 329866 114938 330102 115174
rect 329546 114618 329782 114854
rect 329866 114618 330102 114854
rect 329546 78938 329782 79174
rect 329866 78938 330102 79174
rect 329546 78618 329782 78854
rect 329866 78618 330102 78854
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 333266 550658 333502 550894
rect 333586 550658 333822 550894
rect 333266 550338 333502 550574
rect 333586 550338 333822 550574
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 333266 478658 333502 478894
rect 333586 478658 333822 478894
rect 333266 478338 333502 478574
rect 333586 478338 333822 478574
rect 333266 442658 333502 442894
rect 333586 442658 333822 442894
rect 333266 442338 333502 442574
rect 333586 442338 333822 442574
rect 333266 406658 333502 406894
rect 333586 406658 333822 406894
rect 333266 406338 333502 406574
rect 333586 406338 333822 406574
rect 333266 370658 333502 370894
rect 333586 370658 333822 370894
rect 333266 370338 333502 370574
rect 333586 370338 333822 370574
rect 333266 334658 333502 334894
rect 333586 334658 333822 334894
rect 333266 334338 333502 334574
rect 333586 334338 333822 334574
rect 333266 298658 333502 298894
rect 333586 298658 333822 298894
rect 333266 298338 333502 298574
rect 333586 298338 333822 298574
rect 333266 262658 333502 262894
rect 333586 262658 333822 262894
rect 333266 262338 333502 262574
rect 333586 262338 333822 262574
rect 333266 226658 333502 226894
rect 333586 226658 333822 226894
rect 333266 226338 333502 226574
rect 333586 226338 333822 226574
rect 333266 190658 333502 190894
rect 333586 190658 333822 190894
rect 333266 190338 333502 190574
rect 333586 190338 333822 190574
rect 333266 154658 333502 154894
rect 333586 154658 333822 154894
rect 333266 154338 333502 154574
rect 333586 154338 333822 154574
rect 333266 118658 333502 118894
rect 333586 118658 333822 118894
rect 333266 118338 333502 118574
rect 333586 118338 333822 118574
rect 333266 82658 333502 82894
rect 333586 82658 333822 82894
rect 333266 82338 333502 82574
rect 333586 82338 333822 82574
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 336986 518378 337222 518614
rect 337306 518378 337542 518614
rect 336986 518058 337222 518294
rect 337306 518058 337542 518294
rect 336986 482378 337222 482614
rect 337306 482378 337542 482614
rect 336986 482058 337222 482294
rect 337306 482058 337542 482294
rect 336986 446378 337222 446614
rect 337306 446378 337542 446614
rect 336986 446058 337222 446294
rect 337306 446058 337542 446294
rect 336986 410378 337222 410614
rect 337306 410378 337542 410614
rect 336986 410058 337222 410294
rect 337306 410058 337542 410294
rect 336986 374378 337222 374614
rect 337306 374378 337542 374614
rect 336986 374058 337222 374294
rect 337306 374058 337542 374294
rect 336986 338378 337222 338614
rect 337306 338378 337542 338614
rect 336986 338058 337222 338294
rect 337306 338058 337542 338294
rect 336986 302378 337222 302614
rect 337306 302378 337542 302614
rect 336986 302058 337222 302294
rect 337306 302058 337542 302294
rect 336986 266378 337222 266614
rect 337306 266378 337542 266614
rect 336986 266058 337222 266294
rect 337306 266058 337542 266294
rect 336986 230378 337222 230614
rect 337306 230378 337542 230614
rect 336986 230058 337222 230294
rect 337306 230058 337542 230294
rect 336986 194378 337222 194614
rect 337306 194378 337542 194614
rect 336986 194058 337222 194294
rect 337306 194058 337542 194294
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 336986 122378 337222 122614
rect 337306 122378 337542 122614
rect 336986 122058 337222 122294
rect 337306 122058 337542 122294
rect 336986 86378 337222 86614
rect 337306 86378 337542 86614
rect 336986 86058 337222 86294
rect 337306 86058 337542 86294
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 347546 564938 347782 565174
rect 347866 564938 348102 565174
rect 347546 564618 347782 564854
rect 347866 564618 348102 564854
rect 347546 528938 347782 529174
rect 347866 528938 348102 529174
rect 347546 528618 347782 528854
rect 347866 528618 348102 528854
rect 347546 492938 347782 493174
rect 347866 492938 348102 493174
rect 347546 492618 347782 492854
rect 347866 492618 348102 492854
rect 347546 456938 347782 457174
rect 347866 456938 348102 457174
rect 347546 456618 347782 456854
rect 347866 456618 348102 456854
rect 347546 420938 347782 421174
rect 347866 420938 348102 421174
rect 347546 420618 347782 420854
rect 347866 420618 348102 420854
rect 347546 384938 347782 385174
rect 347866 384938 348102 385174
rect 347546 384618 347782 384854
rect 347866 384618 348102 384854
rect 347546 348938 347782 349174
rect 347866 348938 348102 349174
rect 347546 348618 347782 348854
rect 347866 348618 348102 348854
rect 347546 312938 347782 313174
rect 347866 312938 348102 313174
rect 347546 312618 347782 312854
rect 347866 312618 348102 312854
rect 347546 276938 347782 277174
rect 347866 276938 348102 277174
rect 347546 276618 347782 276854
rect 347866 276618 348102 276854
rect 347546 240938 347782 241174
rect 347866 240938 348102 241174
rect 347546 240618 347782 240854
rect 347866 240618 348102 240854
rect 347546 204938 347782 205174
rect 347866 204938 348102 205174
rect 347546 204618 347782 204854
rect 347866 204618 348102 204854
rect 347546 168938 347782 169174
rect 347866 168938 348102 169174
rect 347546 168618 347782 168854
rect 347866 168618 348102 168854
rect 347546 132938 347782 133174
rect 347866 132938 348102 133174
rect 347546 132618 347782 132854
rect 347866 132618 348102 132854
rect 347546 96938 347782 97174
rect 347866 96938 348102 97174
rect 347546 96618 347782 96854
rect 347866 96618 348102 96854
rect 347546 60938 347782 61174
rect 347866 60938 348102 61174
rect 347546 60618 347782 60854
rect 347866 60618 348102 60854
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 351266 568658 351502 568894
rect 351586 568658 351822 568894
rect 351266 568338 351502 568574
rect 351586 568338 351822 568574
rect 351266 532658 351502 532894
rect 351586 532658 351822 532894
rect 351266 532338 351502 532574
rect 351586 532338 351822 532574
rect 351266 496658 351502 496894
rect 351586 496658 351822 496894
rect 351266 496338 351502 496574
rect 351586 496338 351822 496574
rect 351266 460658 351502 460894
rect 351586 460658 351822 460894
rect 351266 460338 351502 460574
rect 351586 460338 351822 460574
rect 351266 424658 351502 424894
rect 351586 424658 351822 424894
rect 351266 424338 351502 424574
rect 351586 424338 351822 424574
rect 351266 388658 351502 388894
rect 351586 388658 351822 388894
rect 351266 388338 351502 388574
rect 351586 388338 351822 388574
rect 351266 352658 351502 352894
rect 351586 352658 351822 352894
rect 351266 352338 351502 352574
rect 351586 352338 351822 352574
rect 351266 316658 351502 316894
rect 351586 316658 351822 316894
rect 351266 316338 351502 316574
rect 351586 316338 351822 316574
rect 351266 280658 351502 280894
rect 351586 280658 351822 280894
rect 351266 280338 351502 280574
rect 351586 280338 351822 280574
rect 351266 244658 351502 244894
rect 351586 244658 351822 244894
rect 351266 244338 351502 244574
rect 351586 244338 351822 244574
rect 351266 208658 351502 208894
rect 351586 208658 351822 208894
rect 351266 208338 351502 208574
rect 351586 208338 351822 208574
rect 351266 172658 351502 172894
rect 351586 172658 351822 172894
rect 351266 172338 351502 172574
rect 351586 172338 351822 172574
rect 351266 136658 351502 136894
rect 351586 136658 351822 136894
rect 351266 136338 351502 136574
rect 351586 136338 351822 136574
rect 351266 100658 351502 100894
rect 351586 100658 351822 100894
rect 351266 100338 351502 100574
rect 351586 100338 351822 100574
rect 351266 64658 351502 64894
rect 351586 64658 351822 64894
rect 351266 64338 351502 64574
rect 351586 64338 351822 64574
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 354986 536378 355222 536614
rect 355306 536378 355542 536614
rect 354986 536058 355222 536294
rect 355306 536058 355542 536294
rect 354986 500378 355222 500614
rect 355306 500378 355542 500614
rect 354986 500058 355222 500294
rect 355306 500058 355542 500294
rect 354986 464378 355222 464614
rect 355306 464378 355542 464614
rect 354986 464058 355222 464294
rect 355306 464058 355542 464294
rect 354986 428378 355222 428614
rect 355306 428378 355542 428614
rect 354986 428058 355222 428294
rect 355306 428058 355542 428294
rect 354986 392378 355222 392614
rect 355306 392378 355542 392614
rect 354986 392058 355222 392294
rect 355306 392058 355542 392294
rect 354986 356378 355222 356614
rect 355306 356378 355542 356614
rect 354986 356058 355222 356294
rect 355306 356058 355542 356294
rect 354986 320378 355222 320614
rect 355306 320378 355542 320614
rect 354986 320058 355222 320294
rect 355306 320058 355542 320294
rect 354986 284378 355222 284614
rect 355306 284378 355542 284614
rect 354986 284058 355222 284294
rect 355306 284058 355542 284294
rect 354986 248378 355222 248614
rect 355306 248378 355542 248614
rect 354986 248058 355222 248294
rect 355306 248058 355542 248294
rect 354986 212378 355222 212614
rect 355306 212378 355542 212614
rect 354986 212058 355222 212294
rect 355306 212058 355542 212294
rect 354986 176378 355222 176614
rect 355306 176378 355542 176614
rect 354986 176058 355222 176294
rect 355306 176058 355542 176294
rect 354986 140378 355222 140614
rect 355306 140378 355542 140614
rect 354986 140058 355222 140294
rect 355306 140058 355542 140294
rect 354986 104378 355222 104614
rect 355306 104378 355542 104614
rect 354986 104058 355222 104294
rect 355306 104058 355542 104294
rect 354986 68378 355222 68614
rect 355306 68378 355542 68614
rect 354986 68058 355222 68294
rect 355306 68058 355542 68294
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 365546 366938 365782 367174
rect 365866 366938 366102 367174
rect 365546 366618 365782 366854
rect 365866 366618 366102 366854
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 365546 294938 365782 295174
rect 365866 294938 366102 295174
rect 365546 294618 365782 294854
rect 365866 294618 366102 294854
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 369266 298658 369502 298894
rect 369586 298658 369822 298894
rect 369266 298338 369502 298574
rect 369586 298338 369822 298574
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 369266 226658 369502 226894
rect 369586 226658 369822 226894
rect 369266 226338 369502 226574
rect 369586 226338 369822 226574
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 383546 564938 383782 565174
rect 383866 564938 384102 565174
rect 383546 564618 383782 564854
rect 383866 564618 384102 564854
rect 383546 528938 383782 529174
rect 383866 528938 384102 529174
rect 383546 528618 383782 528854
rect 383866 528618 384102 528854
rect 383546 492938 383782 493174
rect 383866 492938 384102 493174
rect 383546 492618 383782 492854
rect 383866 492618 384102 492854
rect 383546 456938 383782 457174
rect 383866 456938 384102 457174
rect 383546 456618 383782 456854
rect 383866 456618 384102 456854
rect 383546 420938 383782 421174
rect 383866 420938 384102 421174
rect 383546 420618 383782 420854
rect 383866 420618 384102 420854
rect 383546 384938 383782 385174
rect 383866 384938 384102 385174
rect 383546 384618 383782 384854
rect 383866 384618 384102 384854
rect 383546 348938 383782 349174
rect 383866 348938 384102 349174
rect 383546 348618 383782 348854
rect 383866 348618 384102 348854
rect 383546 312938 383782 313174
rect 383866 312938 384102 313174
rect 383546 312618 383782 312854
rect 383866 312618 384102 312854
rect 383546 276938 383782 277174
rect 383866 276938 384102 277174
rect 383546 276618 383782 276854
rect 383866 276618 384102 276854
rect 383546 240938 383782 241174
rect 383866 240938 384102 241174
rect 383546 240618 383782 240854
rect 383866 240618 384102 240854
rect 383546 204938 383782 205174
rect 383866 204938 384102 205174
rect 383546 204618 383782 204854
rect 383866 204618 384102 204854
rect 383546 168938 383782 169174
rect 383866 168938 384102 169174
rect 383546 168618 383782 168854
rect 383866 168618 384102 168854
rect 383546 132938 383782 133174
rect 383866 132938 384102 133174
rect 383546 132618 383782 132854
rect 383866 132618 384102 132854
rect 383546 96938 383782 97174
rect 383866 96938 384102 97174
rect 383546 96618 383782 96854
rect 383866 96618 384102 96854
rect 383546 60938 383782 61174
rect 383866 60938 384102 61174
rect 383546 60618 383782 60854
rect 383866 60618 384102 60854
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 387266 568658 387502 568894
rect 387586 568658 387822 568894
rect 387266 568338 387502 568574
rect 387586 568338 387822 568574
rect 387266 532658 387502 532894
rect 387586 532658 387822 532894
rect 387266 532338 387502 532574
rect 387586 532338 387822 532574
rect 387266 496658 387502 496894
rect 387586 496658 387822 496894
rect 387266 496338 387502 496574
rect 387586 496338 387822 496574
rect 387266 460658 387502 460894
rect 387586 460658 387822 460894
rect 387266 460338 387502 460574
rect 387586 460338 387822 460574
rect 387266 424658 387502 424894
rect 387586 424658 387822 424894
rect 387266 424338 387502 424574
rect 387586 424338 387822 424574
rect 387266 388658 387502 388894
rect 387586 388658 387822 388894
rect 387266 388338 387502 388574
rect 387586 388338 387822 388574
rect 387266 352658 387502 352894
rect 387586 352658 387822 352894
rect 387266 352338 387502 352574
rect 387586 352338 387822 352574
rect 387266 316658 387502 316894
rect 387586 316658 387822 316894
rect 387266 316338 387502 316574
rect 387586 316338 387822 316574
rect 387266 280658 387502 280894
rect 387586 280658 387822 280894
rect 387266 280338 387502 280574
rect 387586 280338 387822 280574
rect 387266 244658 387502 244894
rect 387586 244658 387822 244894
rect 387266 244338 387502 244574
rect 387586 244338 387822 244574
rect 387266 208658 387502 208894
rect 387586 208658 387822 208894
rect 387266 208338 387502 208574
rect 387586 208338 387822 208574
rect 387266 172658 387502 172894
rect 387586 172658 387822 172894
rect 387266 172338 387502 172574
rect 387586 172338 387822 172574
rect 387266 136658 387502 136894
rect 387586 136658 387822 136894
rect 387266 136338 387502 136574
rect 387586 136338 387822 136574
rect 387266 100658 387502 100894
rect 387586 100658 387822 100894
rect 387266 100338 387502 100574
rect 387586 100338 387822 100574
rect 387266 64658 387502 64894
rect 387586 64658 387822 64894
rect 387266 64338 387502 64574
rect 387586 64338 387822 64574
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 390986 536378 391222 536614
rect 391306 536378 391542 536614
rect 390986 536058 391222 536294
rect 391306 536058 391542 536294
rect 390986 500378 391222 500614
rect 391306 500378 391542 500614
rect 390986 500058 391222 500294
rect 391306 500058 391542 500294
rect 390986 464378 391222 464614
rect 391306 464378 391542 464614
rect 390986 464058 391222 464294
rect 391306 464058 391542 464294
rect 390986 428378 391222 428614
rect 391306 428378 391542 428614
rect 390986 428058 391222 428294
rect 391306 428058 391542 428294
rect 390986 392378 391222 392614
rect 391306 392378 391542 392614
rect 390986 392058 391222 392294
rect 391306 392058 391542 392294
rect 390986 356378 391222 356614
rect 391306 356378 391542 356614
rect 390986 356058 391222 356294
rect 391306 356058 391542 356294
rect 390986 320378 391222 320614
rect 391306 320378 391542 320614
rect 390986 320058 391222 320294
rect 391306 320058 391542 320294
rect 390986 284378 391222 284614
rect 391306 284378 391542 284614
rect 390986 284058 391222 284294
rect 391306 284058 391542 284294
rect 390986 248378 391222 248614
rect 391306 248378 391542 248614
rect 390986 248058 391222 248294
rect 391306 248058 391542 248294
rect 390986 212378 391222 212614
rect 391306 212378 391542 212614
rect 390986 212058 391222 212294
rect 391306 212058 391542 212294
rect 390986 176378 391222 176614
rect 391306 176378 391542 176614
rect 390986 176058 391222 176294
rect 391306 176058 391542 176294
rect 390986 140378 391222 140614
rect 391306 140378 391542 140614
rect 390986 140058 391222 140294
rect 391306 140058 391542 140294
rect 390986 104378 391222 104614
rect 391306 104378 391542 104614
rect 390986 104058 391222 104294
rect 391306 104058 391542 104294
rect 390986 68378 391222 68614
rect 391306 68378 391542 68614
rect 390986 68058 391222 68294
rect 391306 68058 391542 68294
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 401546 438938 401782 439174
rect 401866 438938 402102 439174
rect 401546 438618 401782 438854
rect 401866 438618 402102 438854
rect 401546 402938 401782 403174
rect 401866 402938 402102 403174
rect 401546 402618 401782 402854
rect 401866 402618 402102 402854
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 401546 330938 401782 331174
rect 401866 330938 402102 331174
rect 401546 330618 401782 330854
rect 401866 330618 402102 330854
rect 401546 294938 401782 295174
rect 401866 294938 402102 295174
rect 401546 294618 401782 294854
rect 401866 294618 402102 294854
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 401546 222938 401782 223174
rect 401866 222938 402102 223174
rect 401546 222618 401782 222854
rect 401866 222618 402102 222854
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 405266 442658 405502 442894
rect 405586 442658 405822 442894
rect 405266 442338 405502 442574
rect 405586 442338 405822 442574
rect 405266 406658 405502 406894
rect 405586 406658 405822 406894
rect 405266 406338 405502 406574
rect 405586 406338 405822 406574
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 405266 334658 405502 334894
rect 405586 334658 405822 334894
rect 405266 334338 405502 334574
rect 405586 334338 405822 334574
rect 405266 298658 405502 298894
rect 405586 298658 405822 298894
rect 405266 298338 405502 298574
rect 405586 298338 405822 298574
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 405266 226658 405502 226894
rect 405586 226658 405822 226894
rect 405266 226338 405502 226574
rect 405586 226338 405822 226574
rect 405266 190658 405502 190894
rect 405586 190658 405822 190894
rect 405266 190338 405502 190574
rect 405586 190338 405822 190574
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 405266 118658 405502 118894
rect 405586 118658 405822 118894
rect 405266 118338 405502 118574
rect 405586 118338 405822 118574
rect 405266 82658 405502 82894
rect 405586 82658 405822 82894
rect 405266 82338 405502 82574
rect 405586 82338 405822 82574
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 408986 446378 409222 446614
rect 409306 446378 409542 446614
rect 408986 446058 409222 446294
rect 409306 446058 409542 446294
rect 408986 410378 409222 410614
rect 409306 410378 409542 410614
rect 408986 410058 409222 410294
rect 409306 410058 409542 410294
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 408986 338378 409222 338614
rect 409306 338378 409542 338614
rect 408986 338058 409222 338294
rect 409306 338058 409542 338294
rect 408986 302378 409222 302614
rect 409306 302378 409542 302614
rect 408986 302058 409222 302294
rect 409306 302058 409542 302294
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 408986 230378 409222 230614
rect 409306 230378 409542 230614
rect 408986 230058 409222 230294
rect 409306 230058 409542 230294
rect 408986 194378 409222 194614
rect 409306 194378 409542 194614
rect 408986 194058 409222 194294
rect 409306 194058 409542 194294
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 408986 86378 409222 86614
rect 409306 86378 409542 86614
rect 408986 86058 409222 86294
rect 409306 86058 409542 86294
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 419546 564938 419782 565174
rect 419866 564938 420102 565174
rect 419546 564618 419782 564854
rect 419866 564618 420102 564854
rect 419546 528938 419782 529174
rect 419866 528938 420102 529174
rect 419546 528618 419782 528854
rect 419866 528618 420102 528854
rect 419546 492938 419782 493174
rect 419866 492938 420102 493174
rect 419546 492618 419782 492854
rect 419866 492618 420102 492854
rect 419546 456938 419782 457174
rect 419866 456938 420102 457174
rect 419546 456618 419782 456854
rect 419866 456618 420102 456854
rect 419546 420938 419782 421174
rect 419866 420938 420102 421174
rect 419546 420618 419782 420854
rect 419866 420618 420102 420854
rect 419546 384938 419782 385174
rect 419866 384938 420102 385174
rect 419546 384618 419782 384854
rect 419866 384618 420102 384854
rect 419546 348938 419782 349174
rect 419866 348938 420102 349174
rect 419546 348618 419782 348854
rect 419866 348618 420102 348854
rect 419546 312938 419782 313174
rect 419866 312938 420102 313174
rect 419546 312618 419782 312854
rect 419866 312618 420102 312854
rect 419546 276938 419782 277174
rect 419866 276938 420102 277174
rect 419546 276618 419782 276854
rect 419866 276618 420102 276854
rect 419546 240938 419782 241174
rect 419866 240938 420102 241174
rect 419546 240618 419782 240854
rect 419866 240618 420102 240854
rect 419546 204938 419782 205174
rect 419866 204938 420102 205174
rect 419546 204618 419782 204854
rect 419866 204618 420102 204854
rect 419546 168938 419782 169174
rect 419866 168938 420102 169174
rect 419546 168618 419782 168854
rect 419866 168618 420102 168854
rect 419546 132938 419782 133174
rect 419866 132938 420102 133174
rect 419546 132618 419782 132854
rect 419866 132618 420102 132854
rect 419546 96938 419782 97174
rect 419866 96938 420102 97174
rect 419546 96618 419782 96854
rect 419866 96618 420102 96854
rect 419546 60938 419782 61174
rect 419866 60938 420102 61174
rect 419546 60618 419782 60854
rect 419866 60618 420102 60854
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 423266 568658 423502 568894
rect 423586 568658 423822 568894
rect 423266 568338 423502 568574
rect 423586 568338 423822 568574
rect 423266 532658 423502 532894
rect 423586 532658 423822 532894
rect 423266 532338 423502 532574
rect 423586 532338 423822 532574
rect 423266 496658 423502 496894
rect 423586 496658 423822 496894
rect 423266 496338 423502 496574
rect 423586 496338 423822 496574
rect 423266 460658 423502 460894
rect 423586 460658 423822 460894
rect 423266 460338 423502 460574
rect 423586 460338 423822 460574
rect 423266 424658 423502 424894
rect 423586 424658 423822 424894
rect 423266 424338 423502 424574
rect 423586 424338 423822 424574
rect 423266 388658 423502 388894
rect 423586 388658 423822 388894
rect 423266 388338 423502 388574
rect 423586 388338 423822 388574
rect 423266 352658 423502 352894
rect 423586 352658 423822 352894
rect 423266 352338 423502 352574
rect 423586 352338 423822 352574
rect 423266 316658 423502 316894
rect 423586 316658 423822 316894
rect 423266 316338 423502 316574
rect 423586 316338 423822 316574
rect 423266 280658 423502 280894
rect 423586 280658 423822 280894
rect 423266 280338 423502 280574
rect 423586 280338 423822 280574
rect 423266 244658 423502 244894
rect 423586 244658 423822 244894
rect 423266 244338 423502 244574
rect 423586 244338 423822 244574
rect 423266 208658 423502 208894
rect 423586 208658 423822 208894
rect 423266 208338 423502 208574
rect 423586 208338 423822 208574
rect 423266 172658 423502 172894
rect 423586 172658 423822 172894
rect 423266 172338 423502 172574
rect 423586 172338 423822 172574
rect 423266 136658 423502 136894
rect 423586 136658 423822 136894
rect 423266 136338 423502 136574
rect 423586 136338 423822 136574
rect 423266 100658 423502 100894
rect 423586 100658 423822 100894
rect 423266 100338 423502 100574
rect 423586 100338 423822 100574
rect 423266 64658 423502 64894
rect 423586 64658 423822 64894
rect 423266 64338 423502 64574
rect 423586 64338 423822 64574
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 426986 572378 427222 572614
rect 427306 572378 427542 572614
rect 426986 572058 427222 572294
rect 427306 572058 427542 572294
rect 426986 536378 427222 536614
rect 427306 536378 427542 536614
rect 426986 536058 427222 536294
rect 427306 536058 427542 536294
rect 426986 500378 427222 500614
rect 427306 500378 427542 500614
rect 426986 500058 427222 500294
rect 427306 500058 427542 500294
rect 426986 464378 427222 464614
rect 427306 464378 427542 464614
rect 426986 464058 427222 464294
rect 427306 464058 427542 464294
rect 426986 428378 427222 428614
rect 427306 428378 427542 428614
rect 426986 428058 427222 428294
rect 427306 428058 427542 428294
rect 426986 392378 427222 392614
rect 427306 392378 427542 392614
rect 426986 392058 427222 392294
rect 427306 392058 427542 392294
rect 426986 356378 427222 356614
rect 427306 356378 427542 356614
rect 426986 356058 427222 356294
rect 427306 356058 427542 356294
rect 426986 320378 427222 320614
rect 427306 320378 427542 320614
rect 426986 320058 427222 320294
rect 427306 320058 427542 320294
rect 426986 284378 427222 284614
rect 427306 284378 427542 284614
rect 426986 284058 427222 284294
rect 427306 284058 427542 284294
rect 426986 248378 427222 248614
rect 427306 248378 427542 248614
rect 426986 248058 427222 248294
rect 427306 248058 427542 248294
rect 426986 212378 427222 212614
rect 427306 212378 427542 212614
rect 426986 212058 427222 212294
rect 427306 212058 427542 212294
rect 426986 176378 427222 176614
rect 427306 176378 427542 176614
rect 426986 176058 427222 176294
rect 427306 176058 427542 176294
rect 426986 140378 427222 140614
rect 427306 140378 427542 140614
rect 426986 140058 427222 140294
rect 427306 140058 427542 140294
rect 426986 104378 427222 104614
rect 427306 104378 427542 104614
rect 426986 104058 427222 104294
rect 427306 104058 427542 104294
rect 426986 68378 427222 68614
rect 427306 68378 427542 68614
rect 426986 68058 427222 68294
rect 427306 68058 427542 68294
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 437546 438938 437782 439174
rect 437866 438938 438102 439174
rect 437546 438618 437782 438854
rect 437866 438618 438102 438854
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 437546 294938 437782 295174
rect 437866 294938 438102 295174
rect 437546 294618 437782 294854
rect 437866 294618 438102 294854
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 437546 114938 437782 115174
rect 437866 114938 438102 115174
rect 437546 114618 437782 114854
rect 437866 114618 438102 114854
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 441266 442658 441502 442894
rect 441586 442658 441822 442894
rect 441266 442338 441502 442574
rect 441586 442338 441822 442574
rect 441266 406658 441502 406894
rect 441586 406658 441822 406894
rect 441266 406338 441502 406574
rect 441586 406338 441822 406574
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 441266 334658 441502 334894
rect 441586 334658 441822 334894
rect 441266 334338 441502 334574
rect 441586 334338 441822 334574
rect 441266 298658 441502 298894
rect 441586 298658 441822 298894
rect 441266 298338 441502 298574
rect 441586 298338 441822 298574
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 441266 226658 441502 226894
rect 441586 226658 441822 226894
rect 441266 226338 441502 226574
rect 441586 226338 441822 226574
rect 441266 190658 441502 190894
rect 441586 190658 441822 190894
rect 441266 190338 441502 190574
rect 441586 190338 441822 190574
rect 441266 154658 441502 154894
rect 441586 154658 441822 154894
rect 441266 154338 441502 154574
rect 441586 154338 441822 154574
rect 441266 118658 441502 118894
rect 441586 118658 441822 118894
rect 441266 118338 441502 118574
rect 441586 118338 441822 118574
rect 441266 82658 441502 82894
rect 441586 82658 441822 82894
rect 441266 82338 441502 82574
rect 441586 82338 441822 82574
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 444986 410378 445222 410614
rect 445306 410378 445542 410614
rect 444986 410058 445222 410294
rect 445306 410058 445542 410294
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 444986 302378 445222 302614
rect 445306 302378 445542 302614
rect 444986 302058 445222 302294
rect 445306 302058 445542 302294
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 444986 122378 445222 122614
rect 445306 122378 445542 122614
rect 444986 122058 445222 122294
rect 445306 122058 445542 122294
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 455546 528938 455782 529174
rect 455866 528938 456102 529174
rect 455546 528618 455782 528854
rect 455866 528618 456102 528854
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 455546 456938 455782 457174
rect 455866 456938 456102 457174
rect 455546 456618 455782 456854
rect 455866 456618 456102 456854
rect 455546 420938 455782 421174
rect 455866 420938 456102 421174
rect 455546 420618 455782 420854
rect 455866 420618 456102 420854
rect 455546 384938 455782 385174
rect 455866 384938 456102 385174
rect 455546 384618 455782 384854
rect 455866 384618 456102 384854
rect 455546 348938 455782 349174
rect 455866 348938 456102 349174
rect 455546 348618 455782 348854
rect 455866 348618 456102 348854
rect 455546 312938 455782 313174
rect 455866 312938 456102 313174
rect 455546 312618 455782 312854
rect 455866 312618 456102 312854
rect 455546 276938 455782 277174
rect 455866 276938 456102 277174
rect 455546 276618 455782 276854
rect 455866 276618 456102 276854
rect 455546 240938 455782 241174
rect 455866 240938 456102 241174
rect 455546 240618 455782 240854
rect 455866 240618 456102 240854
rect 455546 204938 455782 205174
rect 455866 204938 456102 205174
rect 455546 204618 455782 204854
rect 455866 204618 456102 204854
rect 455546 168938 455782 169174
rect 455866 168938 456102 169174
rect 455546 168618 455782 168854
rect 455866 168618 456102 168854
rect 455546 132938 455782 133174
rect 455866 132938 456102 133174
rect 455546 132618 455782 132854
rect 455866 132618 456102 132854
rect 455546 96938 455782 97174
rect 455866 96938 456102 97174
rect 455546 96618 455782 96854
rect 455866 96618 456102 96854
rect 455546 60938 455782 61174
rect 455866 60938 456102 61174
rect 455546 60618 455782 60854
rect 455866 60618 456102 60854
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 459266 532658 459502 532894
rect 459586 532658 459822 532894
rect 459266 532338 459502 532574
rect 459586 532338 459822 532574
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 459266 460658 459502 460894
rect 459586 460658 459822 460894
rect 459266 460338 459502 460574
rect 459586 460338 459822 460574
rect 459266 424658 459502 424894
rect 459586 424658 459822 424894
rect 459266 424338 459502 424574
rect 459586 424338 459822 424574
rect 459266 388658 459502 388894
rect 459586 388658 459822 388894
rect 459266 388338 459502 388574
rect 459586 388338 459822 388574
rect 459266 352658 459502 352894
rect 459586 352658 459822 352894
rect 459266 352338 459502 352574
rect 459586 352338 459822 352574
rect 459266 316658 459502 316894
rect 459586 316658 459822 316894
rect 459266 316338 459502 316574
rect 459586 316338 459822 316574
rect 459266 280658 459502 280894
rect 459586 280658 459822 280894
rect 459266 280338 459502 280574
rect 459586 280338 459822 280574
rect 459266 244658 459502 244894
rect 459586 244658 459822 244894
rect 459266 244338 459502 244574
rect 459586 244338 459822 244574
rect 459266 208658 459502 208894
rect 459586 208658 459822 208894
rect 459266 208338 459502 208574
rect 459586 208338 459822 208574
rect 459266 172658 459502 172894
rect 459586 172658 459822 172894
rect 459266 172338 459502 172574
rect 459586 172338 459822 172574
rect 459266 136658 459502 136894
rect 459586 136658 459822 136894
rect 459266 136338 459502 136574
rect 459586 136338 459822 136574
rect 459266 100658 459502 100894
rect 459586 100658 459822 100894
rect 459266 100338 459502 100574
rect 459586 100338 459822 100574
rect 459266 64658 459502 64894
rect 459586 64658 459822 64894
rect 459266 64338 459502 64574
rect 459586 64338 459822 64574
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 462986 536378 463222 536614
rect 463306 536378 463542 536614
rect 462986 536058 463222 536294
rect 463306 536058 463542 536294
rect 462986 500378 463222 500614
rect 463306 500378 463542 500614
rect 462986 500058 463222 500294
rect 463306 500058 463542 500294
rect 462986 464378 463222 464614
rect 463306 464378 463542 464614
rect 462986 464058 463222 464294
rect 463306 464058 463542 464294
rect 462986 428378 463222 428614
rect 463306 428378 463542 428614
rect 462986 428058 463222 428294
rect 463306 428058 463542 428294
rect 462986 392378 463222 392614
rect 463306 392378 463542 392614
rect 462986 392058 463222 392294
rect 463306 392058 463542 392294
rect 462986 356378 463222 356614
rect 463306 356378 463542 356614
rect 462986 356058 463222 356294
rect 463306 356058 463542 356294
rect 462986 320378 463222 320614
rect 463306 320378 463542 320614
rect 462986 320058 463222 320294
rect 463306 320058 463542 320294
rect 462986 284378 463222 284614
rect 463306 284378 463542 284614
rect 462986 284058 463222 284294
rect 463306 284058 463542 284294
rect 462986 248378 463222 248614
rect 463306 248378 463542 248614
rect 462986 248058 463222 248294
rect 463306 248058 463542 248294
rect 462986 212378 463222 212614
rect 463306 212378 463542 212614
rect 462986 212058 463222 212294
rect 463306 212058 463542 212294
rect 462986 176378 463222 176614
rect 463306 176378 463542 176614
rect 462986 176058 463222 176294
rect 463306 176058 463542 176294
rect 462986 140378 463222 140614
rect 463306 140378 463542 140614
rect 462986 140058 463222 140294
rect 463306 140058 463542 140294
rect 462986 104378 463222 104614
rect 463306 104378 463542 104614
rect 462986 104058 463222 104294
rect 463306 104058 463542 104294
rect 462986 68378 463222 68614
rect 463306 68378 463542 68614
rect 462986 68058 463222 68294
rect 463306 68058 463542 68294
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 477266 334658 477502 334894
rect 477586 334658 477822 334894
rect 477266 334338 477502 334574
rect 477586 334338 477822 334574
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 477266 226658 477502 226894
rect 477586 226658 477822 226894
rect 477266 226338 477502 226574
rect 477586 226338 477822 226574
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 480986 410378 481222 410614
rect 481306 410378 481542 410614
rect 480986 410058 481222 410294
rect 481306 410058 481542 410294
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 480986 338378 481222 338614
rect 481306 338378 481542 338614
rect 480986 338058 481222 338294
rect 481306 338058 481542 338294
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 491546 456938 491782 457174
rect 491866 456938 492102 457174
rect 491546 456618 491782 456854
rect 491866 456618 492102 456854
rect 491546 420938 491782 421174
rect 491866 420938 492102 421174
rect 491546 420618 491782 420854
rect 491866 420618 492102 420854
rect 491546 384938 491782 385174
rect 491866 384938 492102 385174
rect 491546 384618 491782 384854
rect 491866 384618 492102 384854
rect 491546 348938 491782 349174
rect 491866 348938 492102 349174
rect 491546 348618 491782 348854
rect 491866 348618 492102 348854
rect 491546 312938 491782 313174
rect 491866 312938 492102 313174
rect 491546 312618 491782 312854
rect 491866 312618 492102 312854
rect 491546 276938 491782 277174
rect 491866 276938 492102 277174
rect 491546 276618 491782 276854
rect 491866 276618 492102 276854
rect 491546 240938 491782 241174
rect 491866 240938 492102 241174
rect 491546 240618 491782 240854
rect 491866 240618 492102 240854
rect 491546 204938 491782 205174
rect 491866 204938 492102 205174
rect 491546 204618 491782 204854
rect 491866 204618 492102 204854
rect 491546 168938 491782 169174
rect 491866 168938 492102 169174
rect 491546 168618 491782 168854
rect 491866 168618 492102 168854
rect 491546 132938 491782 133174
rect 491866 132938 492102 133174
rect 491546 132618 491782 132854
rect 491866 132618 492102 132854
rect 491546 96938 491782 97174
rect 491866 96938 492102 97174
rect 491546 96618 491782 96854
rect 491866 96618 492102 96854
rect 491546 60938 491782 61174
rect 491866 60938 492102 61174
rect 491546 60618 491782 60854
rect 491866 60618 492102 60854
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 495266 460658 495502 460894
rect 495586 460658 495822 460894
rect 495266 460338 495502 460574
rect 495586 460338 495822 460574
rect 495266 424658 495502 424894
rect 495586 424658 495822 424894
rect 495266 424338 495502 424574
rect 495586 424338 495822 424574
rect 495266 388658 495502 388894
rect 495586 388658 495822 388894
rect 495266 388338 495502 388574
rect 495586 388338 495822 388574
rect 495266 352658 495502 352894
rect 495586 352658 495822 352894
rect 495266 352338 495502 352574
rect 495586 352338 495822 352574
rect 495266 316658 495502 316894
rect 495586 316658 495822 316894
rect 495266 316338 495502 316574
rect 495586 316338 495822 316574
rect 495266 280658 495502 280894
rect 495586 280658 495822 280894
rect 495266 280338 495502 280574
rect 495586 280338 495822 280574
rect 495266 244658 495502 244894
rect 495586 244658 495822 244894
rect 495266 244338 495502 244574
rect 495586 244338 495822 244574
rect 495266 208658 495502 208894
rect 495586 208658 495822 208894
rect 495266 208338 495502 208574
rect 495586 208338 495822 208574
rect 495266 172658 495502 172894
rect 495586 172658 495822 172894
rect 495266 172338 495502 172574
rect 495586 172338 495822 172574
rect 495266 136658 495502 136894
rect 495586 136658 495822 136894
rect 495266 136338 495502 136574
rect 495586 136338 495822 136574
rect 495266 100658 495502 100894
rect 495586 100658 495822 100894
rect 495266 100338 495502 100574
rect 495586 100338 495822 100574
rect 495266 64658 495502 64894
rect 495586 64658 495822 64894
rect 495266 64338 495502 64574
rect 495586 64338 495822 64574
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 498986 608378 499222 608614
rect 499306 608378 499542 608614
rect 498986 608058 499222 608294
rect 499306 608058 499542 608294
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 498986 464378 499222 464614
rect 499306 464378 499542 464614
rect 498986 464058 499222 464294
rect 499306 464058 499542 464294
rect 498986 428378 499222 428614
rect 499306 428378 499542 428614
rect 498986 428058 499222 428294
rect 499306 428058 499542 428294
rect 498986 392378 499222 392614
rect 499306 392378 499542 392614
rect 498986 392058 499222 392294
rect 499306 392058 499542 392294
rect 498986 356378 499222 356614
rect 499306 356378 499542 356614
rect 498986 356058 499222 356294
rect 499306 356058 499542 356294
rect 498986 320378 499222 320614
rect 499306 320378 499542 320614
rect 498986 320058 499222 320294
rect 499306 320058 499542 320294
rect 498986 284378 499222 284614
rect 499306 284378 499542 284614
rect 498986 284058 499222 284294
rect 499306 284058 499542 284294
rect 498986 248378 499222 248614
rect 499306 248378 499542 248614
rect 498986 248058 499222 248294
rect 499306 248058 499542 248294
rect 498986 212378 499222 212614
rect 499306 212378 499542 212614
rect 498986 212058 499222 212294
rect 499306 212058 499542 212294
rect 498986 176378 499222 176614
rect 499306 176378 499542 176614
rect 498986 176058 499222 176294
rect 499306 176058 499542 176294
rect 498986 140378 499222 140614
rect 499306 140378 499542 140614
rect 498986 140058 499222 140294
rect 499306 140058 499542 140294
rect 498986 104378 499222 104614
rect 499306 104378 499542 104614
rect 498986 104058 499222 104294
rect 499306 104058 499542 104294
rect 498986 68378 499222 68614
rect 499306 68378 499542 68614
rect 498986 68058 499222 68294
rect 499306 68058 499542 68294
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 77686 561454
rect 77922 561218 85617 561454
rect 85853 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 77686 561134
rect 77922 560898 85617 561134
rect 85853 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73721 543454
rect 73957 543218 81651 543454
rect 81887 543218 89582 543454
rect 89818 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73721 543134
rect 73957 542898 81651 543134
rect 81887 542898 89582 543134
rect 89818 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 88380 417454
rect 88616 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 88380 417134
rect 88616 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73020 399454
rect 73256 399218 103740 399454
rect 103976 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73020 399134
rect 73256 398898 103740 399134
rect 103976 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 197818 291454
rect 198054 291218 228538 291454
rect 228774 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 197818 291134
rect 198054 290898 228538 291134
rect 228774 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 79019 273454
rect 79255 273218 88283 273454
rect 88519 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 213178 273454
rect 213414 273218 243898 273454
rect 244134 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 79019 273134
rect 79255 272898 88283 273134
rect 88519 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 213178 273134
rect 213414 272898 243898 273134
rect 244134 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 74387 255454
rect 74623 255218 83651 255454
rect 83887 255218 92915 255454
rect 93151 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 197818 255454
rect 198054 255218 228538 255454
rect 228774 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 74387 255134
rect 74623 254898 83651 255134
rect 83887 254898 92915 255134
rect 93151 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 197818 255134
rect 198054 254898 228538 255134
rect 228774 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 102986 176614
rect 103222 176378 103306 176614
rect 103542 176378 138986 176614
rect 139222 176378 139306 176614
rect 139542 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 102986 176294
rect 103222 176058 103306 176294
rect 103542 176058 138986 176294
rect 139222 176058 139306 176294
rect 139542 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 99266 172894
rect 99502 172658 99586 172894
rect 99822 172658 135266 172894
rect 135502 172658 135586 172894
rect 135822 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 279266 172894
rect 279502 172658 279586 172894
rect 279822 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 99266 172574
rect 99502 172338 99586 172574
rect 99822 172338 135266 172574
rect 135502 172338 135586 172574
rect 135822 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 279266 172574
rect 279502 172338 279586 172574
rect 279822 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 95546 169174
rect 95782 168938 95866 169174
rect 96102 168938 131546 169174
rect 131782 168938 131866 169174
rect 132102 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 275546 169174
rect 275782 168938 275866 169174
rect 276102 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 95546 168854
rect 95782 168618 95866 168854
rect 96102 168618 131546 168854
rect 131782 168618 131866 168854
rect 132102 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 275546 168854
rect 275782 168618 275866 168854
rect 276102 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 102986 140614
rect 103222 140378 103306 140614
rect 103542 140378 138986 140614
rect 139222 140378 139306 140614
rect 139542 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 102986 140294
rect 103222 140058 103306 140294
rect 103542 140058 138986 140294
rect 139222 140058 139306 140294
rect 139542 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 99266 136894
rect 99502 136658 99586 136894
rect 99822 136658 135266 136894
rect 135502 136658 135586 136894
rect 135822 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 279266 136894
rect 279502 136658 279586 136894
rect 279822 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 99266 136574
rect 99502 136338 99586 136574
rect 99822 136338 135266 136574
rect 135502 136338 135586 136574
rect 135822 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 279266 136574
rect 279502 136338 279586 136574
rect 279822 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 131546 133174
rect 131782 132938 131866 133174
rect 132102 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 131546 132854
rect 131782 132618 131866 132854
rect 132102 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 77686 129454
rect 77922 129218 85617 129454
rect 85853 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 204306 129454
rect 204542 129218 214058 129454
rect 214294 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 77686 129134
rect 77922 128898 85617 129134
rect 85853 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 204306 129134
rect 204542 128898 214058 129134
rect 214294 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73721 111454
rect 73957 111218 81651 111454
rect 81887 111218 89582 111454
rect 89818 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 199430 111454
rect 199666 111218 209182 111454
rect 209418 111218 218934 111454
rect 219170 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73721 111134
rect 73957 110898 81651 111134
rect 81887 110898 89582 111134
rect 89818 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 199430 111134
rect 199666 110898 209182 111134
rect 209418 110898 218934 111134
rect 219170 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 102986 104614
rect 103222 104378 103306 104614
rect 103542 104378 138986 104614
rect 139222 104378 139306 104614
rect 139542 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 102986 104294
rect 103222 104058 103306 104294
rect 103542 104058 138986 104294
rect 139222 104058 139306 104294
rect 139542 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 99266 100894
rect 99502 100658 99586 100894
rect 99822 100658 135266 100894
rect 135502 100658 135586 100894
rect 135822 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 279266 100894
rect 279502 100658 279586 100894
rect 279822 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 99266 100574
rect 99502 100338 99586 100574
rect 99822 100338 135266 100574
rect 135502 100338 135586 100574
rect 135822 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 279266 100574
rect 279502 100338 279586 100574
rect 279822 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 131546 97174
rect 131782 96938 131866 97174
rect 132102 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 131546 96854
rect 131782 96618 131866 96854
rect 132102 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use zube_wrapped_project  zube_wrapped_project_5
timestamp 1635266113
transform 1 0 193568 0 1 241592
box 0 0 60000 60000
use wrapped_ws2812  wrapped_ws2812_4
timestamp 1635266113
transform 1 0 193568 0 1 92782
box 0 0 31475 48253
use wrapped_vga_clock  wrapped_vga_clock_2
timestamp 1635266113
transform 1 0 68770 0 1 390356
box 0 0 44000 44000
use wrapped_tpm2137  wrapped_tpm2137_3
timestamp 1635266113
transform 1 0 68770 0 1 539166
box 0 0 26000 42000
use wrapped_rgb_mixer  wrapped_rgb_mixer_0
timestamp 1635266113
transform 1 0 68770 0 1 92782
box 0 0 26000 42000
use wrapped_frequency_counter  wrapped_frequency_counter_1
timestamp 1635266113
transform 1 0 68770 0 1 241592
box 0 0 30000 42000
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 90782 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 90782 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 136782 74414 239592 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 143035 218414 239592 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 239592 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 285592 74414 388356 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 388356 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 436356 74414 537166 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 583166 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 436356 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 303592 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 303592 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 90782 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 90782 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 136782 78134 239592 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 143035 222134 239592 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 285592 78134 388356 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 388356 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 436356 78134 537166 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 583166 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 436356 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 303592 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 90782 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 90782 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 136782 81854 239592 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 143035 225854 239592 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 285592 81854 388356 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 436356 81854 537166 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 583166 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 303592 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 90782 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 90782 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 136782 85574 239592 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 143035 193574 239592 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 239592 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 285592 85574 388356 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 436356 85574 537166 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 583166 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 303592 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 303592 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 90782 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 239592 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 143035 207854 239592 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 239592 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 285592 99854 388356 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 436356 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 303592 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 303592 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 90782 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 90782 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 136782 67574 239592 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 143035 211574 239592 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 239592 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 285592 67574 388356 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 388356 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 436356 67574 537166 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 583166 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 436356 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 303592 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 303592 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 90782 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 90782 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 136782 92414 239592 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 143035 200414 239592 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 239592 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 285592 92414 388356 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 436356 92414 537166 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 583166 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 303592 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 303592 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 90782 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 90782 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 136782 96134 239592 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 143035 204134 239592 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 239592 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 285592 96134 388356 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 436356 96134 537166 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 583166 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 303592 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 303592 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
